// Generator : SpinalHDL dev    git head : c796d9fc761d68c4391d98f72d852457e34aeb32
// Component : EndeavourSoc
// Git hash  : 7bccf9e9ef87ac7526360a482416657e6df0b62b

`timescale 1ns/1ps

module EndeavourSoc (
  input  wire          io_nreset,
  input  wire          io_clk_in,
  output wire          io_plla_i2c_scl,
  inout  wire          io_plla_i2c_sda,
  input  wire          io_plla_clk0,
  input  wire          io_plla_clk1,
  input  wire          io_plla_clk2,
  output wire          io_pllb_i2c_scl,
  inout  wire          io_pllb_i2c_sda,
  input  wire          io_pllb_clk0,
  input  wire          io_pllb_clk1,
  input  wire          io_pllb_clk2,
  output wire [2:0]    io_leds,
  input  wire [1:0]    io_keys,
  output wire          io_audio_shdn,
  output wire          io_audio_i2c_scl,
  inout  wire          io_audio_i2c_sda,
  input  wire          io_uart_rx,
  output wire          io_uart_tx,
  output wire          io_dvi_tmds0p,
  output wire          io_dvi_tmds0m,
  output wire          io_dvi_tmds1p,
  output wire          io_dvi_tmds1m,
  output wire          io_dvi_tmds2p,
  output wire          io_dvi_tmds2m,
  output wire          io_dvi_tmdsCp,
  output wire          io_dvi_tmdsCm,
  output wire          io_sdcard_clk,
  inout  wire          io_sdcard_cmd,
  inout  wire [3:0]    io_sdcard_data,
  input  wire          io_sdcard_ndetect,
  output wire          io_ddr_sdram_ck_p,
  output wire          io_ddr_sdram_ck_n,
  output wire          io_ddr_sdram_cke,
  output wire          io_ddr_sdram_ras_n,
  output wire          io_ddr_sdram_cas_n,
  output wire          io_ddr_sdram_we_n,
  output wire [1:0]    io_ddr_sdram_ba,
  output wire [13:0]   io_ddr_sdram_a,
  output wire [1:0]    io_ddr_sdram_dm,
  inout  wire [1:0]    io_ddr_sdram_dqs,
  inout  wire [15:0]   io_ddr_sdram_dq,
  inout  wire          io_usb1_dp,
  inout  wire          io_usb1_dn,
  inout  wire          io_usb2_dp,
  inout  wire          io_usb2_dn
);
  localparam A_PUT_FULL_DATA = 3'd0;
  localparam A_PUT_PARTIAL_DATA = 3'd1;
  localparam A_GET = 3'd4;
  localparam A_ACQUIRE_BLOCK = 3'd6;
  localparam A_ACQUIRE_PERM = 3'd7;
  localparam D_ACCESS_ACK = 3'd0;
  localparam D_ACCESS_ACK_DATA = 3'd1;
  localparam D_GRANT = 3'd4;
  localparam D_GRANT_DATA = 3'd5;
  localparam D_RELEASE_ACK = 3'd6;

  wire       [4:0]    board_ctrl_apb_PADDR;
  wire       [4:0]    video_ctrl_apb_PADDR;
  wire       [3:0]    peripheral_uart_ctrl_apb_PADDR;
  wire       [2:0]    peripheral_audio_ctrl_apb_PADDR;
  wire       [4:0]    peripheral_sdcard_ctrl_apb_PADDR;
  wire       [11:0]   peripheral_usb_ctrl_io_apb_ctrl_PADDR;
  wire       [11:0]   peripheral_usb_ctrl_io_apb_dma_PADDR;
  wire       [18:0]   peripheral_apb_bridge_input_PADDR;
  wire                vexiiRiscv_1_PrivilegedPlugin_logic_harts_0_int_m_timer;
  wire                vexiiRiscv_1_PrivilegedPlugin_logic_harts_0_int_m_software;
  wire                vexiiRiscv_1_PrivilegedPlugin_logic_harts_0_int_m_external;
  wire                vexiiRiscv_1_PrivilegedPlugin_logic_harts_0_int_s_external;
  wire                board_ctrl_plla_i2c_scl;
  wire                board_ctrl_pllb_i2c_scl;
  wire                board_ctrl_reset_cpu;
  wire                board_ctrl_reset_ram;
  wire                board_ctrl_reset_peripheral;
  wire                board_ctrl_clk_cpu;
  wire                board_ctrl_clk_ram;
  wire                board_ctrl_clk_ram_bus;
  wire                board_ctrl_clk_peripheral;
  wire       [63:0]   board_ctrl_utime;
  wire                board_ctrl_timer_interrupt;
  wire                board_ctrl_clk_tmds_pixel;
  wire                board_ctrl_clk_tmds_x5;
  wire       [2:0]    board_ctrl_leds;
  wire                board_ctrl_apb_PREADY;
  wire       [31:0]   board_ctrl_apb_PRDATA;
  wire       [1:0]    video_ctrl_video_mode_out;
  wire                video_ctrl_dvi_tmds0p;
  wire                video_ctrl_dvi_tmds0m;
  wire                video_ctrl_dvi_tmds1p;
  wire                video_ctrl_dvi_tmds1m;
  wire                video_ctrl_dvi_tmds2p;
  wire                video_ctrl_dvi_tmds2m;
  wire                video_ctrl_dvi_tmdsCp;
  wire                video_ctrl_dvi_tmdsCm;
  wire                video_ctrl_apb_PREADY;
  wire       [31:0]   video_ctrl_apb_PRDATA;
  wire                video_ctrl_axi_ar_valid;
  wire       [31:0]   video_ctrl_axi_ar_payload_addr;
  wire       [7:0]    video_ctrl_axi_ar_payload_len;
  wire       [1:0]    video_ctrl_axi_ar_payload_burst;
  wire                video_ctrl_axi_r_ready;
  wire                peripheral_uart_ctrl_uart_tx;
  wire                peripheral_uart_ctrl_interrupt;
  wire                peripheral_uart_ctrl_apb_PREADY;
  wire       [31:0]   peripheral_uart_ctrl_apb_PRDATA;
  wire                peripheral_audio_ctrl_shdn;
  wire                peripheral_audio_ctrl_i2c_scl;
  wire                peripheral_audio_ctrl_apb_PREADY;
  wire       [31:0]   peripheral_audio_ctrl_apb_PRDATA;
  wire                peripheral_sdcard_ctrl_sdcard_clk;
  wire                peripheral_sdcard_ctrl_interrupt;
  wire                peripheral_sdcard_ctrl_apb_PREADY;
  wire       [31:0]   peripheral_sdcard_ctrl_apb_PRDATA;
  wire                peripheral_usb_ctrl_io_apb_ctrl_PREADY;
  wire       [31:0]   peripheral_usb_ctrl_io_apb_ctrl_PRDATA;
  wire                peripheral_usb_ctrl_io_apb_dma_PREADY;
  wire       [31:0]   peripheral_usb_ctrl_io_apb_dma_PRDATA;
  wire                peripheral_usb_ctrl_io_interrupt;
  wire                peripheral_usb_ctrl__zz_io_interrupt;
  wire                peripheral_apb_decoder_io_input_PREADY;
  wire       [31:0]   peripheral_apb_decoder_io_input_PRDATA;
  wire       [18:0]   peripheral_apb_decoder_io_output_PADDR;
  wire       [4:0]    peripheral_apb_decoder_io_output_PSEL;
  wire                peripheral_apb_decoder_io_output_PENABLE;
  wire                peripheral_apb_decoder_io_output_PWRITE;
  wire       [31:0]   peripheral_apb_decoder_io_output_PWDATA;
  wire                apb3Router_2_io_input_PREADY;
  wire       [31:0]   apb3Router_2_io_input_PRDATA;
  wire       [18:0]   apb3Router_2_io_outputs_0_PADDR;
  wire       [0:0]    apb3Router_2_io_outputs_0_PSEL;
  wire                apb3Router_2_io_outputs_0_PENABLE;
  wire                apb3Router_2_io_outputs_0_PWRITE;
  wire       [31:0]   apb3Router_2_io_outputs_0_PWDATA;
  wire       [18:0]   apb3Router_2_io_outputs_1_PADDR;
  wire       [0:0]    apb3Router_2_io_outputs_1_PSEL;
  wire                apb3Router_2_io_outputs_1_PENABLE;
  wire                apb3Router_2_io_outputs_1_PWRITE;
  wire       [31:0]   apb3Router_2_io_outputs_1_PWDATA;
  wire       [18:0]   apb3Router_2_io_outputs_2_PADDR;
  wire       [0:0]    apb3Router_2_io_outputs_2_PSEL;
  wire                apb3Router_2_io_outputs_2_PENABLE;
  wire                apb3Router_2_io_outputs_2_PWRITE;
  wire       [31:0]   apb3Router_2_io_outputs_2_PWDATA;
  wire       [18:0]   apb3Router_2_io_outputs_3_PADDR;
  wire       [0:0]    apb3Router_2_io_outputs_3_PSEL;
  wire                apb3Router_2_io_outputs_3_PENABLE;
  wire                apb3Router_2_io_outputs_3_PWRITE;
  wire       [31:0]   apb3Router_2_io_outputs_3_PWDATA;
  wire       [18:0]   apb3Router_2_io_outputs_4_PADDR;
  wire       [0:0]    apb3Router_2_io_outputs_4_PSEL;
  wire                apb3Router_2_io_outputs_4_PENABLE;
  wire                apb3Router_2_io_outputs_4_PWRITE;
  wire       [31:0]   apb3Router_2_io_outputs_4_PWDATA;
  wire                peripheral_apb_bridge_input_PREADY;
  wire       [31:0]   peripheral_apb_bridge_input_PRDATA;
  wire       [18:0]   peripheral_apb_bridge_output_PADDR;
  wire       [0:0]    peripheral_apb_bridge_output_PSEL;
  wire                peripheral_apb_bridge_output_PENABLE;
  wire                peripheral_apb_bridge_output_PWRITE;
  wire       [31:0]   peripheral_apb_bridge_output_PWDATA;
  wire                vexiiRiscv_1_FetchL1TileLinkPlugin_logic_down_a_valid;
  wire       [2:0]    vexiiRiscv_1_FetchL1TileLinkPlugin_logic_down_a_payload_opcode;
  wire       [2:0]    vexiiRiscv_1_FetchL1TileLinkPlugin_logic_down_a_payload_param;
  wire       [31:0]   vexiiRiscv_1_FetchL1TileLinkPlugin_logic_down_a_payload_address;
  wire       [2:0]    vexiiRiscv_1_FetchL1TileLinkPlugin_logic_down_a_payload_size;
  wire                vexiiRiscv_1_FetchL1TileLinkPlugin_logic_down_d_ready;
  wire                vexiiRiscv_1_LsuL1TileLinkPlugin_logic_down_a_valid;
  wire       [2:0]    vexiiRiscv_1_LsuL1TileLinkPlugin_logic_down_a_payload_opcode;
  wire       [2:0]    vexiiRiscv_1_LsuL1TileLinkPlugin_logic_down_a_payload_param;
  wire       [0:0]    vexiiRiscv_1_LsuL1TileLinkPlugin_logic_down_a_payload_source;
  wire       [31:0]   vexiiRiscv_1_LsuL1TileLinkPlugin_logic_down_a_payload_address;
  wire       [2:0]    vexiiRiscv_1_LsuL1TileLinkPlugin_logic_down_a_payload_size;
  wire       [7:0]    vexiiRiscv_1_LsuL1TileLinkPlugin_logic_down_a_payload_mask;
  wire       [63:0]   vexiiRiscv_1_LsuL1TileLinkPlugin_logic_down_a_payload_data;
  wire                vexiiRiscv_1_LsuL1TileLinkPlugin_logic_down_a_payload_corrupt;
  wire                vexiiRiscv_1_LsuL1TileLinkPlugin_logic_down_d_ready;
  wire                vexiiRiscv_1_LsuTileLinkPlugin_logic_bridge_down_a_valid;
  wire       [2:0]    vexiiRiscv_1_LsuTileLinkPlugin_logic_bridge_down_a_payload_opcode;
  wire       [2:0]    vexiiRiscv_1_LsuTileLinkPlugin_logic_bridge_down_a_payload_param;
  wire       [31:0]   vexiiRiscv_1_LsuTileLinkPlugin_logic_bridge_down_a_payload_address;
  wire       [1:0]    vexiiRiscv_1_LsuTileLinkPlugin_logic_bridge_down_a_payload_size;
  wire       [3:0]    vexiiRiscv_1_LsuTileLinkPlugin_logic_bridge_down_a_payload_mask;
  wire       [31:0]   vexiiRiscv_1_LsuTileLinkPlugin_logic_bridge_down_a_payload_data;
  wire                vexiiRiscv_1_LsuTileLinkPlugin_logic_bridge_down_a_payload_corrupt;
  wire                vexiiRiscv_1_LsuTileLinkPlugin_logic_bridge_down_d_ready;
  wire                arbiter_1_io_ups_0_a_ready;
  wire                arbiter_1_io_ups_0_d_valid;
  wire       [2:0]    arbiter_1_io_ups_0_d_payload_opcode;
  wire       [2:0]    arbiter_1_io_ups_0_d_payload_param;
  wire       [2:0]    arbiter_1_io_ups_0_d_payload_size;
  wire                arbiter_1_io_ups_0_d_payload_denied;
  wire       [63:0]   arbiter_1_io_ups_0_d_payload_data;
  wire                arbiter_1_io_ups_0_d_payload_corrupt;
  wire                arbiter_1_io_ups_1_a_ready;
  wire                arbiter_1_io_ups_1_d_valid;
  wire       [2:0]    arbiter_1_io_ups_1_d_payload_opcode;
  wire       [2:0]    arbiter_1_io_ups_1_d_payload_param;
  wire       [1:0]    arbiter_1_io_ups_1_d_payload_size;
  wire                arbiter_1_io_ups_1_d_payload_denied;
  wire       [63:0]   arbiter_1_io_ups_1_d_payload_data;
  wire                arbiter_1_io_ups_1_d_payload_corrupt;
  wire                arbiter_1_io_ups_2_a_ready;
  wire                arbiter_1_io_ups_2_d_valid;
  wire       [2:0]    arbiter_1_io_ups_2_d_payload_opcode;
  wire       [2:0]    arbiter_1_io_ups_2_d_payload_param;
  wire       [0:0]    arbiter_1_io_ups_2_d_payload_source;
  wire       [2:0]    arbiter_1_io_ups_2_d_payload_size;
  wire                arbiter_1_io_ups_2_d_payload_denied;
  wire       [63:0]   arbiter_1_io_ups_2_d_payload_data;
  wire                arbiter_1_io_ups_2_d_payload_corrupt;
  wire                arbiter_1_io_down_a_valid;
  wire       [2:0]    arbiter_1_io_down_a_payload_opcode;
  wire       [2:0]    arbiter_1_io_down_a_payload_param;
  wire       [2:0]    arbiter_1_io_down_a_payload_source;
  wire       [31:0]   arbiter_1_io_down_a_payload_address;
  wire       [2:0]    arbiter_1_io_down_a_payload_size;
  wire       [7:0]    arbiter_1_io_down_a_payload_mask;
  wire       [63:0]   arbiter_1_io_down_a_payload_data;
  wire                arbiter_1_io_down_a_payload_corrupt;
  wire                arbiter_1_io_down_d_ready;
  wire                ramBridge_logic_bridge_io_up_a_ready;
  wire                ramBridge_logic_bridge_io_up_d_valid;
  wire       [2:0]    ramBridge_logic_bridge_io_up_d_payload_opcode;
  wire       [2:0]    ramBridge_logic_bridge_io_up_d_payload_param;
  wire       [2:0]    ramBridge_logic_bridge_io_up_d_payload_source;
  wire       [2:0]    ramBridge_logic_bridge_io_up_d_payload_size;
  wire                ramBridge_logic_bridge_io_up_d_payload_denied;
  wire       [63:0]   ramBridge_logic_bridge_io_up_d_payload_data;
  wire                ramBridge_logic_bridge_io_up_d_payload_corrupt;
  wire                ramBridge_logic_bridge_io_down_ar_valid;
  wire       [26:0]   ramBridge_logic_bridge_io_down_ar_payload_addr;
  wire       [2:0]    ramBridge_logic_bridge_io_down_ar_payload_id;
  wire       [7:0]    ramBridge_logic_bridge_io_down_ar_payload_len;
  wire       [2:0]    ramBridge_logic_bridge_io_down_ar_payload_size;
  wire       [1:0]    ramBridge_logic_bridge_io_down_ar_payload_burst;
  wire                ramBridge_logic_bridge_io_down_aw_valid;
  wire       [26:0]   ramBridge_logic_bridge_io_down_aw_payload_addr;
  wire       [2:0]    ramBridge_logic_bridge_io_down_aw_payload_id;
  wire       [7:0]    ramBridge_logic_bridge_io_down_aw_payload_len;
  wire       [2:0]    ramBridge_logic_bridge_io_down_aw_payload_size;
  wire       [1:0]    ramBridge_logic_bridge_io_down_aw_payload_burst;
  wire                ramBridge_logic_bridge_io_down_aw_payload_allStrb;
  wire                ramBridge_logic_bridge_io_down_w_valid;
  wire       [63:0]   ramBridge_logic_bridge_io_down_w_payload_data;
  wire       [7:0]    ramBridge_logic_bridge_io_down_w_payload_strb;
  wire                ramBridge_logic_bridge_io_down_w_payload_last;
  wire                ramBridge_logic_bridge_io_down_r_ready;
  wire                ramBridge_logic_bridge_io_down_b_ready;
  wire                widthAdapter_2_io_up_a_ready;
  wire                widthAdapter_2_io_up_d_valid;
  wire       [2:0]    widthAdapter_2_io_up_d_payload_opcode;
  wire       [2:0]    widthAdapter_2_io_up_d_payload_param;
  wire       [1:0]    widthAdapter_2_io_up_d_payload_size;
  wire                widthAdapter_2_io_up_d_payload_denied;
  wire       [31:0]   widthAdapter_2_io_up_d_payload_data;
  wire                widthAdapter_2_io_up_d_payload_corrupt;
  wire                widthAdapter_2_io_down_a_valid;
  wire       [2:0]    widthAdapter_2_io_down_a_payload_opcode;
  wire       [2:0]    widthAdapter_2_io_down_a_payload_param;
  wire       [31:0]   widthAdapter_2_io_down_a_payload_address;
  wire       [1:0]    widthAdapter_2_io_down_a_payload_size;
  wire       [7:0]    widthAdapter_2_io_down_a_payload_mask;
  wire       [63:0]   widthAdapter_2_io_down_a_payload_data;
  wire                widthAdapter_2_io_down_a_payload_corrupt;
  wire                widthAdapter_2_io_down_d_ready;
  wire                streamArbiter_10_io_inputs_0_ready;
  wire                streamArbiter_10_io_inputs_1_ready;
  wire                streamArbiter_10_io_output_valid;
  wire       [26:0]   streamArbiter_10_io_output_payload_addr;
  wire       [2:0]    streamArbiter_10_io_output_payload_id;
  wire       [7:0]    streamArbiter_10_io_output_payload_len;
  wire       [2:0]    streamArbiter_10_io_output_payload_size;
  wire       [1:0]    streamArbiter_10_io_output_payload_burst;
  wire                streamArbiter_10_io_output_payload_allStrb;
  wire       [0:0]    streamArbiter_10_io_chosen;
  wire       [1:0]    streamArbiter_10_io_chosenOH;
  wire                ram_ddr_ctrl_arw_ready;
  wire                ram_ddr_ctrl_wready;
  wire                ram_ddr_ctrl_bvalid;
  wire       [2:0]    ram_ddr_ctrl_bid;
  wire       [1:0]    ram_ddr_ctrl_bresp;
  wire                ram_ddr_ctrl_rvalid;
  wire       [63:0]   ram_ddr_ctrl_rdata;
  wire       [2:0]    ram_ddr_ctrl_rid;
  wire       [1:0]    ram_ddr_ctrl_rresp;
  wire                ram_ddr_ctrl_rlast;
  wire                ram_ddr_ctrl_ddr_ck_p;
  wire                ram_ddr_ctrl_ddr_ck_n;
  wire                ram_ddr_ctrl_ddr_cke;
  wire                ram_ddr_ctrl_ddr_ras_n;
  wire                ram_ddr_ctrl_ddr_cas_n;
  wire                ram_ddr_ctrl_ddr_we_n;
  wire       [1:0]    ram_ddr_ctrl_ddr_ba;
  wire       [13:0]   ram_ddr_ctrl_ddr_a;
  wire       [1:0]    ram_ddr_ctrl_ddr_dm;
  wire                ram_axi_cc_io_input_arw_ready;
  wire                ram_axi_cc_io_input_w_ready;
  wire                ram_axi_cc_io_input_b_valid;
  wire       [2:0]    ram_axi_cc_io_input_b_payload_id;
  wire       [1:0]    ram_axi_cc_io_input_b_payload_resp;
  wire                ram_axi_cc_io_input_r_valid;
  wire       [63:0]   ram_axi_cc_io_input_r_payload_data;
  wire       [2:0]    ram_axi_cc_io_input_r_payload_id;
  wire       [1:0]    ram_axi_cc_io_input_r_payload_resp;
  wire                ram_axi_cc_io_input_r_payload_last;
  wire                ram_axi_cc_io_output_arw_valid;
  wire       [26:0]   ram_axi_cc_io_output_arw_payload_addr;
  wire       [2:0]    ram_axi_cc_io_output_arw_payload_id;
  wire       [7:0]    ram_axi_cc_io_output_arw_payload_len;
  wire       [2:0]    ram_axi_cc_io_output_arw_payload_size;
  wire       [1:0]    ram_axi_cc_io_output_arw_payload_burst;
  wire                ram_axi_cc_io_output_arw_payload_allStrb;
  wire                ram_axi_cc_io_output_arw_payload_write;
  wire                ram_axi_cc_io_output_w_valid;
  wire       [63:0]   ram_axi_cc_io_output_w_payload_data;
  wire       [7:0]    ram_axi_cc_io_output_w_payload_strb;
  wire                ram_axi_cc_io_output_w_payload_last;
  wire                ram_axi_cc_io_output_b_ready;
  wire                ram_axi_cc_io_output_r_ready;
  wire                decoder_2_io_up_a_ready;
  wire                decoder_2_io_up_d_valid;
  wire       [2:0]    decoder_2_io_up_d_payload_opcode;
  wire       [2:0]    decoder_2_io_up_d_payload_param;
  wire       [2:0]    decoder_2_io_up_d_payload_source;
  wire       [2:0]    decoder_2_io_up_d_payload_size;
  wire                decoder_2_io_up_d_payload_denied;
  wire       [63:0]   decoder_2_io_up_d_payload_data;
  wire                decoder_2_io_up_d_payload_corrupt;
  wire                decoder_2_io_downs_0_a_valid;
  wire       [2:0]    decoder_2_io_downs_0_a_payload_opcode;
  wire       [2:0]    decoder_2_io_downs_0_a_payload_param;
  wire       [2:0]    decoder_2_io_downs_0_a_payload_source;
  wire       [30:0]   decoder_2_io_downs_0_a_payload_address;
  wire       [2:0]    decoder_2_io_downs_0_a_payload_size;
  wire       [7:0]    decoder_2_io_downs_0_a_payload_mask;
  wire       [63:0]   decoder_2_io_downs_0_a_payload_data;
  wire                decoder_2_io_downs_0_a_payload_corrupt;
  wire                decoder_2_io_downs_0_d_ready;
  wire                decoder_2_io_downs_1_a_valid;
  wire       [2:0]    decoder_2_io_downs_1_a_payload_opcode;
  wire       [2:0]    decoder_2_io_downs_1_a_payload_param;
  wire       [2:0]    decoder_2_io_downs_1_a_payload_source;
  wire       [26:0]   decoder_2_io_downs_1_a_payload_address;
  wire       [2:0]    decoder_2_io_downs_1_a_payload_size;
  wire       [7:0]    decoder_2_io_downs_1_a_payload_mask;
  wire       [63:0]   decoder_2_io_downs_1_a_payload_data;
  wire                decoder_2_io_downs_1_a_payload_corrupt;
  wire                decoder_2_io_downs_1_d_ready;
  wire                toApb_logic_bridge_io_up_a_ready;
  wire                toApb_logic_bridge_io_up_d_valid;
  wire       [2:0]    toApb_logic_bridge_io_up_d_payload_opcode;
  wire       [2:0]    toApb_logic_bridge_io_up_d_payload_param;
  wire       [2:0]    toApb_logic_bridge_io_up_d_payload_source;
  wire       [2:0]    toApb_logic_bridge_io_up_d_payload_size;
  wire                toApb_logic_bridge_io_up_d_payload_denied;
  wire       [31:0]   toApb_logic_bridge_io_up_d_payload_data;
  wire                toApb_logic_bridge_io_up_d_payload_corrupt;
  wire       [26:0]   toApb_logic_bridge_io_down_PADDR;
  wire       [0:0]    toApb_logic_bridge_io_down_PSEL;
  wire                toApb_logic_bridge_io_down_PENABLE;
  wire                toApb_logic_bridge_io_down_PWRITE;
  wire       [31:0]   toApb_logic_bridge_io_down_PWDATA;
  wire                internalRam_thread_logic_io_up_a_ready;
  wire                internalRam_thread_logic_io_up_d_valid;
  wire       [2:0]    internalRam_thread_logic_io_up_d_payload_opcode;
  wire       [2:0]    internalRam_thread_logic_io_up_d_payload_param;
  wire       [2:0]    internalRam_thread_logic_io_up_d_payload_source;
  wire       [2:0]    internalRam_thread_logic_io_up_d_payload_size;
  wire                internalRam_thread_logic_io_up_d_payload_denied;
  wire       [31:0]   internalRam_thread_logic_io_up_d_payload_data;
  wire                internalRam_thread_logic_io_up_d_payload_corrupt;
  wire                widthAdapter_3_io_up_a_ready;
  wire                widthAdapter_3_io_up_d_valid;
  wire       [2:0]    widthAdapter_3_io_up_d_payload_opcode;
  wire       [2:0]    widthAdapter_3_io_up_d_payload_param;
  wire       [2:0]    widthAdapter_3_io_up_d_payload_source;
  wire       [2:0]    widthAdapter_3_io_up_d_payload_size;
  wire                widthAdapter_3_io_up_d_payload_denied;
  wire       [63:0]   widthAdapter_3_io_up_d_payload_data;
  wire                widthAdapter_3_io_up_d_payload_corrupt;
  wire                widthAdapter_3_io_down_a_valid;
  wire       [2:0]    widthAdapter_3_io_down_a_payload_opcode;
  wire       [2:0]    widthAdapter_3_io_down_a_payload_param;
  wire       [2:0]    widthAdapter_3_io_down_a_payload_source;
  wire       [30:0]   widthAdapter_3_io_down_a_payload_address;
  wire       [2:0]    widthAdapter_3_io_down_a_payload_size;
  wire       [3:0]    widthAdapter_3_io_down_a_payload_mask;
  wire       [31:0]   widthAdapter_3_io_down_a_payload_data;
  wire                widthAdapter_3_io_down_a_payload_corrupt;
  wire                widthAdapter_3_io_down_d_ready;
  wire                decoder_3_io_up_a_ready;
  wire                decoder_3_io_up_d_valid;
  wire       [2:0]    decoder_3_io_up_d_payload_opcode;
  wire       [2:0]    decoder_3_io_up_d_payload_param;
  wire       [2:0]    decoder_3_io_up_d_payload_source;
  wire       [2:0]    decoder_3_io_up_d_payload_size;
  wire                decoder_3_io_up_d_payload_denied;
  wire       [31:0]   decoder_3_io_up_d_payload_data;
  wire                decoder_3_io_up_d_payload_corrupt;
  wire                decoder_3_io_downs_0_a_valid;
  wire       [2:0]    decoder_3_io_downs_0_a_payload_opcode;
  wire       [2:0]    decoder_3_io_downs_0_a_payload_param;
  wire       [2:0]    decoder_3_io_downs_0_a_payload_source;
  wire       [26:0]   decoder_3_io_downs_0_a_payload_address;
  wire       [2:0]    decoder_3_io_downs_0_a_payload_size;
  wire       [3:0]    decoder_3_io_downs_0_a_payload_mask;
  wire       [31:0]   decoder_3_io_downs_0_a_payload_data;
  wire                decoder_3_io_downs_0_a_payload_corrupt;
  wire                decoder_3_io_downs_0_d_ready;
  wire                decoder_3_io_downs_1_a_valid;
  wire       [2:0]    decoder_3_io_downs_1_a_payload_opcode;
  wire       [2:0]    decoder_3_io_downs_1_a_payload_param;
  wire       [2:0]    decoder_3_io_downs_1_a_payload_source;
  wire       [13:0]   decoder_3_io_downs_1_a_payload_address;
  wire       [2:0]    decoder_3_io_downs_1_a_payload_size;
  wire       [3:0]    decoder_3_io_downs_1_a_payload_mask;
  wire       [31:0]   decoder_3_io_downs_1_a_payload_data;
  wire                decoder_3_io_downs_1_a_payload_corrupt;
  wire                decoder_3_io_downs_1_d_ready;
  wire                toApb_down_decoder_io_input_PREADY;
  wire       [31:0]   toApb_down_decoder_io_input_PRDATA;
  wire                toApb_down_decoder_io_input_PSLVERROR;
  wire       [26:0]   toApb_down_decoder_io_output_PADDR;
  wire       [3:0]    toApb_down_decoder_io_output_PSEL;
  wire                toApb_down_decoder_io_output_PENABLE;
  wire                toApb_down_decoder_io_output_PWRITE;
  wire       [31:0]   toApb_down_decoder_io_output_PWDATA;
  wire                apb3Router_3_io_input_PREADY;
  wire       [31:0]   apb3Router_3_io_input_PRDATA;
  wire                apb3Router_3_io_input_PSLVERROR;
  wire       [26:0]   apb3Router_3_io_outputs_0_PADDR;
  wire       [0:0]    apb3Router_3_io_outputs_0_PSEL;
  wire                apb3Router_3_io_outputs_0_PENABLE;
  wire                apb3Router_3_io_outputs_0_PWRITE;
  wire       [31:0]   apb3Router_3_io_outputs_0_PWDATA;
  wire       [26:0]   apb3Router_3_io_outputs_1_PADDR;
  wire       [0:0]    apb3Router_3_io_outputs_1_PSEL;
  wire                apb3Router_3_io_outputs_1_PENABLE;
  wire                apb3Router_3_io_outputs_1_PWRITE;
  wire       [31:0]   apb3Router_3_io_outputs_1_PWDATA;
  wire       [26:0]   apb3Router_3_io_outputs_2_PADDR;
  wire       [0:0]    apb3Router_3_io_outputs_2_PSEL;
  wire                apb3Router_3_io_outputs_2_PENABLE;
  wire                apb3Router_3_io_outputs_2_PWRITE;
  wire       [31:0]   apb3Router_3_io_outputs_2_PWDATA;
  wire       [26:0]   apb3Router_3_io_outputs_3_PADDR;
  wire       [0:0]    apb3Router_3_io_outputs_3_PSEL;
  wire                apb3Router_3_io_outputs_3_PENABLE;
  wire                apb3Router_3_io_outputs_3_PWRITE;
  wire       [31:0]   apb3Router_3_io_outputs_3_PWDATA;
  wire       [18:0]   peripheral_apb_PADDR;
  wire       [0:0]    peripheral_apb_PSEL;
  wire                peripheral_apb_PENABLE;
  wire                peripheral_apb_PREADY;
  wire                peripheral_apb_PWRITE;
  wire       [31:0]   peripheral_apb_PWDATA;
  wire       [31:0]   peripheral_apb_PRDATA;
  (* async_reg = "true" *) reg                 usb_interrupt;
  wire       [0:0]    plic_gateways_0_priority;
  reg                 plic_gateways_0_ip;
  reg                 plic_gateways_0_waitCompletion;
  wire                when_PlicGateway_l21;
  wire       [0:0]    plic_gateways_1_priority;
  reg                 plic_gateways_1_ip;
  reg                 plic_gateways_1_waitCompletion;
  wire                when_PlicGateway_l21_1;
  wire       [0:0]    plic_gateways_2_priority;
  reg                 plic_gateways_2_ip;
  reg                 plic_gateways_2_waitCompletion;
  wire                when_PlicGateway_l21_2;
  wire                plic_target_ie_0;
  wire                plic_target_ie_1;
  wire                plic_target_ie_2;
  wire       [0:0]    plic_target_threshold;
  wire       [0:0]    plic_target_requests_0_priority;
  wire       [1:0]    plic_target_requests_0_id;
  wire                plic_target_requests_0_valid;
  wire       [0:0]    plic_target_requests_1_priority;
  wire       [1:0]    plic_target_requests_1_id;
  wire                plic_target_requests_1_valid;
  wire       [0:0]    plic_target_requests_2_priority;
  wire       [1:0]    plic_target_requests_2_id;
  wire                plic_target_requests_2_valid;
  wire       [0:0]    plic_target_requests_3_priority;
  wire       [1:0]    plic_target_requests_3_id;
  wire                plic_target_requests_3_valid;
  wire                _zz_plic_target_bestRequest_id;
  wire       [0:0]    _zz_plic_target_bestRequest_priority;
  wire                _zz_plic_target_bestRequest_valid;
  wire                _zz_plic_target_bestRequest_id_1;
  wire       [0:0]    _zz_plic_target_bestRequest_priority_1;
  wire                _zz_plic_target_bestRequest_valid_1;
  wire                _zz_plic_target_bestRequest_priority_2;
  reg        [0:0]    plic_target_bestRequest_priority;
  reg        [1:0]    plic_target_bestRequest_id;
  reg                 plic_target_bestRequest_valid;
  wire                plic_target_iep;
  wire       [1:0]    plic_target_claim;
  wire       [25:0]   plic_apb_PADDR;
  wire       [0:0]    plic_apb_PSEL;
  wire                plic_apb_PENABLE;
  reg                 plic_apb_PREADY;
  wire                plic_apb_PWRITE;
  wire       [31:0]   plic_apb_PWDATA;
  reg        [31:0]   plic_apb_PRDATA;
  wire                _zz_1;
  wire                _zz_2;
  wire                _zz_3;
  wire                _zz_4;
  reg        [0:0]    _zz_plic_gateways_0_priority;
  reg        [0:0]    _zz_plic_gateways_1_priority;
  reg        [0:0]    _zz_plic_gateways_2_priority;
  reg                 plic_claim_valid;
  reg        [1:0]    plic_claim_payload;
  reg                 plic_completion_valid;
  reg        [1:0]    plic_completion_payload;
  reg                 plic_coherencyStall_willIncrement;
  wire                plic_coherencyStall_willClear;
  reg        [0:0]    plic_coherencyStall_valueNext;
  reg        [0:0]    plic_coherencyStall_value;
  wire                plic_coherencyStall_willOverflowIfInc;
  wire                plic_coherencyStall_willOverflow;
  wire                when_PlicMapper_l122;
  reg        [0:0]    _zz_plic_target_threshold;
  reg                 plic_targetMapping_0_targetCompletion_valid;
  wire       [1:0]    plic_targetMapping_0_targetCompletion_payload;
  reg                 _zz_plic_target_ie_0;
  reg                 _zz_plic_target_ie_1;
  reg                 _zz_plic_target_ie_2;
  wire                when_Apb3SlaveFactory_l81;
  wire                _zz_FetchL1TileLinkPlugin_logic_down_a_ready;
  wire       [2:0]    _zz_io_ups_0_a_payload_opcode;
  wire       [2:0]    _zz_FetchL1TileLinkPlugin_logic_down_d_payload_opcode;
  wire       [2:0]    _zz_io_ups_0_a_payload_opcode_1;
  reg                 _zz_io_ups_0_d_ready;
  wire       [2:0]    _zz_FetchL1TileLinkPlugin_logic_down_d_payload_opcode_1;
  wire                _zz_5;
  wire                _zz_6;
  wire       [2:0]    _zz_io_ups_0_a_payload_opcode_2;
  reg                 _zz_FetchL1TileLinkPlugin_logic_down_a_ready_1;
  reg        [2:0]    _zz_io_ups_0_a_payload_opcode_3;
  reg        [2:0]    _zz_io_ups_0_a_payload_param;
  reg        [31:0]   _zz_io_ups_0_a_payload_address;
  reg        [2:0]    _zz_io_ups_0_a_payload_size;
  wire                _zz_io_ups_0_a_valid;
  wire       [2:0]    _zz_io_ups_0_a_payload_opcode_4;
  reg                 _zz_io_ups_0_a_valid_1;
  reg        [2:0]    _zz_io_ups_0_a_payload_opcode_5;
  reg        [2:0]    _zz_io_ups_0_a_payload_param_1;
  reg        [31:0]   _zz_io_ups_0_a_payload_address_1;
  reg        [2:0]    _zz_io_ups_0_a_payload_size_1;
  wire                _zz_when_Stream_l393;
  wire       [2:0]    _zz_FetchL1TileLinkPlugin_logic_down_d_payload_opcode_2;
  reg                 _zz_when_Stream_l393_1;
  reg        [2:0]    _zz_FetchL1TileLinkPlugin_logic_down_d_payload_opcode_3;
  reg        [2:0]    _zz_FetchL1TileLinkPlugin_logic_down_d_payload_param;
  reg        [2:0]    _zz_FetchL1TileLinkPlugin_logic_down_d_payload_size;
  reg                 _zz_FetchL1TileLinkPlugin_logic_down_d_payload_denied;
  reg        [63:0]   _zz_FetchL1TileLinkPlugin_logic_down_d_payload_data;
  reg                 _zz_FetchL1TileLinkPlugin_logic_down_d_payload_corrupt;
  wire                when_Stream_l393;
  wire                _zz_LsuTileLinkPlugin_logic_bridge_down_a_ready;
  wire       [2:0]    _zz_io_up_a_payload_opcode;
  wire       [2:0]    _zz_LsuTileLinkPlugin_logic_bridge_down_d_payload_opcode;
  wire       [2:0]    _zz_io_up_a_payload_opcode_1;
  reg                 _zz_io_up_d_ready;
  wire       [2:0]    _zz_LsuTileLinkPlugin_logic_bridge_down_d_payload_opcode_1;
  wire                _zz_io_up_a_valid;
  wire       [2:0]    _zz_io_up_a_payload_opcode_2;
  reg                 _zz_LsuTileLinkPlugin_logic_bridge_down_a_ready_1;
  reg        [2:0]    _zz_io_up_a_payload_opcode_3;
  reg        [2:0]    _zz_io_up_a_payload_param;
  reg        [31:0]   _zz_io_up_a_payload_address;
  reg        [1:0]    _zz_io_up_a_payload_size;
  reg        [3:0]    _zz_io_up_a_payload_mask;
  reg        [31:0]   _zz_io_up_a_payload_data;
  reg                 _zz_io_up_a_payload_corrupt;
  wire                _zz_when_Stream_l393_2;
  wire       [2:0]    _zz_LsuTileLinkPlugin_logic_bridge_down_d_payload_opcode_2;
  (* keep , syn_keep *) reg                 _zz_when_Stream_l393_3 /* synthesis syn_keep = 1 */ ;
  (* keep , syn_keep *) reg        [2:0]    _zz_LsuTileLinkPlugin_logic_bridge_down_d_payload_opcode_3 /* synthesis syn_keep = 1 */ ;
  (* keep , syn_keep *) reg        [2:0]    _zz_LsuTileLinkPlugin_logic_bridge_down_d_payload_param /* synthesis syn_keep = 1 */ ;
  (* keep , syn_keep *) reg        [1:0]    _zz_LsuTileLinkPlugin_logic_bridge_down_d_payload_size /* synthesis syn_keep = 1 */ ;
  (* keep , syn_keep *) reg                 _zz_LsuTileLinkPlugin_logic_bridge_down_d_payload_denied /* synthesis syn_keep = 1 */ ;
  (* keep , syn_keep *) reg        [31:0]   _zz_LsuTileLinkPlugin_logic_bridge_down_d_payload_data /* synthesis syn_keep = 1 */ ;
  (* keep , syn_keep *) reg                 _zz_LsuTileLinkPlugin_logic_bridge_down_d_payload_corrupt /* synthesis syn_keep = 1 */ ;
  wire                when_Stream_l393_1;
  wire                _zz_LsuL1TileLinkPlugin_logic_down_a_ready;
  wire       [2:0]    _zz_io_ups_2_a_payload_opcode;
  wire       [2:0]    _zz_LsuL1TileLinkPlugin_logic_down_d_payload_opcode;
  wire       [2:0]    _zz_io_ups_2_a_payload_opcode_1;
  reg                 _zz_io_ups_2_d_ready;
  wire       [2:0]    _zz_LsuL1TileLinkPlugin_logic_down_d_payload_opcode_1;
  wire                _zz_io_ups_2_a_valid;
  wire       [2:0]    _zz_io_ups_2_a_payload_opcode_2;
  reg                 _zz_LsuL1TileLinkPlugin_logic_down_a_ready_1;
  reg        [2:0]    _zz_io_ups_2_a_payload_opcode_3;
  reg        [2:0]    _zz_io_ups_2_a_payload_param;
  reg        [0:0]    _zz_io_ups_2_a_payload_source;
  reg        [31:0]   _zz_io_ups_2_a_payload_address;
  reg        [2:0]    _zz_io_ups_2_a_payload_size;
  reg        [7:0]    _zz_io_ups_2_a_payload_mask;
  reg        [63:0]   _zz_io_ups_2_a_payload_data;
  reg                 _zz_io_ups_2_a_payload_corrupt;
  wire                _zz_when_Stream_l393_4;
  wire       [2:0]    _zz_LsuL1TileLinkPlugin_logic_down_d_payload_opcode_2;
  (* keep , syn_keep *) reg                 _zz_when_Stream_l393_5 /* synthesis syn_keep = 1 */ ;
  (* keep , syn_keep *) reg        [2:0]    _zz_LsuL1TileLinkPlugin_logic_down_d_payload_opcode_3 /* synthesis syn_keep = 1 */ ;
  (* keep , syn_keep *) reg        [2:0]    _zz_LsuL1TileLinkPlugin_logic_down_d_payload_param /* synthesis syn_keep = 1 */ ;
  (* keep , syn_keep *) reg        [0:0]    _zz_LsuL1TileLinkPlugin_logic_down_d_payload_source /* synthesis syn_keep = 1 */ ;
  (* keep , syn_keep *) reg        [2:0]    _zz_LsuL1TileLinkPlugin_logic_down_d_payload_size /* synthesis syn_keep = 1 */ ;
  (* keep , syn_keep *) reg                 _zz_LsuL1TileLinkPlugin_logic_down_d_payload_denied /* synthesis syn_keep = 1 */ ;
  (* keep , syn_keep *) reg        [63:0]   _zz_LsuL1TileLinkPlugin_logic_down_d_payload_data /* synthesis syn_keep = 1 */ ;
  (* keep , syn_keep *) reg                 _zz_LsuL1TileLinkPlugin_logic_down_d_payload_corrupt /* synthesis syn_keep = 1 */ ;
  wire                when_Stream_l393_2;
  wire       [2:0]    _zz_io_up_a_payload_opcode_4;
  wire       [2:0]    _zz_io_down_d_payload_opcode;
  wire       [2:0]    _zz_io_ups_0_a_payload_opcode_6;
  wire       [2:0]    _zz_FetchL1TileLinkPlugin_logic_down_d_payload_opcode_4;
  wire       [2:0]    _zz_io_ups_1_a_payload_opcode;
  wire       [2:0]    _zz_io_down_d_payload_opcode_1;
  wire       [2:0]    _zz_io_ups_2_a_payload_opcode_4;
  wire       [2:0]    _zz_LsuL1TileLinkPlugin_logic_down_d_payload_opcode_4;
  wire       [2:0]    _zz_io_up_a_payload_opcode_5;
  wire       [2:0]    _zz_io_down_d_payload_opcode_2;
  wire       [2:0]    _zz_io_up_a_payload_opcode_6;
  wire       [2:0]    _zz_io_down_d_payload_opcode_3;
  wire                ramBridge_up_bus_a_valid;
  wire                ramBridge_up_bus_a_ready;
  wire       [2:0]    ramBridge_up_bus_a_payload_opcode;
  wire       [2:0]    ramBridge_up_bus_a_payload_param;
  wire       [2:0]    ramBridge_up_bus_a_payload_source;
  wire       [26:0]   ramBridge_up_bus_a_payload_address;
  wire       [2:0]    ramBridge_up_bus_a_payload_size;
  wire       [7:0]    ramBridge_up_bus_a_payload_mask;
  wire       [63:0]   ramBridge_up_bus_a_payload_data;
  wire                ramBridge_up_bus_a_payload_corrupt;
  wire                ramBridge_up_bus_d_valid;
  wire                ramBridge_up_bus_d_ready;
  wire       [2:0]    ramBridge_up_bus_d_payload_opcode;
  wire       [2:0]    ramBridge_up_bus_d_payload_param;
  wire       [2:0]    ramBridge_up_bus_d_payload_source;
  wire       [2:0]    ramBridge_up_bus_d_payload_size;
  wire                ramBridge_up_bus_d_payload_denied;
  wire       [63:0]   ramBridge_up_bus_d_payload_data;
  wire                ramBridge_up_bus_d_payload_corrupt;
  wire       [2:0]    _zz_ramBridge_up_bus_a_payload_opcode;
  wire       [2:0]    _zz_io_downs_1_d_payload_opcode;
  wire       [2:0]    _zz_io_ups_0_a_payload_opcode_7;
  wire       [2:0]    _zz_FetchL1TileLinkPlugin_logic_down_d_payload_opcode_5;
  wire       [2:0]    _zz_io_up_a_payload_opcode_7;
  wire       [2:0]    _zz_LsuTileLinkPlugin_logic_bridge_down_d_payload_opcode_4;
  wire       [2:0]    _zz_io_ups_2_a_payload_opcode_5;
  wire       [2:0]    _zz_LsuL1TileLinkPlugin_logic_down_d_payload_opcode_5;
  wire                ramBridge_down_aw_valid;
  wire                ramBridge_down_aw_ready;
  wire       [26:0]   ramBridge_down_aw_payload_addr;
  wire       [2:0]    ramBridge_down_aw_payload_id;
  wire       [7:0]    ramBridge_down_aw_payload_len;
  wire       [2:0]    ramBridge_down_aw_payload_size;
  wire       [1:0]    ramBridge_down_aw_payload_burst;
  wire                ramBridge_down_aw_payload_allStrb;
  wire                ramBridge_down_w_valid;
  wire                ramBridge_down_w_ready;
  wire       [63:0]   ramBridge_down_w_payload_data;
  wire       [7:0]    ramBridge_down_w_payload_strb;
  wire                ramBridge_down_w_payload_last;
  wire                ramBridge_down_b_valid;
  wire                ramBridge_down_b_ready;
  wire       [2:0]    ramBridge_down_b_payload_id;
  wire       [1:0]    ramBridge_down_b_payload_resp;
  wire                ramBridge_down_ar_valid;
  wire                ramBridge_down_ar_ready;
  wire       [26:0]   ramBridge_down_ar_payload_addr;
  wire       [2:0]    ramBridge_down_ar_payload_id;
  wire       [7:0]    ramBridge_down_ar_payload_len;
  wire       [2:0]    ramBridge_down_ar_payload_size;
  wire       [1:0]    ramBridge_down_ar_payload_burst;
  wire                ramBridge_down_r_valid;
  wire                ramBridge_down_r_ready;
  wire       [63:0]   ramBridge_down_r_payload_data;
  wire       [2:0]    ramBridge_down_r_payload_id;
  wire       [1:0]    ramBridge_down_r_payload_resp;
  wire                ramBridge_down_r_payload_last;
  wire                toApb_up_bus_a_valid;
  wire                toApb_up_bus_a_ready;
  wire       [2:0]    toApb_up_bus_a_payload_opcode;
  wire       [2:0]    toApb_up_bus_a_payload_param;
  wire       [2:0]    toApb_up_bus_a_payload_source;
  wire       [26:0]   toApb_up_bus_a_payload_address;
  wire       [2:0]    toApb_up_bus_a_payload_size;
  wire       [3:0]    toApb_up_bus_a_payload_mask;
  wire       [31:0]   toApb_up_bus_a_payload_data;
  wire                toApb_up_bus_a_payload_corrupt;
  wire                toApb_up_bus_d_valid;
  wire                toApb_up_bus_d_ready;
  wire       [2:0]    toApb_up_bus_d_payload_opcode;
  wire       [2:0]    toApb_up_bus_d_payload_param;
  wire       [2:0]    toApb_up_bus_d_payload_source;
  wire       [2:0]    toApb_up_bus_d_payload_size;
  wire                toApb_up_bus_d_payload_denied;
  wire       [31:0]   toApb_up_bus_d_payload_data;
  wire                toApb_up_bus_d_payload_corrupt;
  wire       [2:0]    _zz_toApb_up_bus_a_payload_opcode;
  wire       [2:0]    _zz_io_downs_0_d_payload_opcode;
  wire                internalRam_up_bus_a_valid;
  wire                internalRam_up_bus_a_ready;
  wire       [2:0]    internalRam_up_bus_a_payload_opcode;
  wire       [2:0]    internalRam_up_bus_a_payload_param;
  wire       [2:0]    internalRam_up_bus_a_payload_source;
  wire       [13:0]   internalRam_up_bus_a_payload_address;
  wire       [2:0]    internalRam_up_bus_a_payload_size;
  wire       [3:0]    internalRam_up_bus_a_payload_mask;
  wire       [31:0]   internalRam_up_bus_a_payload_data;
  wire                internalRam_up_bus_a_payload_corrupt;
  wire                internalRam_up_bus_d_valid;
  wire                internalRam_up_bus_d_ready;
  wire       [2:0]    internalRam_up_bus_d_payload_opcode;
  wire       [2:0]    internalRam_up_bus_d_payload_param;
  wire       [2:0]    internalRam_up_bus_d_payload_source;
  wire       [2:0]    internalRam_up_bus_d_payload_size;
  wire                internalRam_up_bus_d_payload_denied;
  wire       [31:0]   internalRam_up_bus_d_payload_data;
  wire                internalRam_up_bus_d_payload_corrupt;
  wire       [2:0]    _zz_internalRam_up_bus_a_payload_opcode;
  wire       [2:0]    _zz_io_downs_1_d_payload_opcode_1;
  wire                ram_axi_arw_valid;
  wire                ram_axi_arw_ready;
  wire       [26:0]   ram_axi_arw_payload_addr;
  wire       [2:0]    ram_axi_arw_payload_id;
  wire       [7:0]    ram_axi_arw_payload_len;
  wire       [2:0]    ram_axi_arw_payload_size;
  wire       [1:0]    ram_axi_arw_payload_burst;
  wire                ram_axi_arw_payload_allStrb;
  wire                ram_axi_arw_payload_write;
  wire                ram_axi_w_valid;
  wire                ram_axi_w_ready;
  wire       [63:0]   ram_axi_w_payload_data;
  wire       [7:0]    ram_axi_w_payload_strb;
  wire                ram_axi_w_payload_last;
  wire                ram_axi_b_valid;
  wire                ram_axi_b_ready;
  wire       [2:0]    ram_axi_b_payload_id;
  wire       [1:0]    ram_axi_b_payload_resp;
  wire                ram_axi_r_valid;
  wire                ram_axi_r_ready;
  wire       [63:0]   ram_axi_r_payload_data;
  wire       [2:0]    ram_axi_r_payload_id;
  wire       [1:0]    ram_axi_r_payload_resp;
  wire                ram_axi_r_payload_last;
  wire       [2:0]    _zz_io_up_a_payload_opcode_8;
  wire       [2:0]    _zz_io_downs_0_d_payload_opcode_1;
  wire       [2:0]    _zz_ramBridge_up_bus_a_payload_opcode_1;
  wire       [2:0]    _zz_io_downs_1_d_payload_opcode_2;
  wire       [26:0]   toApb_down_PADDR;
  wire       [0:0]    toApb_down_PSEL;
  wire                toApb_down_PENABLE;
  wire                toApb_down_PREADY;
  wire                toApb_down_PWRITE;
  wire       [31:0]   toApb_down_PWDATA;
  wire       [31:0]   toApb_down_PRDATA;
  wire                toApb_down_PSLVERROR;
  wire       [2:0]    _zz_toApb_up_bus_a_payload_opcode_1;
  wire       [2:0]    _zz_io_downs_0_d_payload_opcode_2;
  wire       [2:0]    _zz_internalRam_up_bus_a_payload_opcode_1;
  wire       [2:0]    _zz_io_downs_1_d_payload_opcode_3;
  `ifndef SYNTHESIS
  reg [127:0] _zz_io_ups_0_a_payload_opcode_string;
  reg [119:0] _zz_FetchL1TileLinkPlugin_logic_down_d_payload_opcode_string;
  reg [127:0] _zz_io_ups_0_a_payload_opcode_1_string;
  reg [119:0] _zz_FetchL1TileLinkPlugin_logic_down_d_payload_opcode_1_string;
  reg [127:0] _zz_io_ups_0_a_payload_opcode_2_string;
  reg [127:0] _zz_io_ups_0_a_payload_opcode_3_string;
  reg [127:0] _zz_io_ups_0_a_payload_opcode_4_string;
  reg [127:0] _zz_io_ups_0_a_payload_opcode_5_string;
  reg [119:0] _zz_FetchL1TileLinkPlugin_logic_down_d_payload_opcode_2_string;
  reg [119:0] _zz_FetchL1TileLinkPlugin_logic_down_d_payload_opcode_3_string;
  reg [127:0] _zz_io_up_a_payload_opcode_string;
  reg [119:0] _zz_LsuTileLinkPlugin_logic_bridge_down_d_payload_opcode_string;
  reg [127:0] _zz_io_up_a_payload_opcode_1_string;
  reg [119:0] _zz_LsuTileLinkPlugin_logic_bridge_down_d_payload_opcode_1_string;
  reg [127:0] _zz_io_up_a_payload_opcode_2_string;
  reg [127:0] _zz_io_up_a_payload_opcode_3_string;
  reg [119:0] _zz_LsuTileLinkPlugin_logic_bridge_down_d_payload_opcode_2_string;
  reg [119:0] _zz_LsuTileLinkPlugin_logic_bridge_down_d_payload_opcode_3_string;
  reg [127:0] _zz_io_ups_2_a_payload_opcode_string;
  reg [119:0] _zz_LsuL1TileLinkPlugin_logic_down_d_payload_opcode_string;
  reg [127:0] _zz_io_ups_2_a_payload_opcode_1_string;
  reg [119:0] _zz_LsuL1TileLinkPlugin_logic_down_d_payload_opcode_1_string;
  reg [127:0] _zz_io_ups_2_a_payload_opcode_2_string;
  reg [127:0] _zz_io_ups_2_a_payload_opcode_3_string;
  reg [119:0] _zz_LsuL1TileLinkPlugin_logic_down_d_payload_opcode_2_string;
  reg [119:0] _zz_LsuL1TileLinkPlugin_logic_down_d_payload_opcode_3_string;
  reg [127:0] _zz_io_up_a_payload_opcode_4_string;
  reg [119:0] _zz_io_down_d_payload_opcode_string;
  reg [127:0] _zz_io_ups_0_a_payload_opcode_6_string;
  reg [119:0] _zz_FetchL1TileLinkPlugin_logic_down_d_payload_opcode_4_string;
  reg [127:0] _zz_io_ups_1_a_payload_opcode_string;
  reg [119:0] _zz_io_down_d_payload_opcode_1_string;
  reg [127:0] _zz_io_ups_2_a_payload_opcode_4_string;
  reg [119:0] _zz_LsuL1TileLinkPlugin_logic_down_d_payload_opcode_4_string;
  reg [127:0] _zz_io_up_a_payload_opcode_5_string;
  reg [119:0] _zz_io_down_d_payload_opcode_2_string;
  reg [127:0] _zz_io_up_a_payload_opcode_6_string;
  reg [119:0] _zz_io_down_d_payload_opcode_3_string;
  reg [127:0] ramBridge_up_bus_a_payload_opcode_string;
  reg [119:0] ramBridge_up_bus_d_payload_opcode_string;
  reg [127:0] _zz_ramBridge_up_bus_a_payload_opcode_string;
  reg [119:0] _zz_io_downs_1_d_payload_opcode_string;
  reg [127:0] _zz_io_ups_0_a_payload_opcode_7_string;
  reg [119:0] _zz_FetchL1TileLinkPlugin_logic_down_d_payload_opcode_5_string;
  reg [127:0] _zz_io_up_a_payload_opcode_7_string;
  reg [119:0] _zz_LsuTileLinkPlugin_logic_bridge_down_d_payload_opcode_4_string;
  reg [127:0] _zz_io_ups_2_a_payload_opcode_5_string;
  reg [119:0] _zz_LsuL1TileLinkPlugin_logic_down_d_payload_opcode_5_string;
  reg [127:0] toApb_up_bus_a_payload_opcode_string;
  reg [119:0] toApb_up_bus_d_payload_opcode_string;
  reg [127:0] _zz_toApb_up_bus_a_payload_opcode_string;
  reg [119:0] _zz_io_downs_0_d_payload_opcode_string;
  reg [127:0] internalRam_up_bus_a_payload_opcode_string;
  reg [119:0] internalRam_up_bus_d_payload_opcode_string;
  reg [127:0] _zz_internalRam_up_bus_a_payload_opcode_string;
  reg [119:0] _zz_io_downs_1_d_payload_opcode_1_string;
  reg [127:0] _zz_io_up_a_payload_opcode_8_string;
  reg [119:0] _zz_io_downs_0_d_payload_opcode_1_string;
  reg [127:0] _zz_ramBridge_up_bus_a_payload_opcode_1_string;
  reg [119:0] _zz_io_downs_1_d_payload_opcode_2_string;
  reg [127:0] _zz_toApb_up_bus_a_payload_opcode_1_string;
  reg [119:0] _zz_io_downs_0_d_payload_opcode_2_string;
  reg [127:0] _zz_internalRam_up_bus_a_payload_opcode_1_string;
  reg [119:0] _zz_io_downs_1_d_payload_opcode_3_string;
  `endif


  BoardController board_ctrl (
    .nreset_in        (io_nreset                             ), //i
    .clk_in           (io_clk_in                             ), //i
    .plla_i2c_scl     (board_ctrl_plla_i2c_scl               ), //o
    .plla_i2c_sda     (io_plla_i2c_sda                       ), //~
    .plla_clk0        (io_plla_clk0                          ), //i
    .plla_clk1        (io_plla_clk1                          ), //i
    .plla_clk2        (io_plla_clk2                          ), //i
    .pllb_i2c_scl     (board_ctrl_pllb_i2c_scl               ), //o
    .pllb_i2c_sda     (io_pllb_i2c_sda                       ), //~
    .pllb_clk0        (io_pllb_clk0                          ), //i
    .pllb_clk1        (io_pllb_clk1                          ), //i
    .pllb_clk2        (io_pllb_clk2                          ), //i
    .reset_cpu        (board_ctrl_reset_cpu                  ), //o
    .reset_ram        (board_ctrl_reset_ram                  ), //o
    .reset_peripheral (board_ctrl_reset_peripheral           ), //o
    .clk_cpu          (board_ctrl_clk_cpu                    ), //o
    .clk_ram          (board_ctrl_clk_ram                    ), //o
    .clk_ram_bus      (board_ctrl_clk_ram_bus                ), //o
    .clk_peripheral   (board_ctrl_clk_peripheral             ), //o
    .utime            (board_ctrl_utime[63:0]                ), //o
    .timer_interrupt  (board_ctrl_timer_interrupt            ), //o
    .video_mode       (video_ctrl_video_mode_out[1:0]        ), //i
    .clk_tmds_pixel   (board_ctrl_clk_tmds_pixel             ), //o
    .clk_tmds_x5      (board_ctrl_clk_tmds_x5                ), //o
    .leds             (board_ctrl_leds[2:0]                  ), //o
    .keys             (io_keys[1:0]                          ), //i
    .apb_PADDR        (board_ctrl_apb_PADDR[4:0]             ), //i
    .apb_PSEL         (apb3Router_3_io_outputs_1_PSEL        ), //i
    .apb_PENABLE      (apb3Router_3_io_outputs_1_PENABLE     ), //i
    .apb_PREADY       (board_ctrl_apb_PREADY                 ), //o
    .apb_PWRITE       (apb3Router_3_io_outputs_1_PWRITE      ), //i
    .apb_PWDATA       (apb3Router_3_io_outputs_1_PWDATA[31:0]), //i
    .apb_PRDATA       (board_ctrl_apb_PRDATA[31:0]           )  //o
  );
  VideoController video_ctrl (
    .clk                  (board_ctrl_clk_cpu                    ), //i
    .reset                (board_ctrl_reset_cpu                  ), //i
    .video_mode_out       (video_ctrl_video_mode_out[1:0]        ), //o
    .tmds_pixel_clk       (board_ctrl_clk_tmds_pixel             ), //i
    .tmds_x5_clk          (board_ctrl_clk_tmds_x5                ), //i
    .dvi_tmds0p           (video_ctrl_dvi_tmds0p                 ), //o
    .dvi_tmds0m           (video_ctrl_dvi_tmds0m                 ), //o
    .dvi_tmds1p           (video_ctrl_dvi_tmds1p                 ), //o
    .dvi_tmds1m           (video_ctrl_dvi_tmds1m                 ), //o
    .dvi_tmds2p           (video_ctrl_dvi_tmds2p                 ), //o
    .dvi_tmds2m           (video_ctrl_dvi_tmds2m                 ), //o
    .dvi_tmdsCp           (video_ctrl_dvi_tmdsCp                 ), //o
    .dvi_tmdsCm           (video_ctrl_dvi_tmdsCm                 ), //o
    .apb_PADDR            (video_ctrl_apb_PADDR[4:0]             ), //i
    .apb_PSEL             (apb3Router_3_io_outputs_2_PSEL        ), //i
    .apb_PENABLE          (apb3Router_3_io_outputs_2_PENABLE     ), //i
    .apb_PREADY           (video_ctrl_apb_PREADY                 ), //o
    .apb_PWRITE           (apb3Router_3_io_outputs_2_PWRITE      ), //i
    .apb_PWDATA           (apb3Router_3_io_outputs_2_PWDATA[31:0]), //i
    .apb_PRDATA           (video_ctrl_apb_PRDATA[31:0]           ), //o
    .axi_ar_valid         (video_ctrl_axi_ar_valid               ), //o
    .axi_ar_ready         (1'b0                                  ), //i
    .axi_ar_payload_addr  (video_ctrl_axi_ar_payload_addr[31:0]  ), //o
    .axi_ar_payload_len   (video_ctrl_axi_ar_payload_len[7:0]    ), //o
    .axi_ar_payload_burst (video_ctrl_axi_ar_payload_burst[1:0]  ), //o
    .axi_r_valid          (1'b0                                  ), //i
    .axi_r_ready          (video_ctrl_axi_r_ready                ), //o
    .axi_r_payload_data   (32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx  ), //i
    .axi_r_payload_last   (1'bx                                  )  //i
  );
  UartController peripheral_uart_ctrl (
    .clk         (board_ctrl_clk_peripheral             ), //i
    .reset       (board_ctrl_reset_peripheral           ), //i
    .uart_rx     (io_uart_rx                            ), //i
    .uart_tx     (peripheral_uart_ctrl_uart_tx          ), //o
    .interrupt   (peripheral_uart_ctrl_interrupt        ), //o
    .apb_PADDR   (peripheral_uart_ctrl_apb_PADDR[3:0]   ), //i
    .apb_PSEL    (apb3Router_2_io_outputs_0_PSEL        ), //i
    .apb_PENABLE (apb3Router_2_io_outputs_0_PENABLE     ), //i
    .apb_PREADY  (peripheral_uart_ctrl_apb_PREADY       ), //o
    .apb_PWRITE  (apb3Router_2_io_outputs_0_PWRITE      ), //i
    .apb_PWDATA  (apb3Router_2_io_outputs_0_PWDATA[31:0]), //i
    .apb_PRDATA  (peripheral_uart_ctrl_apb_PRDATA[31:0] )  //o
  );
  AudioController peripheral_audio_ctrl (
    .clk         (board_ctrl_clk_peripheral             ), //i
    .reset       (board_ctrl_reset_peripheral           ), //i
    .shdn        (peripheral_audio_ctrl_shdn            ), //o
    .i2c_scl     (peripheral_audio_ctrl_i2c_scl         ), //o
    .i2c_sda     (io_audio_i2c_sda                      ), //~
    .apb_PADDR   (peripheral_audio_ctrl_apb_PADDR[2:0]  ), //i
    .apb_PSEL    (apb3Router_2_io_outputs_1_PSEL        ), //i
    .apb_PENABLE (apb3Router_2_io_outputs_1_PENABLE     ), //i
    .apb_PREADY  (peripheral_audio_ctrl_apb_PREADY      ), //o
    .apb_PWRITE  (apb3Router_2_io_outputs_1_PWRITE      ), //i
    .apb_PWDATA  (apb3Router_2_io_outputs_1_PWDATA[31:0]), //i
    .apb_PRDATA  (peripheral_audio_ctrl_apb_PRDATA[31:0])  //o
  );
  SdcardController peripheral_sdcard_ctrl (
    .clk            (board_ctrl_clk_peripheral              ), //i
    .reset          (board_ctrl_reset_peripheral            ), //i
    .sdcard_clk     (peripheral_sdcard_ctrl_sdcard_clk      ), //o
    .sdcard_cmd     (io_sdcard_cmd                          ), //~
    .sdcard_data    (io_sdcard_data                         ), //~
    .sdcard_ndetect (io_sdcard_ndetect                      ), //i
    .interrupt      (peripheral_sdcard_ctrl_interrupt       ), //o
    .apb_PADDR      (peripheral_sdcard_ctrl_apb_PADDR[4:0]  ), //i
    .apb_PSEL       (apb3Router_2_io_outputs_2_PSEL         ), //i
    .apb_PENABLE    (apb3Router_2_io_outputs_2_PENABLE      ), //i
    .apb_PREADY     (peripheral_sdcard_ctrl_apb_PREADY      ), //o
    .apb_PWRITE     (apb3Router_2_io_outputs_2_PWRITE       ), //i
    .apb_PWDATA     (apb3Router_2_io_outputs_2_PWDATA[31:0] ), //i
    .apb_PRDATA     (peripheral_sdcard_ctrl_apb_PRDATA[31:0])  //o
  );
  EndeavourUSB peripheral_usb_ctrl (
    .io_usb1_dp          (io_usb1_dp                                  ), //~
    .io_usb1_dn          (io_usb1_dn                                  ), //~
    .io_usb2_dp          (io_usb2_dp                                  ), //~
    .io_usb2_dn          (io_usb2_dn                                  ), //~
    .io_apb_ctrl_PADDR   (peripheral_usb_ctrl_io_apb_ctrl_PADDR[11:0] ), //i
    .io_apb_ctrl_PSEL    (apb3Router_2_io_outputs_3_PSEL              ), //i
    .io_apb_ctrl_PENABLE (apb3Router_2_io_outputs_3_PENABLE           ), //i
    .io_apb_ctrl_PREADY  (peripheral_usb_ctrl_io_apb_ctrl_PREADY      ), //o
    .io_apb_ctrl_PWRITE  (apb3Router_2_io_outputs_3_PWRITE            ), //i
    .io_apb_ctrl_PWDATA  (apb3Router_2_io_outputs_3_PWDATA[31:0]      ), //i
    .io_apb_ctrl_PRDATA  (peripheral_usb_ctrl_io_apb_ctrl_PRDATA[31:0]), //o
    .io_apb_dma_PADDR    (peripheral_usb_ctrl_io_apb_dma_PADDR[11:0]  ), //i
    .io_apb_dma_PSEL     (apb3Router_2_io_outputs_4_PSEL              ), //i
    .io_apb_dma_PENABLE  (apb3Router_2_io_outputs_4_PENABLE           ), //i
    .io_apb_dma_PREADY   (peripheral_usb_ctrl_io_apb_dma_PREADY       ), //o
    .io_apb_dma_PWRITE   (apb3Router_2_io_outputs_4_PWRITE            ), //i
    .io_apb_dma_PWDATA   (apb3Router_2_io_outputs_4_PWDATA[31:0]      ), //i
    .io_apb_dma_PRDATA   (peripheral_usb_ctrl_io_apb_dma_PRDATA[31:0] ), //o
    .io_interrupt        (peripheral_usb_ctrl_io_interrupt            ), //o
    ._zz_io_interrupt    (peripheral_usb_ctrl__zz_io_interrupt        ), //o
    .clk_peripheral      (board_ctrl_clk_peripheral                   ), //i
    .reset_peripheral    (board_ctrl_reset_peripheral                 )  //i
  );
  Apb3Decoder peripheral_apb_decoder (
    .io_input_PADDR    (peripheral_apb_PADDR[18:0]                   ), //i
    .io_input_PSEL     (peripheral_apb_PSEL                          ), //i
    .io_input_PENABLE  (peripheral_apb_PENABLE                       ), //i
    .io_input_PREADY   (peripheral_apb_decoder_io_input_PREADY       ), //o
    .io_input_PWRITE   (peripheral_apb_PWRITE                        ), //i
    .io_input_PWDATA   (peripheral_apb_PWDATA[31:0]                  ), //i
    .io_input_PRDATA   (peripheral_apb_decoder_io_input_PRDATA[31:0] ), //o
    .io_output_PADDR   (peripheral_apb_decoder_io_output_PADDR[18:0] ), //o
    .io_output_PSEL    (peripheral_apb_decoder_io_output_PSEL[4:0]   ), //o
    .io_output_PENABLE (peripheral_apb_decoder_io_output_PENABLE     ), //o
    .io_output_PREADY  (apb3Router_2_io_input_PREADY                 ), //i
    .io_output_PWRITE  (peripheral_apb_decoder_io_output_PWRITE      ), //o
    .io_output_PWDATA  (peripheral_apb_decoder_io_output_PWDATA[31:0]), //o
    .io_output_PRDATA  (apb3Router_2_io_input_PRDATA[31:0]           )  //i
  );
  Apb3Router apb3Router_2 (
    .io_input_PADDR       (peripheral_apb_decoder_io_output_PADDR[18:0] ), //i
    .io_input_PSEL        (peripheral_apb_decoder_io_output_PSEL[4:0]   ), //i
    .io_input_PENABLE     (peripheral_apb_decoder_io_output_PENABLE     ), //i
    .io_input_PREADY      (apb3Router_2_io_input_PREADY                 ), //o
    .io_input_PWRITE      (peripheral_apb_decoder_io_output_PWRITE      ), //i
    .io_input_PWDATA      (peripheral_apb_decoder_io_output_PWDATA[31:0]), //i
    .io_input_PRDATA      (apb3Router_2_io_input_PRDATA[31:0]           ), //o
    .io_outputs_0_PADDR   (apb3Router_2_io_outputs_0_PADDR[18:0]        ), //o
    .io_outputs_0_PSEL    (apb3Router_2_io_outputs_0_PSEL               ), //o
    .io_outputs_0_PENABLE (apb3Router_2_io_outputs_0_PENABLE            ), //o
    .io_outputs_0_PREADY  (peripheral_uart_ctrl_apb_PREADY              ), //i
    .io_outputs_0_PWRITE  (apb3Router_2_io_outputs_0_PWRITE             ), //o
    .io_outputs_0_PWDATA  (apb3Router_2_io_outputs_0_PWDATA[31:0]       ), //o
    .io_outputs_0_PRDATA  (peripheral_uart_ctrl_apb_PRDATA[31:0]        ), //i
    .io_outputs_1_PADDR   (apb3Router_2_io_outputs_1_PADDR[18:0]        ), //o
    .io_outputs_1_PSEL    (apb3Router_2_io_outputs_1_PSEL               ), //o
    .io_outputs_1_PENABLE (apb3Router_2_io_outputs_1_PENABLE            ), //o
    .io_outputs_1_PREADY  (peripheral_audio_ctrl_apb_PREADY             ), //i
    .io_outputs_1_PWRITE  (apb3Router_2_io_outputs_1_PWRITE             ), //o
    .io_outputs_1_PWDATA  (apb3Router_2_io_outputs_1_PWDATA[31:0]       ), //o
    .io_outputs_1_PRDATA  (peripheral_audio_ctrl_apb_PRDATA[31:0]       ), //i
    .io_outputs_2_PADDR   (apb3Router_2_io_outputs_2_PADDR[18:0]        ), //o
    .io_outputs_2_PSEL    (apb3Router_2_io_outputs_2_PSEL               ), //o
    .io_outputs_2_PENABLE (apb3Router_2_io_outputs_2_PENABLE            ), //o
    .io_outputs_2_PREADY  (peripheral_sdcard_ctrl_apb_PREADY            ), //i
    .io_outputs_2_PWRITE  (apb3Router_2_io_outputs_2_PWRITE             ), //o
    .io_outputs_2_PWDATA  (apb3Router_2_io_outputs_2_PWDATA[31:0]       ), //o
    .io_outputs_2_PRDATA  (peripheral_sdcard_ctrl_apb_PRDATA[31:0]      ), //i
    .io_outputs_3_PADDR   (apb3Router_2_io_outputs_3_PADDR[18:0]        ), //o
    .io_outputs_3_PSEL    (apb3Router_2_io_outputs_3_PSEL               ), //o
    .io_outputs_3_PENABLE (apb3Router_2_io_outputs_3_PENABLE            ), //o
    .io_outputs_3_PREADY  (peripheral_usb_ctrl_io_apb_ctrl_PREADY       ), //i
    .io_outputs_3_PWRITE  (apb3Router_2_io_outputs_3_PWRITE             ), //o
    .io_outputs_3_PWDATA  (apb3Router_2_io_outputs_3_PWDATA[31:0]       ), //o
    .io_outputs_3_PRDATA  (peripheral_usb_ctrl_io_apb_ctrl_PRDATA[31:0] ), //i
    .io_outputs_4_PADDR   (apb3Router_2_io_outputs_4_PADDR[18:0]        ), //o
    .io_outputs_4_PSEL    (apb3Router_2_io_outputs_4_PSEL               ), //o
    .io_outputs_4_PENABLE (apb3Router_2_io_outputs_4_PENABLE            ), //o
    .io_outputs_4_PREADY  (peripheral_usb_ctrl_io_apb_dma_PREADY        ), //i
    .io_outputs_4_PWRITE  (apb3Router_2_io_outputs_4_PWRITE             ), //o
    .io_outputs_4_PWDATA  (apb3Router_2_io_outputs_4_PWDATA[31:0]       ), //o
    .io_outputs_4_PRDATA  (peripheral_usb_ctrl_io_apb_dma_PRDATA[31:0]  ), //i
    .clk_peripheral       (board_ctrl_clk_peripheral                    ), //i
    .reset_peripheral     (board_ctrl_reset_peripheral                  )  //i
  );
  ApbClockBridge #(
    .AWIDTH (19)
  ) peripheral_apb_bridge (
    .clk_input      (board_ctrl_clk_cpu                       ), //i
    .clk_output     (board_ctrl_clk_peripheral                ), //i
    .input_PADDR    (peripheral_apb_bridge_input_PADDR[18:0]  ), //i
    .input_PSEL     (apb3Router_3_io_outputs_0_PSEL           ), //i
    .input_PENABLE  (apb3Router_3_io_outputs_0_PENABLE        ), //i
    .input_PREADY   (peripheral_apb_bridge_input_PREADY       ), //o
    .input_PWRITE   (apb3Router_3_io_outputs_0_PWRITE         ), //i
    .input_PWDATA   (apb3Router_3_io_outputs_0_PWDATA[31:0]   ), //i
    .input_PRDATA   (peripheral_apb_bridge_input_PRDATA[31:0] ), //o
    .output_PADDR   (peripheral_apb_bridge_output_PADDR[18:0] ), //o
    .output_PSEL    (peripheral_apb_bridge_output_PSEL        ), //o
    .output_PENABLE (peripheral_apb_bridge_output_PENABLE     ), //o
    .output_PREADY  (peripheral_apb_PREADY                    ), //i
    .output_PWRITE  (peripheral_apb_bridge_output_PWRITE      ), //o
    .output_PWDATA  (peripheral_apb_bridge_output_PWDATA[31:0]), //o
    .output_PRDATA  (peripheral_apb_PRDATA[31:0]              )  //i
  );
  VexiiRiscv vexiiRiscv_1 (
    .PrivilegedPlugin_logic_rdtime                         (board_ctrl_utime[63:0]                                                  ), //i
    .PrivilegedPlugin_logic_harts_0_int_m_timer            (vexiiRiscv_1_PrivilegedPlugin_logic_harts_0_int_m_timer                 ), //i
    .PrivilegedPlugin_logic_harts_0_int_m_software         (vexiiRiscv_1_PrivilegedPlugin_logic_harts_0_int_m_software              ), //i
    .PrivilegedPlugin_logic_harts_0_int_m_external         (vexiiRiscv_1_PrivilegedPlugin_logic_harts_0_int_m_external              ), //i
    .PrivilegedPlugin_logic_harts_0_int_s_external         (vexiiRiscv_1_PrivilegedPlugin_logic_harts_0_int_s_external              ), //i
    .FetchL1TileLinkPlugin_logic_down_a_valid              (vexiiRiscv_1_FetchL1TileLinkPlugin_logic_down_a_valid                   ), //o
    .FetchL1TileLinkPlugin_logic_down_a_ready              (_zz_FetchL1TileLinkPlugin_logic_down_a_ready                            ), //i
    .FetchL1TileLinkPlugin_logic_down_a_payload_opcode     (vexiiRiscv_1_FetchL1TileLinkPlugin_logic_down_a_payload_opcode[2:0]     ), //o
    .FetchL1TileLinkPlugin_logic_down_a_payload_param      (vexiiRiscv_1_FetchL1TileLinkPlugin_logic_down_a_payload_param[2:0]      ), //o
    .FetchL1TileLinkPlugin_logic_down_a_payload_address    (vexiiRiscv_1_FetchL1TileLinkPlugin_logic_down_a_payload_address[31:0]   ), //o
    .FetchL1TileLinkPlugin_logic_down_a_payload_size       (vexiiRiscv_1_FetchL1TileLinkPlugin_logic_down_a_payload_size[2:0]       ), //o
    .FetchL1TileLinkPlugin_logic_down_d_valid              (_zz_when_Stream_l393                                                    ), //i
    .FetchL1TileLinkPlugin_logic_down_d_ready              (vexiiRiscv_1_FetchL1TileLinkPlugin_logic_down_d_ready                   ), //o
    .FetchL1TileLinkPlugin_logic_down_d_payload_opcode     (_zz_FetchL1TileLinkPlugin_logic_down_d_payload_opcode[2:0]              ), //i
    .FetchL1TileLinkPlugin_logic_down_d_payload_param      (_zz_FetchL1TileLinkPlugin_logic_down_d_payload_param[2:0]               ), //i
    .FetchL1TileLinkPlugin_logic_down_d_payload_size       (_zz_FetchL1TileLinkPlugin_logic_down_d_payload_size[2:0]                ), //i
    .FetchL1TileLinkPlugin_logic_down_d_payload_denied     (_zz_FetchL1TileLinkPlugin_logic_down_d_payload_denied                   ), //i
    .FetchL1TileLinkPlugin_logic_down_d_payload_data       (_zz_FetchL1TileLinkPlugin_logic_down_d_payload_data[63:0]               ), //i
    .FetchL1TileLinkPlugin_logic_down_d_payload_corrupt    (_zz_FetchL1TileLinkPlugin_logic_down_d_payload_corrupt                  ), //i
    .LsuL1TileLinkPlugin_logic_down_a_valid                (vexiiRiscv_1_LsuL1TileLinkPlugin_logic_down_a_valid                     ), //o
    .LsuL1TileLinkPlugin_logic_down_a_ready                (_zz_LsuL1TileLinkPlugin_logic_down_a_ready                              ), //i
    .LsuL1TileLinkPlugin_logic_down_a_payload_opcode       (vexiiRiscv_1_LsuL1TileLinkPlugin_logic_down_a_payload_opcode[2:0]       ), //o
    .LsuL1TileLinkPlugin_logic_down_a_payload_param        (vexiiRiscv_1_LsuL1TileLinkPlugin_logic_down_a_payload_param[2:0]        ), //o
    .LsuL1TileLinkPlugin_logic_down_a_payload_source       (vexiiRiscv_1_LsuL1TileLinkPlugin_logic_down_a_payload_source            ), //o
    .LsuL1TileLinkPlugin_logic_down_a_payload_address      (vexiiRiscv_1_LsuL1TileLinkPlugin_logic_down_a_payload_address[31:0]     ), //o
    .LsuL1TileLinkPlugin_logic_down_a_payload_size         (vexiiRiscv_1_LsuL1TileLinkPlugin_logic_down_a_payload_size[2:0]         ), //o
    .LsuL1TileLinkPlugin_logic_down_a_payload_mask         (vexiiRiscv_1_LsuL1TileLinkPlugin_logic_down_a_payload_mask[7:0]         ), //o
    .LsuL1TileLinkPlugin_logic_down_a_payload_data         (vexiiRiscv_1_LsuL1TileLinkPlugin_logic_down_a_payload_data[63:0]        ), //o
    .LsuL1TileLinkPlugin_logic_down_a_payload_corrupt      (vexiiRiscv_1_LsuL1TileLinkPlugin_logic_down_a_payload_corrupt           ), //o
    .LsuL1TileLinkPlugin_logic_down_d_valid                (_zz_when_Stream_l393_4                                                  ), //i
    .LsuL1TileLinkPlugin_logic_down_d_ready                (vexiiRiscv_1_LsuL1TileLinkPlugin_logic_down_d_ready                     ), //o
    .LsuL1TileLinkPlugin_logic_down_d_payload_opcode       (_zz_LsuL1TileLinkPlugin_logic_down_d_payload_opcode[2:0]                ), //i
    .LsuL1TileLinkPlugin_logic_down_d_payload_param        (_zz_LsuL1TileLinkPlugin_logic_down_d_payload_param[2:0]                 ), //i
    .LsuL1TileLinkPlugin_logic_down_d_payload_source       (_zz_LsuL1TileLinkPlugin_logic_down_d_payload_source                     ), //i
    .LsuL1TileLinkPlugin_logic_down_d_payload_size         (_zz_LsuL1TileLinkPlugin_logic_down_d_payload_size[2:0]                  ), //i
    .LsuL1TileLinkPlugin_logic_down_d_payload_denied       (_zz_LsuL1TileLinkPlugin_logic_down_d_payload_denied                     ), //i
    .LsuL1TileLinkPlugin_logic_down_d_payload_data         (_zz_LsuL1TileLinkPlugin_logic_down_d_payload_data[63:0]                 ), //i
    .LsuL1TileLinkPlugin_logic_down_d_payload_corrupt      (_zz_LsuL1TileLinkPlugin_logic_down_d_payload_corrupt                    ), //i
    .LsuTileLinkPlugin_logic_bridge_down_a_valid           (vexiiRiscv_1_LsuTileLinkPlugin_logic_bridge_down_a_valid                ), //o
    .LsuTileLinkPlugin_logic_bridge_down_a_ready           (_zz_LsuTileLinkPlugin_logic_bridge_down_a_ready                         ), //i
    .LsuTileLinkPlugin_logic_bridge_down_a_payload_opcode  (vexiiRiscv_1_LsuTileLinkPlugin_logic_bridge_down_a_payload_opcode[2:0]  ), //o
    .LsuTileLinkPlugin_logic_bridge_down_a_payload_param   (vexiiRiscv_1_LsuTileLinkPlugin_logic_bridge_down_a_payload_param[2:0]   ), //o
    .LsuTileLinkPlugin_logic_bridge_down_a_payload_address (vexiiRiscv_1_LsuTileLinkPlugin_logic_bridge_down_a_payload_address[31:0]), //o
    .LsuTileLinkPlugin_logic_bridge_down_a_payload_size    (vexiiRiscv_1_LsuTileLinkPlugin_logic_bridge_down_a_payload_size[1:0]    ), //o
    .LsuTileLinkPlugin_logic_bridge_down_a_payload_mask    (vexiiRiscv_1_LsuTileLinkPlugin_logic_bridge_down_a_payload_mask[3:0]    ), //o
    .LsuTileLinkPlugin_logic_bridge_down_a_payload_data    (vexiiRiscv_1_LsuTileLinkPlugin_logic_bridge_down_a_payload_data[31:0]   ), //o
    .LsuTileLinkPlugin_logic_bridge_down_a_payload_corrupt (vexiiRiscv_1_LsuTileLinkPlugin_logic_bridge_down_a_payload_corrupt      ), //o
    .LsuTileLinkPlugin_logic_bridge_down_d_valid           (_zz_when_Stream_l393_2                                                  ), //i
    .LsuTileLinkPlugin_logic_bridge_down_d_ready           (vexiiRiscv_1_LsuTileLinkPlugin_logic_bridge_down_d_ready                ), //o
    .LsuTileLinkPlugin_logic_bridge_down_d_payload_opcode  (_zz_LsuTileLinkPlugin_logic_bridge_down_d_payload_opcode[2:0]           ), //i
    .LsuTileLinkPlugin_logic_bridge_down_d_payload_param   (_zz_LsuTileLinkPlugin_logic_bridge_down_d_payload_param[2:0]            ), //i
    .LsuTileLinkPlugin_logic_bridge_down_d_payload_size    (_zz_LsuTileLinkPlugin_logic_bridge_down_d_payload_size[1:0]             ), //i
    .LsuTileLinkPlugin_logic_bridge_down_d_payload_denied  (_zz_LsuTileLinkPlugin_logic_bridge_down_d_payload_denied                ), //i
    .LsuTileLinkPlugin_logic_bridge_down_d_payload_data    (_zz_LsuTileLinkPlugin_logic_bridge_down_d_payload_data[31:0]            ), //i
    .LsuTileLinkPlugin_logic_bridge_down_d_payload_corrupt (_zz_LsuTileLinkPlugin_logic_bridge_down_d_payload_corrupt               ), //i
    .clk_cpu                                               (board_ctrl_clk_cpu                                                      ), //i
    .reset_cpu                                             (board_ctrl_reset_cpu                                                    )  //i
  );
  Arbiter arbiter_1 (
    .io_ups_0_a_valid           (_zz_io_ups_0_a_valid                          ), //i
    .io_ups_0_a_ready           (arbiter_1_io_ups_0_a_ready                    ), //o
    .io_ups_0_a_payload_opcode  (_zz_io_ups_0_a_payload_opcode_6[2:0]          ), //i
    .io_ups_0_a_payload_param   (_zz_io_ups_0_a_payload_param_1[2:0]           ), //i
    .io_ups_0_a_payload_address (_zz_io_ups_0_a_payload_address_1[31:0]        ), //i
    .io_ups_0_a_payload_size    (_zz_io_ups_0_a_payload_size_1[2:0]            ), //i
    .io_ups_0_d_valid           (arbiter_1_io_ups_0_d_valid                    ), //o
    .io_ups_0_d_ready           (_zz_io_ups_0_d_ready                          ), //i
    .io_ups_0_d_payload_opcode  (arbiter_1_io_ups_0_d_payload_opcode[2:0]      ), //o
    .io_ups_0_d_payload_param   (arbiter_1_io_ups_0_d_payload_param[2:0]       ), //o
    .io_ups_0_d_payload_size    (arbiter_1_io_ups_0_d_payload_size[2:0]        ), //o
    .io_ups_0_d_payload_denied  (arbiter_1_io_ups_0_d_payload_denied           ), //o
    .io_ups_0_d_payload_data    (arbiter_1_io_ups_0_d_payload_data[63:0]       ), //o
    .io_ups_0_d_payload_corrupt (arbiter_1_io_ups_0_d_payload_corrupt          ), //o
    .io_ups_1_a_valid           (widthAdapter_2_io_down_a_valid                ), //i
    .io_ups_1_a_ready           (arbiter_1_io_ups_1_a_ready                    ), //o
    .io_ups_1_a_payload_opcode  (_zz_io_ups_1_a_payload_opcode[2:0]            ), //i
    .io_ups_1_a_payload_param   (widthAdapter_2_io_down_a_payload_param[2:0]   ), //i
    .io_ups_1_a_payload_address (widthAdapter_2_io_down_a_payload_address[31:0]), //i
    .io_ups_1_a_payload_size    (widthAdapter_2_io_down_a_payload_size[1:0]    ), //i
    .io_ups_1_a_payload_mask    (widthAdapter_2_io_down_a_payload_mask[7:0]    ), //i
    .io_ups_1_a_payload_data    (widthAdapter_2_io_down_a_payload_data[63:0]   ), //i
    .io_ups_1_a_payload_corrupt (widthAdapter_2_io_down_a_payload_corrupt      ), //i
    .io_ups_1_d_valid           (arbiter_1_io_ups_1_d_valid                    ), //o
    .io_ups_1_d_ready           (widthAdapter_2_io_down_d_ready                ), //i
    .io_ups_1_d_payload_opcode  (arbiter_1_io_ups_1_d_payload_opcode[2:0]      ), //o
    .io_ups_1_d_payload_param   (arbiter_1_io_ups_1_d_payload_param[2:0]       ), //o
    .io_ups_1_d_payload_size    (arbiter_1_io_ups_1_d_payload_size[1:0]        ), //o
    .io_ups_1_d_payload_denied  (arbiter_1_io_ups_1_d_payload_denied           ), //o
    .io_ups_1_d_payload_data    (arbiter_1_io_ups_1_d_payload_data[63:0]       ), //o
    .io_ups_1_d_payload_corrupt (arbiter_1_io_ups_1_d_payload_corrupt          ), //o
    .io_ups_2_a_valid           (_zz_io_ups_2_a_valid                          ), //i
    .io_ups_2_a_ready           (arbiter_1_io_ups_2_a_ready                    ), //o
    .io_ups_2_a_payload_opcode  (_zz_io_ups_2_a_payload_opcode_4[2:0]          ), //i
    .io_ups_2_a_payload_param   (_zz_io_ups_2_a_payload_param[2:0]             ), //i
    .io_ups_2_a_payload_source  (_zz_io_ups_2_a_payload_source                 ), //i
    .io_ups_2_a_payload_address (_zz_io_ups_2_a_payload_address[31:0]          ), //i
    .io_ups_2_a_payload_size    (_zz_io_ups_2_a_payload_size[2:0]              ), //i
    .io_ups_2_a_payload_mask    (_zz_io_ups_2_a_payload_mask[7:0]              ), //i
    .io_ups_2_a_payload_data    (_zz_io_ups_2_a_payload_data[63:0]             ), //i
    .io_ups_2_a_payload_corrupt (_zz_io_ups_2_a_payload_corrupt                ), //i
    .io_ups_2_d_valid           (arbiter_1_io_ups_2_d_valid                    ), //o
    .io_ups_2_d_ready           (_zz_io_ups_2_d_ready                          ), //i
    .io_ups_2_d_payload_opcode  (arbiter_1_io_ups_2_d_payload_opcode[2:0]      ), //o
    .io_ups_2_d_payload_param   (arbiter_1_io_ups_2_d_payload_param[2:0]       ), //o
    .io_ups_2_d_payload_source  (arbiter_1_io_ups_2_d_payload_source           ), //o
    .io_ups_2_d_payload_size    (arbiter_1_io_ups_2_d_payload_size[2:0]        ), //o
    .io_ups_2_d_payload_denied  (arbiter_1_io_ups_2_d_payload_denied           ), //o
    .io_ups_2_d_payload_data    (arbiter_1_io_ups_2_d_payload_data[63:0]       ), //o
    .io_ups_2_d_payload_corrupt (arbiter_1_io_ups_2_d_payload_corrupt          ), //o
    .io_down_a_valid            (arbiter_1_io_down_a_valid                     ), //o
    .io_down_a_ready            (decoder_2_io_up_a_ready                       ), //i
    .io_down_a_payload_opcode   (arbiter_1_io_down_a_payload_opcode[2:0]       ), //o
    .io_down_a_payload_param    (arbiter_1_io_down_a_payload_param[2:0]        ), //o
    .io_down_a_payload_source   (arbiter_1_io_down_a_payload_source[2:0]       ), //o
    .io_down_a_payload_address  (arbiter_1_io_down_a_payload_address[31:0]     ), //o
    .io_down_a_payload_size     (arbiter_1_io_down_a_payload_size[2:0]         ), //o
    .io_down_a_payload_mask     (arbiter_1_io_down_a_payload_mask[7:0]         ), //o
    .io_down_a_payload_data     (arbiter_1_io_down_a_payload_data[63:0]        ), //o
    .io_down_a_payload_corrupt  (arbiter_1_io_down_a_payload_corrupt           ), //o
    .io_down_d_valid            (decoder_2_io_up_d_valid                       ), //i
    .io_down_d_ready            (arbiter_1_io_down_d_ready                     ), //o
    .io_down_d_payload_opcode   (_zz_io_down_d_payload_opcode[2:0]             ), //i
    .io_down_d_payload_param    (decoder_2_io_up_d_payload_param[2:0]          ), //i
    .io_down_d_payload_source   (decoder_2_io_up_d_payload_source[2:0]         ), //i
    .io_down_d_payload_size     (decoder_2_io_up_d_payload_size[2:0]           ), //i
    .io_down_d_payload_denied   (decoder_2_io_up_d_payload_denied              ), //i
    .io_down_d_payload_data     (decoder_2_io_up_d_payload_data[63:0]          ), //i
    .io_down_d_payload_corrupt  (decoder_2_io_up_d_payload_corrupt             ), //i
    .clk_cpu                    (board_ctrl_clk_cpu                            ), //i
    .reset_cpu                  (board_ctrl_reset_cpu                          )  //i
  );
  Axi4Bridge ramBridge_logic_bridge (
    .io_up_a_valid              (ramBridge_up_bus_a_valid                            ), //i
    .io_up_a_ready              (ramBridge_logic_bridge_io_up_a_ready                ), //o
    .io_up_a_payload_opcode     (ramBridge_up_bus_a_payload_opcode[2:0]              ), //i
    .io_up_a_payload_param      (ramBridge_up_bus_a_payload_param[2:0]               ), //i
    .io_up_a_payload_source     (ramBridge_up_bus_a_payload_source[2:0]              ), //i
    .io_up_a_payload_address    (ramBridge_up_bus_a_payload_address[26:0]            ), //i
    .io_up_a_payload_size       (ramBridge_up_bus_a_payload_size[2:0]                ), //i
    .io_up_a_payload_mask       (ramBridge_up_bus_a_payload_mask[7:0]                ), //i
    .io_up_a_payload_data       (ramBridge_up_bus_a_payload_data[63:0]               ), //i
    .io_up_a_payload_corrupt    (ramBridge_up_bus_a_payload_corrupt                  ), //i
    .io_up_d_valid              (ramBridge_logic_bridge_io_up_d_valid                ), //o
    .io_up_d_ready              (ramBridge_up_bus_d_ready                            ), //i
    .io_up_d_payload_opcode     (ramBridge_logic_bridge_io_up_d_payload_opcode[2:0]  ), //o
    .io_up_d_payload_param      (ramBridge_logic_bridge_io_up_d_payload_param[2:0]   ), //o
    .io_up_d_payload_source     (ramBridge_logic_bridge_io_up_d_payload_source[2:0]  ), //o
    .io_up_d_payload_size       (ramBridge_logic_bridge_io_up_d_payload_size[2:0]    ), //o
    .io_up_d_payload_denied     (ramBridge_logic_bridge_io_up_d_payload_denied       ), //o
    .io_up_d_payload_data       (ramBridge_logic_bridge_io_up_d_payload_data[63:0]   ), //o
    .io_up_d_payload_corrupt    (ramBridge_logic_bridge_io_up_d_payload_corrupt      ), //o
    .io_down_aw_valid           (ramBridge_logic_bridge_io_down_aw_valid             ), //o
    .io_down_aw_ready           (ramBridge_down_aw_ready                             ), //i
    .io_down_aw_payload_addr    (ramBridge_logic_bridge_io_down_aw_payload_addr[26:0]), //o
    .io_down_aw_payload_id      (ramBridge_logic_bridge_io_down_aw_payload_id[2:0]   ), //o
    .io_down_aw_payload_len     (ramBridge_logic_bridge_io_down_aw_payload_len[7:0]  ), //o
    .io_down_aw_payload_size    (ramBridge_logic_bridge_io_down_aw_payload_size[2:0] ), //o
    .io_down_aw_payload_burst   (ramBridge_logic_bridge_io_down_aw_payload_burst[1:0]), //o
    .io_down_aw_payload_allStrb (ramBridge_logic_bridge_io_down_aw_payload_allStrb   ), //o
    .io_down_w_valid            (ramBridge_logic_bridge_io_down_w_valid              ), //o
    .io_down_w_ready            (ramBridge_down_w_ready                              ), //i
    .io_down_w_payload_data     (ramBridge_logic_bridge_io_down_w_payload_data[63:0] ), //o
    .io_down_w_payload_strb     (ramBridge_logic_bridge_io_down_w_payload_strb[7:0]  ), //o
    .io_down_w_payload_last     (ramBridge_logic_bridge_io_down_w_payload_last       ), //o
    .io_down_b_valid            (ramBridge_down_b_valid                              ), //i
    .io_down_b_ready            (ramBridge_logic_bridge_io_down_b_ready              ), //o
    .io_down_b_payload_id       (ramBridge_down_b_payload_id[2:0]                    ), //i
    .io_down_b_payload_resp     (ramBridge_down_b_payload_resp[1:0]                  ), //i
    .io_down_ar_valid           (ramBridge_logic_bridge_io_down_ar_valid             ), //o
    .io_down_ar_ready           (ramBridge_down_ar_ready                             ), //i
    .io_down_ar_payload_addr    (ramBridge_logic_bridge_io_down_ar_payload_addr[26:0]), //o
    .io_down_ar_payload_id      (ramBridge_logic_bridge_io_down_ar_payload_id[2:0]   ), //o
    .io_down_ar_payload_len     (ramBridge_logic_bridge_io_down_ar_payload_len[7:0]  ), //o
    .io_down_ar_payload_size    (ramBridge_logic_bridge_io_down_ar_payload_size[2:0] ), //o
    .io_down_ar_payload_burst   (ramBridge_logic_bridge_io_down_ar_payload_burst[1:0]), //o
    .io_down_r_valid            (ramBridge_down_r_valid                              ), //i
    .io_down_r_ready            (ramBridge_logic_bridge_io_down_r_ready              ), //o
    .io_down_r_payload_data     (ramBridge_down_r_payload_data[63:0]                 ), //i
    .io_down_r_payload_id       (ramBridge_down_r_payload_id[2:0]                    ), //i
    .io_down_r_payload_resp     (ramBridge_down_r_payload_resp[1:0]                  ), //i
    .io_down_r_payload_last     (ramBridge_down_r_payload_last                       ), //i
    .clk_cpu                    (board_ctrl_clk_cpu                                  ), //i
    .reset_cpu                  (board_ctrl_reset_cpu                                )  //i
  );
  WidthAdapter widthAdapter_2 (
    .io_up_a_valid             (_zz_io_up_a_valid                             ), //i
    .io_up_a_ready             (widthAdapter_2_io_up_a_ready                  ), //o
    .io_up_a_payload_opcode    (_zz_io_up_a_payload_opcode_7[2:0]             ), //i
    .io_up_a_payload_param     (_zz_io_up_a_payload_param[2:0]                ), //i
    .io_up_a_payload_address   (_zz_io_up_a_payload_address[31:0]             ), //i
    .io_up_a_payload_size      (_zz_io_up_a_payload_size[1:0]                 ), //i
    .io_up_a_payload_mask      (_zz_io_up_a_payload_mask[3:0]                 ), //i
    .io_up_a_payload_data      (_zz_io_up_a_payload_data[31:0]                ), //i
    .io_up_a_payload_corrupt   (_zz_io_up_a_payload_corrupt                   ), //i
    .io_up_d_valid             (widthAdapter_2_io_up_d_valid                  ), //o
    .io_up_d_ready             (_zz_io_up_d_ready                             ), //i
    .io_up_d_payload_opcode    (widthAdapter_2_io_up_d_payload_opcode[2:0]    ), //o
    .io_up_d_payload_param     (widthAdapter_2_io_up_d_payload_param[2:0]     ), //o
    .io_up_d_payload_size      (widthAdapter_2_io_up_d_payload_size[1:0]      ), //o
    .io_up_d_payload_denied    (widthAdapter_2_io_up_d_payload_denied         ), //o
    .io_up_d_payload_data      (widthAdapter_2_io_up_d_payload_data[31:0]     ), //o
    .io_up_d_payload_corrupt   (widthAdapter_2_io_up_d_payload_corrupt        ), //o
    .io_down_a_valid           (widthAdapter_2_io_down_a_valid                ), //o
    .io_down_a_ready           (arbiter_1_io_ups_1_a_ready                    ), //i
    .io_down_a_payload_opcode  (widthAdapter_2_io_down_a_payload_opcode[2:0]  ), //o
    .io_down_a_payload_param   (widthAdapter_2_io_down_a_payload_param[2:0]   ), //o
    .io_down_a_payload_address (widthAdapter_2_io_down_a_payload_address[31:0]), //o
    .io_down_a_payload_size    (widthAdapter_2_io_down_a_payload_size[1:0]    ), //o
    .io_down_a_payload_mask    (widthAdapter_2_io_down_a_payload_mask[7:0]    ), //o
    .io_down_a_payload_data    (widthAdapter_2_io_down_a_payload_data[63:0]   ), //o
    .io_down_a_payload_corrupt (widthAdapter_2_io_down_a_payload_corrupt      ), //o
    .io_down_d_valid           (arbiter_1_io_ups_1_d_valid                    ), //i
    .io_down_d_ready           (widthAdapter_2_io_down_d_ready                ), //o
    .io_down_d_payload_opcode  (_zz_io_down_d_payload_opcode_1[2:0]           ), //i
    .io_down_d_payload_param   (arbiter_1_io_ups_1_d_payload_param[2:0]       ), //i
    .io_down_d_payload_size    (arbiter_1_io_ups_1_d_payload_size[1:0]        ), //i
    .io_down_d_payload_denied  (arbiter_1_io_ups_1_d_payload_denied           ), //i
    .io_down_d_payload_data    (arbiter_1_io_ups_1_d_payload_data[63:0]       ), //i
    .io_down_d_payload_corrupt (arbiter_1_io_ups_1_d_payload_corrupt          ), //i
    .clk_cpu                   (board_ctrl_clk_cpu                            ), //i
    .reset_cpu                 (board_ctrl_reset_cpu                          )  //i
  );
  StreamArbiter_9 streamArbiter_10 (
    .io_inputs_0_valid           (ramBridge_down_ar_valid                      ), //i
    .io_inputs_0_ready           (streamArbiter_10_io_inputs_0_ready           ), //o
    .io_inputs_0_payload_addr    (ramBridge_down_ar_payload_addr[26:0]         ), //i
    .io_inputs_0_payload_id      (ramBridge_down_ar_payload_id[2:0]            ), //i
    .io_inputs_0_payload_len     (ramBridge_down_ar_payload_len[7:0]           ), //i
    .io_inputs_0_payload_size    (ramBridge_down_ar_payload_size[2:0]          ), //i
    .io_inputs_0_payload_burst   (ramBridge_down_ar_payload_burst[1:0]         ), //i
    .io_inputs_0_payload_allStrb (1'b0                                         ), //i
    .io_inputs_1_valid           (ramBridge_down_aw_valid                      ), //i
    .io_inputs_1_ready           (streamArbiter_10_io_inputs_1_ready           ), //o
    .io_inputs_1_payload_addr    (ramBridge_down_aw_payload_addr[26:0]         ), //i
    .io_inputs_1_payload_id      (ramBridge_down_aw_payload_id[2:0]            ), //i
    .io_inputs_1_payload_len     (ramBridge_down_aw_payload_len[7:0]           ), //i
    .io_inputs_1_payload_size    (ramBridge_down_aw_payload_size[2:0]          ), //i
    .io_inputs_1_payload_burst   (ramBridge_down_aw_payload_burst[1:0]         ), //i
    .io_inputs_1_payload_allStrb (ramBridge_down_aw_payload_allStrb            ), //i
    .io_output_valid             (streamArbiter_10_io_output_valid             ), //o
    .io_output_ready             (ram_axi_arw_ready                            ), //i
    .io_output_payload_addr      (streamArbiter_10_io_output_payload_addr[26:0]), //o
    .io_output_payload_id        (streamArbiter_10_io_output_payload_id[2:0]   ), //o
    .io_output_payload_len       (streamArbiter_10_io_output_payload_len[7:0]  ), //o
    .io_output_payload_size      (streamArbiter_10_io_output_payload_size[2:0] ), //o
    .io_output_payload_burst     (streamArbiter_10_io_output_payload_burst[1:0]), //o
    .io_output_payload_allStrb   (streamArbiter_10_io_output_payload_allStrb   ), //o
    .io_chosen                   (streamArbiter_10_io_chosen                   ), //o
    .io_chosenOH                 (streamArbiter_10_io_chosenOH[1:0]            ), //o
    .clk_cpu                     (board_ctrl_clk_cpu                           ), //i
    .reset_cpu                   (board_ctrl_reset_cpu                         )  //i
  );
  DDRSdramController #(
    .ROW_BITS (14),
    .COL_BITS (10),
    .ID_WIDTH (3 )
  ) ram_ddr_ctrl (
    .clk         (board_ctrl_clk_ram_bus                     ), //i
    .clk_shifted (board_ctrl_clk_ram                         ), //i
    .reset       (board_ctrl_reset_ram                       ), //i
    .arw_valid   (ram_axi_cc_io_output_arw_valid             ), //i
    .arw_ready   (ram_ddr_ctrl_arw_ready                     ), //o
    .arw_addr    (ram_axi_cc_io_output_arw_payload_addr[26:0]), //i
    .arw_id      (ram_axi_cc_io_output_arw_payload_id[2:0]   ), //i
    .arw_len     (ram_axi_cc_io_output_arw_payload_len[7:0]  ), //i
    .arw_size    (ram_axi_cc_io_output_arw_payload_size[2:0] ), //i
    .arw_burst   (ram_axi_cc_io_output_arw_payload_burst[1:0]), //i
    .arw_allStrb (ram_axi_cc_io_output_arw_payload_allStrb   ), //i
    .arw_write   (ram_axi_cc_io_output_arw_payload_write     ), //i
    .wvalid      (ram_axi_cc_io_output_w_valid               ), //i
    .wready      (ram_ddr_ctrl_wready                        ), //o
    .wdata       (ram_axi_cc_io_output_w_payload_data[63:0]  ), //i
    .wstrb       (ram_axi_cc_io_output_w_payload_strb[7:0]   ), //i
    .wlast       (ram_axi_cc_io_output_w_payload_last        ), //i
    .bvalid      (ram_ddr_ctrl_bvalid                        ), //o
    .bready      (ram_axi_cc_io_output_b_ready               ), //i
    .bid         (ram_ddr_ctrl_bid[2:0]                      ), //o
    .bresp       (ram_ddr_ctrl_bresp[1:0]                    ), //o
    .rvalid      (ram_ddr_ctrl_rvalid                        ), //o
    .rready      (ram_axi_cc_io_output_r_ready               ), //i
    .rdata       (ram_ddr_ctrl_rdata[63:0]                   ), //o
    .rid         (ram_ddr_ctrl_rid[2:0]                      ), //o
    .rresp       (ram_ddr_ctrl_rresp[1:0]                    ), //o
    .rlast       (ram_ddr_ctrl_rlast                         ), //o
    .ddr_ck_p    (ram_ddr_ctrl_ddr_ck_p                      ), //o
    .ddr_ck_n    (ram_ddr_ctrl_ddr_ck_n                      ), //o
    .ddr_cke     (ram_ddr_ctrl_ddr_cke                       ), //o
    .ddr_ras_n   (ram_ddr_ctrl_ddr_ras_n                     ), //o
    .ddr_cas_n   (ram_ddr_ctrl_ddr_cas_n                     ), //o
    .ddr_we_n    (ram_ddr_ctrl_ddr_we_n                      ), //o
    .ddr_ba      (ram_ddr_ctrl_ddr_ba[1:0]                   ), //o
    .ddr_a       (ram_ddr_ctrl_ddr_a[13:0]                   ), //o
    .ddr_dm      (ram_ddr_ctrl_ddr_dm[1:0]                   ), //o
    .ddr_dqs     (io_ddr_sdram_dqs                           ), //~
    .ddr_dq      (io_ddr_sdram_dq                            )  //~
  );
  Axi4SharedCC ram_axi_cc (
    .io_input_arw_valid            (ram_axi_arw_valid                          ), //i
    .io_input_arw_ready            (ram_axi_cc_io_input_arw_ready              ), //o
    .io_input_arw_payload_addr     (ram_axi_arw_payload_addr[26:0]             ), //i
    .io_input_arw_payload_id       (ram_axi_arw_payload_id[2:0]                ), //i
    .io_input_arw_payload_len      (ram_axi_arw_payload_len[7:0]               ), //i
    .io_input_arw_payload_size     (ram_axi_arw_payload_size[2:0]              ), //i
    .io_input_arw_payload_burst    (ram_axi_arw_payload_burst[1:0]             ), //i
    .io_input_arw_payload_allStrb  (ram_axi_arw_payload_allStrb                ), //i
    .io_input_arw_payload_write    (ram_axi_arw_payload_write                  ), //i
    .io_input_w_valid              (ram_axi_w_valid                            ), //i
    .io_input_w_ready              (ram_axi_cc_io_input_w_ready                ), //o
    .io_input_w_payload_data       (ram_axi_w_payload_data[63:0]               ), //i
    .io_input_w_payload_strb       (ram_axi_w_payload_strb[7:0]                ), //i
    .io_input_w_payload_last       (ram_axi_w_payload_last                     ), //i
    .io_input_b_valid              (ram_axi_cc_io_input_b_valid                ), //o
    .io_input_b_ready              (ram_axi_b_ready                            ), //i
    .io_input_b_payload_id         (ram_axi_cc_io_input_b_payload_id[2:0]      ), //o
    .io_input_b_payload_resp       (ram_axi_cc_io_input_b_payload_resp[1:0]    ), //o
    .io_input_r_valid              (ram_axi_cc_io_input_r_valid                ), //o
    .io_input_r_ready              (ram_axi_r_ready                            ), //i
    .io_input_r_payload_data       (ram_axi_cc_io_input_r_payload_data[63:0]   ), //o
    .io_input_r_payload_id         (ram_axi_cc_io_input_r_payload_id[2:0]      ), //o
    .io_input_r_payload_resp       (ram_axi_cc_io_input_r_payload_resp[1:0]    ), //o
    .io_input_r_payload_last       (ram_axi_cc_io_input_r_payload_last         ), //o
    .io_output_arw_valid           (ram_axi_cc_io_output_arw_valid             ), //o
    .io_output_arw_ready           (ram_ddr_ctrl_arw_ready                     ), //i
    .io_output_arw_payload_addr    (ram_axi_cc_io_output_arw_payload_addr[26:0]), //o
    .io_output_arw_payload_id      (ram_axi_cc_io_output_arw_payload_id[2:0]   ), //o
    .io_output_arw_payload_len     (ram_axi_cc_io_output_arw_payload_len[7:0]  ), //o
    .io_output_arw_payload_size    (ram_axi_cc_io_output_arw_payload_size[2:0] ), //o
    .io_output_arw_payload_burst   (ram_axi_cc_io_output_arw_payload_burst[1:0]), //o
    .io_output_arw_payload_allStrb (ram_axi_cc_io_output_arw_payload_allStrb   ), //o
    .io_output_arw_payload_write   (ram_axi_cc_io_output_arw_payload_write     ), //o
    .io_output_w_valid             (ram_axi_cc_io_output_w_valid               ), //o
    .io_output_w_ready             (ram_ddr_ctrl_wready                        ), //i
    .io_output_w_payload_data      (ram_axi_cc_io_output_w_payload_data[63:0]  ), //o
    .io_output_w_payload_strb      (ram_axi_cc_io_output_w_payload_strb[7:0]   ), //o
    .io_output_w_payload_last      (ram_axi_cc_io_output_w_payload_last        ), //o
    .io_output_b_valid             (ram_ddr_ctrl_bvalid                        ), //i
    .io_output_b_ready             (ram_axi_cc_io_output_b_ready               ), //o
    .io_output_b_payload_id        (ram_ddr_ctrl_bid[2:0]                      ), //i
    .io_output_b_payload_resp      (ram_ddr_ctrl_bresp[1:0]                    ), //i
    .io_output_r_valid             (ram_ddr_ctrl_rvalid                        ), //i
    .io_output_r_ready             (ram_axi_cc_io_output_r_ready               ), //o
    .io_output_r_payload_data      (ram_ddr_ctrl_rdata[63:0]                   ), //i
    .io_output_r_payload_id        (ram_ddr_ctrl_rid[2:0]                      ), //i
    .io_output_r_payload_resp      (ram_ddr_ctrl_rresp[1:0]                    ), //i
    .io_output_r_payload_last      (ram_ddr_ctrl_rlast                         ), //i
    .clk_cpu                       (board_ctrl_clk_cpu                         ), //i
    .reset_cpu                     (board_ctrl_reset_cpu                       ), //i
    .clk_ram_bus                   (board_ctrl_clk_ram_bus                     ), //i
    .reset_ram                     (board_ctrl_reset_ram                       )  //i
  );
  Decoder decoder_2 (
    .io_up_a_valid                (arbiter_1_io_down_a_valid                   ), //i
    .io_up_a_ready                (decoder_2_io_up_a_ready                     ), //o
    .io_up_a_payload_opcode       (_zz_io_up_a_payload_opcode_4[2:0]           ), //i
    .io_up_a_payload_param        (arbiter_1_io_down_a_payload_param[2:0]      ), //i
    .io_up_a_payload_source       (arbiter_1_io_down_a_payload_source[2:0]     ), //i
    .io_up_a_payload_address      (arbiter_1_io_down_a_payload_address[31:0]   ), //i
    .io_up_a_payload_size         (arbiter_1_io_down_a_payload_size[2:0]       ), //i
    .io_up_a_payload_mask         (arbiter_1_io_down_a_payload_mask[7:0]       ), //i
    .io_up_a_payload_data         (arbiter_1_io_down_a_payload_data[63:0]      ), //i
    .io_up_a_payload_corrupt      (arbiter_1_io_down_a_payload_corrupt         ), //i
    .io_up_d_valid                (decoder_2_io_up_d_valid                     ), //o
    .io_up_d_ready                (arbiter_1_io_down_d_ready                   ), //i
    .io_up_d_payload_opcode       (decoder_2_io_up_d_payload_opcode[2:0]       ), //o
    .io_up_d_payload_param        (decoder_2_io_up_d_payload_param[2:0]        ), //o
    .io_up_d_payload_source       (decoder_2_io_up_d_payload_source[2:0]       ), //o
    .io_up_d_payload_size         (decoder_2_io_up_d_payload_size[2:0]         ), //o
    .io_up_d_payload_denied       (decoder_2_io_up_d_payload_denied            ), //o
    .io_up_d_payload_data         (decoder_2_io_up_d_payload_data[63:0]        ), //o
    .io_up_d_payload_corrupt      (decoder_2_io_up_d_payload_corrupt           ), //o
    .io_downs_0_a_valid           (decoder_2_io_downs_0_a_valid                ), //o
    .io_downs_0_a_ready           (widthAdapter_3_io_up_a_ready                ), //i
    .io_downs_0_a_payload_opcode  (decoder_2_io_downs_0_a_payload_opcode[2:0]  ), //o
    .io_downs_0_a_payload_param   (decoder_2_io_downs_0_a_payload_param[2:0]   ), //o
    .io_downs_0_a_payload_source  (decoder_2_io_downs_0_a_payload_source[2:0]  ), //o
    .io_downs_0_a_payload_address (decoder_2_io_downs_0_a_payload_address[30:0]), //o
    .io_downs_0_a_payload_size    (decoder_2_io_downs_0_a_payload_size[2:0]    ), //o
    .io_downs_0_a_payload_mask    (decoder_2_io_downs_0_a_payload_mask[7:0]    ), //o
    .io_downs_0_a_payload_data    (decoder_2_io_downs_0_a_payload_data[63:0]   ), //o
    .io_downs_0_a_payload_corrupt (decoder_2_io_downs_0_a_payload_corrupt      ), //o
    .io_downs_0_d_valid           (widthAdapter_3_io_up_d_valid                ), //i
    .io_downs_0_d_ready           (decoder_2_io_downs_0_d_ready                ), //o
    .io_downs_0_d_payload_opcode  (_zz_io_downs_0_d_payload_opcode_1[2:0]      ), //i
    .io_downs_0_d_payload_param   (widthAdapter_3_io_up_d_payload_param[2:0]   ), //i
    .io_downs_0_d_payload_source  (widthAdapter_3_io_up_d_payload_source[2:0]  ), //i
    .io_downs_0_d_payload_size    (widthAdapter_3_io_up_d_payload_size[2:0]    ), //i
    .io_downs_0_d_payload_denied  (widthAdapter_3_io_up_d_payload_denied       ), //i
    .io_downs_0_d_payload_data    (widthAdapter_3_io_up_d_payload_data[63:0]   ), //i
    .io_downs_0_d_payload_corrupt (widthAdapter_3_io_up_d_payload_corrupt      ), //i
    .io_downs_1_a_valid           (decoder_2_io_downs_1_a_valid                ), //o
    .io_downs_1_a_ready           (ramBridge_up_bus_a_ready                    ), //i
    .io_downs_1_a_payload_opcode  (decoder_2_io_downs_1_a_payload_opcode[2:0]  ), //o
    .io_downs_1_a_payload_param   (decoder_2_io_downs_1_a_payload_param[2:0]   ), //o
    .io_downs_1_a_payload_source  (decoder_2_io_downs_1_a_payload_source[2:0]  ), //o
    .io_downs_1_a_payload_address (decoder_2_io_downs_1_a_payload_address[26:0]), //o
    .io_downs_1_a_payload_size    (decoder_2_io_downs_1_a_payload_size[2:0]    ), //o
    .io_downs_1_a_payload_mask    (decoder_2_io_downs_1_a_payload_mask[7:0]    ), //o
    .io_downs_1_a_payload_data    (decoder_2_io_downs_1_a_payload_data[63:0]   ), //o
    .io_downs_1_a_payload_corrupt (decoder_2_io_downs_1_a_payload_corrupt      ), //o
    .io_downs_1_d_valid           (ramBridge_up_bus_d_valid                    ), //i
    .io_downs_1_d_ready           (decoder_2_io_downs_1_d_ready                ), //o
    .io_downs_1_d_payload_opcode  (_zz_io_downs_1_d_payload_opcode_2[2:0]      ), //i
    .io_downs_1_d_payload_param   (ramBridge_up_bus_d_payload_param[2:0]       ), //i
    .io_downs_1_d_payload_source  (ramBridge_up_bus_d_payload_source[2:0]      ), //i
    .io_downs_1_d_payload_size    (ramBridge_up_bus_d_payload_size[2:0]        ), //i
    .io_downs_1_d_payload_denied  (ramBridge_up_bus_d_payload_denied           ), //i
    .io_downs_1_d_payload_data    (ramBridge_up_bus_d_payload_data[63:0]       ), //i
    .io_downs_1_d_payload_corrupt (ramBridge_up_bus_d_payload_corrupt          ), //i
    .clk_cpu                      (board_ctrl_clk_cpu                          ), //i
    .reset_cpu                    (board_ctrl_reset_cpu                        )  //i
  );
  Apb3Bridge toApb_logic_bridge (
    .io_up_a_valid           (toApb_up_bus_a_valid                          ), //i
    .io_up_a_ready           (toApb_logic_bridge_io_up_a_ready              ), //o
    .io_up_a_payload_opcode  (toApb_up_bus_a_payload_opcode[2:0]            ), //i
    .io_up_a_payload_param   (toApb_up_bus_a_payload_param[2:0]             ), //i
    .io_up_a_payload_source  (toApb_up_bus_a_payload_source[2:0]            ), //i
    .io_up_a_payload_address (toApb_up_bus_a_payload_address[26:0]          ), //i
    .io_up_a_payload_size    (toApb_up_bus_a_payload_size[2:0]              ), //i
    .io_up_a_payload_mask    (toApb_up_bus_a_payload_mask[3:0]              ), //i
    .io_up_a_payload_data    (toApb_up_bus_a_payload_data[31:0]             ), //i
    .io_up_a_payload_corrupt (toApb_up_bus_a_payload_corrupt                ), //i
    .io_up_d_valid           (toApb_logic_bridge_io_up_d_valid              ), //o
    .io_up_d_ready           (toApb_up_bus_d_ready                          ), //i
    .io_up_d_payload_opcode  (toApb_logic_bridge_io_up_d_payload_opcode[2:0]), //o
    .io_up_d_payload_param   (toApb_logic_bridge_io_up_d_payload_param[2:0] ), //o
    .io_up_d_payload_source  (toApb_logic_bridge_io_up_d_payload_source[2:0]), //o
    .io_up_d_payload_size    (toApb_logic_bridge_io_up_d_payload_size[2:0]  ), //o
    .io_up_d_payload_denied  (toApb_logic_bridge_io_up_d_payload_denied     ), //o
    .io_up_d_payload_data    (toApb_logic_bridge_io_up_d_payload_data[31:0] ), //o
    .io_up_d_payload_corrupt (toApb_logic_bridge_io_up_d_payload_corrupt    ), //o
    .io_down_PADDR           (toApb_logic_bridge_io_down_PADDR[26:0]        ), //o
    .io_down_PSEL            (toApb_logic_bridge_io_down_PSEL               ), //o
    .io_down_PENABLE         (toApb_logic_bridge_io_down_PENABLE            ), //o
    .io_down_PREADY          (toApb_down_PREADY                             ), //i
    .io_down_PWRITE          (toApb_logic_bridge_io_down_PWRITE             ), //o
    .io_down_PWDATA          (toApb_logic_bridge_io_down_PWDATA[31:0]       ), //o
    .io_down_PRDATA          (toApb_down_PRDATA[31:0]                       ), //i
    .io_down_PSLVERROR       (toApb_down_PSLVERROR                          ), //i
    .clk_cpu                 (board_ctrl_clk_cpu                            ), //i
    .reset_cpu               (board_ctrl_reset_cpu                          )  //i
  );
  Ram internalRam_thread_logic (
    .io_up_a_valid           (internalRam_up_bus_a_valid                          ), //i
    .io_up_a_ready           (internalRam_thread_logic_io_up_a_ready              ), //o
    .io_up_a_payload_opcode  (internalRam_up_bus_a_payload_opcode[2:0]            ), //i
    .io_up_a_payload_param   (internalRam_up_bus_a_payload_param[2:0]             ), //i
    .io_up_a_payload_source  (internalRam_up_bus_a_payload_source[2:0]            ), //i
    .io_up_a_payload_address (internalRam_up_bus_a_payload_address[13:0]          ), //i
    .io_up_a_payload_size    (internalRam_up_bus_a_payload_size[2:0]              ), //i
    .io_up_a_payload_mask    (internalRam_up_bus_a_payload_mask[3:0]              ), //i
    .io_up_a_payload_data    (internalRam_up_bus_a_payload_data[31:0]             ), //i
    .io_up_a_payload_corrupt (internalRam_up_bus_a_payload_corrupt                ), //i
    .io_up_d_valid           (internalRam_thread_logic_io_up_d_valid              ), //o
    .io_up_d_ready           (internalRam_up_bus_d_ready                          ), //i
    .io_up_d_payload_opcode  (internalRam_thread_logic_io_up_d_payload_opcode[2:0]), //o
    .io_up_d_payload_param   (internalRam_thread_logic_io_up_d_payload_param[2:0] ), //o
    .io_up_d_payload_source  (internalRam_thread_logic_io_up_d_payload_source[2:0]), //o
    .io_up_d_payload_size    (internalRam_thread_logic_io_up_d_payload_size[2:0]  ), //o
    .io_up_d_payload_denied  (internalRam_thread_logic_io_up_d_payload_denied     ), //o
    .io_up_d_payload_data    (internalRam_thread_logic_io_up_d_payload_data[31:0] ), //o
    .io_up_d_payload_corrupt (internalRam_thread_logic_io_up_d_payload_corrupt    ), //o
    .clk_cpu                 (board_ctrl_clk_cpu                                  ), //i
    .reset_cpu               (board_ctrl_reset_cpu                                )  //i
  );
  WidthAdapter_1 widthAdapter_3 (
    .io_up_a_valid             (decoder_2_io_downs_0_a_valid                  ), //i
    .io_up_a_ready             (widthAdapter_3_io_up_a_ready                  ), //o
    .io_up_a_payload_opcode    (_zz_io_up_a_payload_opcode_8[2:0]             ), //i
    .io_up_a_payload_param     (decoder_2_io_downs_0_a_payload_param[2:0]     ), //i
    .io_up_a_payload_source    (decoder_2_io_downs_0_a_payload_source[2:0]    ), //i
    .io_up_a_payload_address   (decoder_2_io_downs_0_a_payload_address[30:0]  ), //i
    .io_up_a_payload_size      (decoder_2_io_downs_0_a_payload_size[2:0]      ), //i
    .io_up_a_payload_mask      (decoder_2_io_downs_0_a_payload_mask[7:0]      ), //i
    .io_up_a_payload_data      (decoder_2_io_downs_0_a_payload_data[63:0]     ), //i
    .io_up_a_payload_corrupt   (decoder_2_io_downs_0_a_payload_corrupt        ), //i
    .io_up_d_valid             (widthAdapter_3_io_up_d_valid                  ), //o
    .io_up_d_ready             (decoder_2_io_downs_0_d_ready                  ), //i
    .io_up_d_payload_opcode    (widthAdapter_3_io_up_d_payload_opcode[2:0]    ), //o
    .io_up_d_payload_param     (widthAdapter_3_io_up_d_payload_param[2:0]     ), //o
    .io_up_d_payload_source    (widthAdapter_3_io_up_d_payload_source[2:0]    ), //o
    .io_up_d_payload_size      (widthAdapter_3_io_up_d_payload_size[2:0]      ), //o
    .io_up_d_payload_denied    (widthAdapter_3_io_up_d_payload_denied         ), //o
    .io_up_d_payload_data      (widthAdapter_3_io_up_d_payload_data[63:0]     ), //o
    .io_up_d_payload_corrupt   (widthAdapter_3_io_up_d_payload_corrupt        ), //o
    .io_down_a_valid           (widthAdapter_3_io_down_a_valid                ), //o
    .io_down_a_ready           (decoder_3_io_up_a_ready                       ), //i
    .io_down_a_payload_opcode  (widthAdapter_3_io_down_a_payload_opcode[2:0]  ), //o
    .io_down_a_payload_param   (widthAdapter_3_io_down_a_payload_param[2:0]   ), //o
    .io_down_a_payload_source  (widthAdapter_3_io_down_a_payload_source[2:0]  ), //o
    .io_down_a_payload_address (widthAdapter_3_io_down_a_payload_address[30:0]), //o
    .io_down_a_payload_size    (widthAdapter_3_io_down_a_payload_size[2:0]    ), //o
    .io_down_a_payload_mask    (widthAdapter_3_io_down_a_payload_mask[3:0]    ), //o
    .io_down_a_payload_data    (widthAdapter_3_io_down_a_payload_data[31:0]   ), //o
    .io_down_a_payload_corrupt (widthAdapter_3_io_down_a_payload_corrupt      ), //o
    .io_down_d_valid           (decoder_3_io_up_d_valid                       ), //i
    .io_down_d_ready           (widthAdapter_3_io_down_d_ready                ), //o
    .io_down_d_payload_opcode  (_zz_io_down_d_payload_opcode_3[2:0]           ), //i
    .io_down_d_payload_param   (decoder_3_io_up_d_payload_param[2:0]          ), //i
    .io_down_d_payload_source  (decoder_3_io_up_d_payload_source[2:0]         ), //i
    .io_down_d_payload_size    (decoder_3_io_up_d_payload_size[2:0]           ), //i
    .io_down_d_payload_denied  (decoder_3_io_up_d_payload_denied              ), //i
    .io_down_d_payload_data    (decoder_3_io_up_d_payload_data[31:0]          ), //i
    .io_down_d_payload_corrupt (decoder_3_io_up_d_payload_corrupt             ), //i
    .clk_cpu                   (board_ctrl_clk_cpu                            ), //i
    .reset_cpu                 (board_ctrl_reset_cpu                          )  //i
  );
  Decoder_1 decoder_3 (
    .io_up_a_valid                (widthAdapter_3_io_down_a_valid                ), //i
    .io_up_a_ready                (decoder_3_io_up_a_ready                       ), //o
    .io_up_a_payload_opcode       (_zz_io_up_a_payload_opcode_5[2:0]             ), //i
    .io_up_a_payload_param        (widthAdapter_3_io_down_a_payload_param[2:0]   ), //i
    .io_up_a_payload_source       (widthAdapter_3_io_down_a_payload_source[2:0]  ), //i
    .io_up_a_payload_address      (widthAdapter_3_io_down_a_payload_address[30:0]), //i
    .io_up_a_payload_size         (widthAdapter_3_io_down_a_payload_size[2:0]    ), //i
    .io_up_a_payload_mask         (widthAdapter_3_io_down_a_payload_mask[3:0]    ), //i
    .io_up_a_payload_data         (widthAdapter_3_io_down_a_payload_data[31:0]   ), //i
    .io_up_a_payload_corrupt      (widthAdapter_3_io_down_a_payload_corrupt      ), //i
    .io_up_d_valid                (decoder_3_io_up_d_valid                       ), //o
    .io_up_d_ready                (widthAdapter_3_io_down_d_ready                ), //i
    .io_up_d_payload_opcode       (decoder_3_io_up_d_payload_opcode[2:0]         ), //o
    .io_up_d_payload_param        (decoder_3_io_up_d_payload_param[2:0]          ), //o
    .io_up_d_payload_source       (decoder_3_io_up_d_payload_source[2:0]         ), //o
    .io_up_d_payload_size         (decoder_3_io_up_d_payload_size[2:0]           ), //o
    .io_up_d_payload_denied       (decoder_3_io_up_d_payload_denied              ), //o
    .io_up_d_payload_data         (decoder_3_io_up_d_payload_data[31:0]          ), //o
    .io_up_d_payload_corrupt      (decoder_3_io_up_d_payload_corrupt             ), //o
    .io_downs_0_a_valid           (decoder_3_io_downs_0_a_valid                  ), //o
    .io_downs_0_a_ready           (toApb_up_bus_a_ready                          ), //i
    .io_downs_0_a_payload_opcode  (decoder_3_io_downs_0_a_payload_opcode[2:0]    ), //o
    .io_downs_0_a_payload_param   (decoder_3_io_downs_0_a_payload_param[2:0]     ), //o
    .io_downs_0_a_payload_source  (decoder_3_io_downs_0_a_payload_source[2:0]    ), //o
    .io_downs_0_a_payload_address (decoder_3_io_downs_0_a_payload_address[26:0]  ), //o
    .io_downs_0_a_payload_size    (decoder_3_io_downs_0_a_payload_size[2:0]      ), //o
    .io_downs_0_a_payload_mask    (decoder_3_io_downs_0_a_payload_mask[3:0]      ), //o
    .io_downs_0_a_payload_data    (decoder_3_io_downs_0_a_payload_data[31:0]     ), //o
    .io_downs_0_a_payload_corrupt (decoder_3_io_downs_0_a_payload_corrupt        ), //o
    .io_downs_0_d_valid           (toApb_up_bus_d_valid                          ), //i
    .io_downs_0_d_ready           (decoder_3_io_downs_0_d_ready                  ), //o
    .io_downs_0_d_payload_opcode  (_zz_io_downs_0_d_payload_opcode_2[2:0]        ), //i
    .io_downs_0_d_payload_param   (toApb_up_bus_d_payload_param[2:0]             ), //i
    .io_downs_0_d_payload_source  (toApb_up_bus_d_payload_source[2:0]            ), //i
    .io_downs_0_d_payload_size    (toApb_up_bus_d_payload_size[2:0]              ), //i
    .io_downs_0_d_payload_denied  (toApb_up_bus_d_payload_denied                 ), //i
    .io_downs_0_d_payload_data    (toApb_up_bus_d_payload_data[31:0]             ), //i
    .io_downs_0_d_payload_corrupt (toApb_up_bus_d_payload_corrupt                ), //i
    .io_downs_1_a_valid           (decoder_3_io_downs_1_a_valid                  ), //o
    .io_downs_1_a_ready           (internalRam_up_bus_a_ready                    ), //i
    .io_downs_1_a_payload_opcode  (decoder_3_io_downs_1_a_payload_opcode[2:0]    ), //o
    .io_downs_1_a_payload_param   (decoder_3_io_downs_1_a_payload_param[2:0]     ), //o
    .io_downs_1_a_payload_source  (decoder_3_io_downs_1_a_payload_source[2:0]    ), //o
    .io_downs_1_a_payload_address (decoder_3_io_downs_1_a_payload_address[13:0]  ), //o
    .io_downs_1_a_payload_size    (decoder_3_io_downs_1_a_payload_size[2:0]      ), //o
    .io_downs_1_a_payload_mask    (decoder_3_io_downs_1_a_payload_mask[3:0]      ), //o
    .io_downs_1_a_payload_data    (decoder_3_io_downs_1_a_payload_data[31:0]     ), //o
    .io_downs_1_a_payload_corrupt (decoder_3_io_downs_1_a_payload_corrupt        ), //o
    .io_downs_1_d_valid           (internalRam_up_bus_d_valid                    ), //i
    .io_downs_1_d_ready           (decoder_3_io_downs_1_d_ready                  ), //o
    .io_downs_1_d_payload_opcode  (_zz_io_downs_1_d_payload_opcode_3[2:0]        ), //i
    .io_downs_1_d_payload_param   (internalRam_up_bus_d_payload_param[2:0]       ), //i
    .io_downs_1_d_payload_source  (internalRam_up_bus_d_payload_source[2:0]      ), //i
    .io_downs_1_d_payload_size    (internalRam_up_bus_d_payload_size[2:0]        ), //i
    .io_downs_1_d_payload_denied  (internalRam_up_bus_d_payload_denied           ), //i
    .io_downs_1_d_payload_data    (internalRam_up_bus_d_payload_data[31:0]       ), //i
    .io_downs_1_d_payload_corrupt (internalRam_up_bus_d_payload_corrupt          ), //i
    .clk_cpu                      (board_ctrl_clk_cpu                            ), //i
    .reset_cpu                    (board_ctrl_reset_cpu                          )  //i
  );
  Apb3Decoder_1 toApb_down_decoder (
    .io_input_PADDR      (toApb_down_PADDR[26:0]                   ), //i
    .io_input_PSEL       (toApb_down_PSEL                          ), //i
    .io_input_PENABLE    (toApb_down_PENABLE                       ), //i
    .io_input_PREADY     (toApb_down_decoder_io_input_PREADY       ), //o
    .io_input_PWRITE     (toApb_down_PWRITE                        ), //i
    .io_input_PWDATA     (toApb_down_PWDATA[31:0]                  ), //i
    .io_input_PRDATA     (toApb_down_decoder_io_input_PRDATA[31:0] ), //o
    .io_input_PSLVERROR  (toApb_down_decoder_io_input_PSLVERROR    ), //o
    .io_output_PADDR     (toApb_down_decoder_io_output_PADDR[26:0] ), //o
    .io_output_PSEL      (toApb_down_decoder_io_output_PSEL[3:0]   ), //o
    .io_output_PENABLE   (toApb_down_decoder_io_output_PENABLE     ), //o
    .io_output_PREADY    (apb3Router_3_io_input_PREADY             ), //i
    .io_output_PWRITE    (toApb_down_decoder_io_output_PWRITE      ), //o
    .io_output_PWDATA    (toApb_down_decoder_io_output_PWDATA[31:0]), //o
    .io_output_PRDATA    (apb3Router_3_io_input_PRDATA[31:0]       ), //i
    .io_output_PSLVERROR (apb3Router_3_io_input_PSLVERROR          )  //i
  );
  Apb3Router_1 apb3Router_3 (
    .io_input_PADDR         (toApb_down_decoder_io_output_PADDR[26:0] ), //i
    .io_input_PSEL          (toApb_down_decoder_io_output_PSEL[3:0]   ), //i
    .io_input_PENABLE       (toApb_down_decoder_io_output_PENABLE     ), //i
    .io_input_PREADY        (apb3Router_3_io_input_PREADY             ), //o
    .io_input_PWRITE        (toApb_down_decoder_io_output_PWRITE      ), //i
    .io_input_PWDATA        (toApb_down_decoder_io_output_PWDATA[31:0]), //i
    .io_input_PRDATA        (apb3Router_3_io_input_PRDATA[31:0]       ), //o
    .io_input_PSLVERROR     (apb3Router_3_io_input_PSLVERROR          ), //o
    .io_outputs_0_PADDR     (apb3Router_3_io_outputs_0_PADDR[26:0]    ), //o
    .io_outputs_0_PSEL      (apb3Router_3_io_outputs_0_PSEL           ), //o
    .io_outputs_0_PENABLE   (apb3Router_3_io_outputs_0_PENABLE        ), //o
    .io_outputs_0_PREADY    (peripheral_apb_bridge_input_PREADY       ), //i
    .io_outputs_0_PWRITE    (apb3Router_3_io_outputs_0_PWRITE         ), //o
    .io_outputs_0_PWDATA    (apb3Router_3_io_outputs_0_PWDATA[31:0]   ), //o
    .io_outputs_0_PRDATA    (peripheral_apb_bridge_input_PRDATA[31:0] ), //i
    .io_outputs_0_PSLVERROR (1'b0                                     ), //i
    .io_outputs_1_PADDR     (apb3Router_3_io_outputs_1_PADDR[26:0]    ), //o
    .io_outputs_1_PSEL      (apb3Router_3_io_outputs_1_PSEL           ), //o
    .io_outputs_1_PENABLE   (apb3Router_3_io_outputs_1_PENABLE        ), //o
    .io_outputs_1_PREADY    (board_ctrl_apb_PREADY                    ), //i
    .io_outputs_1_PWRITE    (apb3Router_3_io_outputs_1_PWRITE         ), //o
    .io_outputs_1_PWDATA    (apb3Router_3_io_outputs_1_PWDATA[31:0]   ), //o
    .io_outputs_1_PRDATA    (board_ctrl_apb_PRDATA[31:0]              ), //i
    .io_outputs_1_PSLVERROR (1'b0                                     ), //i
    .io_outputs_2_PADDR     (apb3Router_3_io_outputs_2_PADDR[26:0]    ), //o
    .io_outputs_2_PSEL      (apb3Router_3_io_outputs_2_PSEL           ), //o
    .io_outputs_2_PENABLE   (apb3Router_3_io_outputs_2_PENABLE        ), //o
    .io_outputs_2_PREADY    (video_ctrl_apb_PREADY                    ), //i
    .io_outputs_2_PWRITE    (apb3Router_3_io_outputs_2_PWRITE         ), //o
    .io_outputs_2_PWDATA    (apb3Router_3_io_outputs_2_PWDATA[31:0]   ), //o
    .io_outputs_2_PRDATA    (video_ctrl_apb_PRDATA[31:0]              ), //i
    .io_outputs_2_PSLVERROR (1'b0                                     ), //i
    .io_outputs_3_PADDR     (apb3Router_3_io_outputs_3_PADDR[26:0]    ), //o
    .io_outputs_3_PSEL      (apb3Router_3_io_outputs_3_PSEL           ), //o
    .io_outputs_3_PENABLE   (apb3Router_3_io_outputs_3_PENABLE        ), //o
    .io_outputs_3_PREADY    (plic_apb_PREADY                          ), //i
    .io_outputs_3_PWRITE    (apb3Router_3_io_outputs_3_PWRITE         ), //o
    .io_outputs_3_PWDATA    (apb3Router_3_io_outputs_3_PWDATA[31:0]   ), //o
    .io_outputs_3_PRDATA    (plic_apb_PRDATA[31:0]                    ), //i
    .io_outputs_3_PSLVERROR (1'b0                                     ), //i
    .clk_cpu                (board_ctrl_clk_cpu                       ), //i
    .reset_cpu              (board_ctrl_reset_cpu                     )  //i
  );
  `ifndef SYNTHESIS
  always @(*) begin
    case(_zz_io_ups_0_a_payload_opcode)
      A_PUT_FULL_DATA : _zz_io_ups_0_a_payload_opcode_string = "PUT_FULL_DATA   ";
      A_PUT_PARTIAL_DATA : _zz_io_ups_0_a_payload_opcode_string = "PUT_PARTIAL_DATA";
      A_GET : _zz_io_ups_0_a_payload_opcode_string = "GET             ";
      A_ACQUIRE_BLOCK : _zz_io_ups_0_a_payload_opcode_string = "ACQUIRE_BLOCK   ";
      A_ACQUIRE_PERM : _zz_io_ups_0_a_payload_opcode_string = "ACQUIRE_PERM    ";
      default : _zz_io_ups_0_a_payload_opcode_string = "????????????????";
    endcase
  end
  always @(*) begin
    case(_zz_FetchL1TileLinkPlugin_logic_down_d_payload_opcode)
      D_ACCESS_ACK : _zz_FetchL1TileLinkPlugin_logic_down_d_payload_opcode_string = "ACCESS_ACK     ";
      D_ACCESS_ACK_DATA : _zz_FetchL1TileLinkPlugin_logic_down_d_payload_opcode_string = "ACCESS_ACK_DATA";
      D_GRANT : _zz_FetchL1TileLinkPlugin_logic_down_d_payload_opcode_string = "GRANT          ";
      D_GRANT_DATA : _zz_FetchL1TileLinkPlugin_logic_down_d_payload_opcode_string = "GRANT_DATA     ";
      D_RELEASE_ACK : _zz_FetchL1TileLinkPlugin_logic_down_d_payload_opcode_string = "RELEASE_ACK    ";
      default : _zz_FetchL1TileLinkPlugin_logic_down_d_payload_opcode_string = "???????????????";
    endcase
  end
  always @(*) begin
    case(_zz_io_ups_0_a_payload_opcode_1)
      A_PUT_FULL_DATA : _zz_io_ups_0_a_payload_opcode_1_string = "PUT_FULL_DATA   ";
      A_PUT_PARTIAL_DATA : _zz_io_ups_0_a_payload_opcode_1_string = "PUT_PARTIAL_DATA";
      A_GET : _zz_io_ups_0_a_payload_opcode_1_string = "GET             ";
      A_ACQUIRE_BLOCK : _zz_io_ups_0_a_payload_opcode_1_string = "ACQUIRE_BLOCK   ";
      A_ACQUIRE_PERM : _zz_io_ups_0_a_payload_opcode_1_string = "ACQUIRE_PERM    ";
      default : _zz_io_ups_0_a_payload_opcode_1_string = "????????????????";
    endcase
  end
  always @(*) begin
    case(_zz_FetchL1TileLinkPlugin_logic_down_d_payload_opcode_1)
      D_ACCESS_ACK : _zz_FetchL1TileLinkPlugin_logic_down_d_payload_opcode_1_string = "ACCESS_ACK     ";
      D_ACCESS_ACK_DATA : _zz_FetchL1TileLinkPlugin_logic_down_d_payload_opcode_1_string = "ACCESS_ACK_DATA";
      D_GRANT : _zz_FetchL1TileLinkPlugin_logic_down_d_payload_opcode_1_string = "GRANT          ";
      D_GRANT_DATA : _zz_FetchL1TileLinkPlugin_logic_down_d_payload_opcode_1_string = "GRANT_DATA     ";
      D_RELEASE_ACK : _zz_FetchL1TileLinkPlugin_logic_down_d_payload_opcode_1_string = "RELEASE_ACK    ";
      default : _zz_FetchL1TileLinkPlugin_logic_down_d_payload_opcode_1_string = "???????????????";
    endcase
  end
  always @(*) begin
    case(_zz_io_ups_0_a_payload_opcode_2)
      A_PUT_FULL_DATA : _zz_io_ups_0_a_payload_opcode_2_string = "PUT_FULL_DATA   ";
      A_PUT_PARTIAL_DATA : _zz_io_ups_0_a_payload_opcode_2_string = "PUT_PARTIAL_DATA";
      A_GET : _zz_io_ups_0_a_payload_opcode_2_string = "GET             ";
      A_ACQUIRE_BLOCK : _zz_io_ups_0_a_payload_opcode_2_string = "ACQUIRE_BLOCK   ";
      A_ACQUIRE_PERM : _zz_io_ups_0_a_payload_opcode_2_string = "ACQUIRE_PERM    ";
      default : _zz_io_ups_0_a_payload_opcode_2_string = "????????????????";
    endcase
  end
  always @(*) begin
    case(_zz_io_ups_0_a_payload_opcode_3)
      A_PUT_FULL_DATA : _zz_io_ups_0_a_payload_opcode_3_string = "PUT_FULL_DATA   ";
      A_PUT_PARTIAL_DATA : _zz_io_ups_0_a_payload_opcode_3_string = "PUT_PARTIAL_DATA";
      A_GET : _zz_io_ups_0_a_payload_opcode_3_string = "GET             ";
      A_ACQUIRE_BLOCK : _zz_io_ups_0_a_payload_opcode_3_string = "ACQUIRE_BLOCK   ";
      A_ACQUIRE_PERM : _zz_io_ups_0_a_payload_opcode_3_string = "ACQUIRE_PERM    ";
      default : _zz_io_ups_0_a_payload_opcode_3_string = "????????????????";
    endcase
  end
  always @(*) begin
    case(_zz_io_ups_0_a_payload_opcode_4)
      A_PUT_FULL_DATA : _zz_io_ups_0_a_payload_opcode_4_string = "PUT_FULL_DATA   ";
      A_PUT_PARTIAL_DATA : _zz_io_ups_0_a_payload_opcode_4_string = "PUT_PARTIAL_DATA";
      A_GET : _zz_io_ups_0_a_payload_opcode_4_string = "GET             ";
      A_ACQUIRE_BLOCK : _zz_io_ups_0_a_payload_opcode_4_string = "ACQUIRE_BLOCK   ";
      A_ACQUIRE_PERM : _zz_io_ups_0_a_payload_opcode_4_string = "ACQUIRE_PERM    ";
      default : _zz_io_ups_0_a_payload_opcode_4_string = "????????????????";
    endcase
  end
  always @(*) begin
    case(_zz_io_ups_0_a_payload_opcode_5)
      A_PUT_FULL_DATA : _zz_io_ups_0_a_payload_opcode_5_string = "PUT_FULL_DATA   ";
      A_PUT_PARTIAL_DATA : _zz_io_ups_0_a_payload_opcode_5_string = "PUT_PARTIAL_DATA";
      A_GET : _zz_io_ups_0_a_payload_opcode_5_string = "GET             ";
      A_ACQUIRE_BLOCK : _zz_io_ups_0_a_payload_opcode_5_string = "ACQUIRE_BLOCK   ";
      A_ACQUIRE_PERM : _zz_io_ups_0_a_payload_opcode_5_string = "ACQUIRE_PERM    ";
      default : _zz_io_ups_0_a_payload_opcode_5_string = "????????????????";
    endcase
  end
  always @(*) begin
    case(_zz_FetchL1TileLinkPlugin_logic_down_d_payload_opcode_2)
      D_ACCESS_ACK : _zz_FetchL1TileLinkPlugin_logic_down_d_payload_opcode_2_string = "ACCESS_ACK     ";
      D_ACCESS_ACK_DATA : _zz_FetchL1TileLinkPlugin_logic_down_d_payload_opcode_2_string = "ACCESS_ACK_DATA";
      D_GRANT : _zz_FetchL1TileLinkPlugin_logic_down_d_payload_opcode_2_string = "GRANT          ";
      D_GRANT_DATA : _zz_FetchL1TileLinkPlugin_logic_down_d_payload_opcode_2_string = "GRANT_DATA     ";
      D_RELEASE_ACK : _zz_FetchL1TileLinkPlugin_logic_down_d_payload_opcode_2_string = "RELEASE_ACK    ";
      default : _zz_FetchL1TileLinkPlugin_logic_down_d_payload_opcode_2_string = "???????????????";
    endcase
  end
  always @(*) begin
    case(_zz_FetchL1TileLinkPlugin_logic_down_d_payload_opcode_3)
      D_ACCESS_ACK : _zz_FetchL1TileLinkPlugin_logic_down_d_payload_opcode_3_string = "ACCESS_ACK     ";
      D_ACCESS_ACK_DATA : _zz_FetchL1TileLinkPlugin_logic_down_d_payload_opcode_3_string = "ACCESS_ACK_DATA";
      D_GRANT : _zz_FetchL1TileLinkPlugin_logic_down_d_payload_opcode_3_string = "GRANT          ";
      D_GRANT_DATA : _zz_FetchL1TileLinkPlugin_logic_down_d_payload_opcode_3_string = "GRANT_DATA     ";
      D_RELEASE_ACK : _zz_FetchL1TileLinkPlugin_logic_down_d_payload_opcode_3_string = "RELEASE_ACK    ";
      default : _zz_FetchL1TileLinkPlugin_logic_down_d_payload_opcode_3_string = "???????????????";
    endcase
  end
  always @(*) begin
    case(_zz_io_up_a_payload_opcode)
      A_PUT_FULL_DATA : _zz_io_up_a_payload_opcode_string = "PUT_FULL_DATA   ";
      A_PUT_PARTIAL_DATA : _zz_io_up_a_payload_opcode_string = "PUT_PARTIAL_DATA";
      A_GET : _zz_io_up_a_payload_opcode_string = "GET             ";
      A_ACQUIRE_BLOCK : _zz_io_up_a_payload_opcode_string = "ACQUIRE_BLOCK   ";
      A_ACQUIRE_PERM : _zz_io_up_a_payload_opcode_string = "ACQUIRE_PERM    ";
      default : _zz_io_up_a_payload_opcode_string = "????????????????";
    endcase
  end
  always @(*) begin
    case(_zz_LsuTileLinkPlugin_logic_bridge_down_d_payload_opcode)
      D_ACCESS_ACK : _zz_LsuTileLinkPlugin_logic_bridge_down_d_payload_opcode_string = "ACCESS_ACK     ";
      D_ACCESS_ACK_DATA : _zz_LsuTileLinkPlugin_logic_bridge_down_d_payload_opcode_string = "ACCESS_ACK_DATA";
      D_GRANT : _zz_LsuTileLinkPlugin_logic_bridge_down_d_payload_opcode_string = "GRANT          ";
      D_GRANT_DATA : _zz_LsuTileLinkPlugin_logic_bridge_down_d_payload_opcode_string = "GRANT_DATA     ";
      D_RELEASE_ACK : _zz_LsuTileLinkPlugin_logic_bridge_down_d_payload_opcode_string = "RELEASE_ACK    ";
      default : _zz_LsuTileLinkPlugin_logic_bridge_down_d_payload_opcode_string = "???????????????";
    endcase
  end
  always @(*) begin
    case(_zz_io_up_a_payload_opcode_1)
      A_PUT_FULL_DATA : _zz_io_up_a_payload_opcode_1_string = "PUT_FULL_DATA   ";
      A_PUT_PARTIAL_DATA : _zz_io_up_a_payload_opcode_1_string = "PUT_PARTIAL_DATA";
      A_GET : _zz_io_up_a_payload_opcode_1_string = "GET             ";
      A_ACQUIRE_BLOCK : _zz_io_up_a_payload_opcode_1_string = "ACQUIRE_BLOCK   ";
      A_ACQUIRE_PERM : _zz_io_up_a_payload_opcode_1_string = "ACQUIRE_PERM    ";
      default : _zz_io_up_a_payload_opcode_1_string = "????????????????";
    endcase
  end
  always @(*) begin
    case(_zz_LsuTileLinkPlugin_logic_bridge_down_d_payload_opcode_1)
      D_ACCESS_ACK : _zz_LsuTileLinkPlugin_logic_bridge_down_d_payload_opcode_1_string = "ACCESS_ACK     ";
      D_ACCESS_ACK_DATA : _zz_LsuTileLinkPlugin_logic_bridge_down_d_payload_opcode_1_string = "ACCESS_ACK_DATA";
      D_GRANT : _zz_LsuTileLinkPlugin_logic_bridge_down_d_payload_opcode_1_string = "GRANT          ";
      D_GRANT_DATA : _zz_LsuTileLinkPlugin_logic_bridge_down_d_payload_opcode_1_string = "GRANT_DATA     ";
      D_RELEASE_ACK : _zz_LsuTileLinkPlugin_logic_bridge_down_d_payload_opcode_1_string = "RELEASE_ACK    ";
      default : _zz_LsuTileLinkPlugin_logic_bridge_down_d_payload_opcode_1_string = "???????????????";
    endcase
  end
  always @(*) begin
    case(_zz_io_up_a_payload_opcode_2)
      A_PUT_FULL_DATA : _zz_io_up_a_payload_opcode_2_string = "PUT_FULL_DATA   ";
      A_PUT_PARTIAL_DATA : _zz_io_up_a_payload_opcode_2_string = "PUT_PARTIAL_DATA";
      A_GET : _zz_io_up_a_payload_opcode_2_string = "GET             ";
      A_ACQUIRE_BLOCK : _zz_io_up_a_payload_opcode_2_string = "ACQUIRE_BLOCK   ";
      A_ACQUIRE_PERM : _zz_io_up_a_payload_opcode_2_string = "ACQUIRE_PERM    ";
      default : _zz_io_up_a_payload_opcode_2_string = "????????????????";
    endcase
  end
  always @(*) begin
    case(_zz_io_up_a_payload_opcode_3)
      A_PUT_FULL_DATA : _zz_io_up_a_payload_opcode_3_string = "PUT_FULL_DATA   ";
      A_PUT_PARTIAL_DATA : _zz_io_up_a_payload_opcode_3_string = "PUT_PARTIAL_DATA";
      A_GET : _zz_io_up_a_payload_opcode_3_string = "GET             ";
      A_ACQUIRE_BLOCK : _zz_io_up_a_payload_opcode_3_string = "ACQUIRE_BLOCK   ";
      A_ACQUIRE_PERM : _zz_io_up_a_payload_opcode_3_string = "ACQUIRE_PERM    ";
      default : _zz_io_up_a_payload_opcode_3_string = "????????????????";
    endcase
  end
  always @(*) begin
    case(_zz_LsuTileLinkPlugin_logic_bridge_down_d_payload_opcode_2)
      D_ACCESS_ACK : _zz_LsuTileLinkPlugin_logic_bridge_down_d_payload_opcode_2_string = "ACCESS_ACK     ";
      D_ACCESS_ACK_DATA : _zz_LsuTileLinkPlugin_logic_bridge_down_d_payload_opcode_2_string = "ACCESS_ACK_DATA";
      D_GRANT : _zz_LsuTileLinkPlugin_logic_bridge_down_d_payload_opcode_2_string = "GRANT          ";
      D_GRANT_DATA : _zz_LsuTileLinkPlugin_logic_bridge_down_d_payload_opcode_2_string = "GRANT_DATA     ";
      D_RELEASE_ACK : _zz_LsuTileLinkPlugin_logic_bridge_down_d_payload_opcode_2_string = "RELEASE_ACK    ";
      default : _zz_LsuTileLinkPlugin_logic_bridge_down_d_payload_opcode_2_string = "???????????????";
    endcase
  end
  always @(*) begin
    case(_zz_LsuTileLinkPlugin_logic_bridge_down_d_payload_opcode_3)
      D_ACCESS_ACK : _zz_LsuTileLinkPlugin_logic_bridge_down_d_payload_opcode_3_string = "ACCESS_ACK     ";
      D_ACCESS_ACK_DATA : _zz_LsuTileLinkPlugin_logic_bridge_down_d_payload_opcode_3_string = "ACCESS_ACK_DATA";
      D_GRANT : _zz_LsuTileLinkPlugin_logic_bridge_down_d_payload_opcode_3_string = "GRANT          ";
      D_GRANT_DATA : _zz_LsuTileLinkPlugin_logic_bridge_down_d_payload_opcode_3_string = "GRANT_DATA     ";
      D_RELEASE_ACK : _zz_LsuTileLinkPlugin_logic_bridge_down_d_payload_opcode_3_string = "RELEASE_ACK    ";
      default : _zz_LsuTileLinkPlugin_logic_bridge_down_d_payload_opcode_3_string = "???????????????";
    endcase
  end
  always @(*) begin
    case(_zz_io_ups_2_a_payload_opcode)
      A_PUT_FULL_DATA : _zz_io_ups_2_a_payload_opcode_string = "PUT_FULL_DATA   ";
      A_PUT_PARTIAL_DATA : _zz_io_ups_2_a_payload_opcode_string = "PUT_PARTIAL_DATA";
      A_GET : _zz_io_ups_2_a_payload_opcode_string = "GET             ";
      A_ACQUIRE_BLOCK : _zz_io_ups_2_a_payload_opcode_string = "ACQUIRE_BLOCK   ";
      A_ACQUIRE_PERM : _zz_io_ups_2_a_payload_opcode_string = "ACQUIRE_PERM    ";
      default : _zz_io_ups_2_a_payload_opcode_string = "????????????????";
    endcase
  end
  always @(*) begin
    case(_zz_LsuL1TileLinkPlugin_logic_down_d_payload_opcode)
      D_ACCESS_ACK : _zz_LsuL1TileLinkPlugin_logic_down_d_payload_opcode_string = "ACCESS_ACK     ";
      D_ACCESS_ACK_DATA : _zz_LsuL1TileLinkPlugin_logic_down_d_payload_opcode_string = "ACCESS_ACK_DATA";
      D_GRANT : _zz_LsuL1TileLinkPlugin_logic_down_d_payload_opcode_string = "GRANT          ";
      D_GRANT_DATA : _zz_LsuL1TileLinkPlugin_logic_down_d_payload_opcode_string = "GRANT_DATA     ";
      D_RELEASE_ACK : _zz_LsuL1TileLinkPlugin_logic_down_d_payload_opcode_string = "RELEASE_ACK    ";
      default : _zz_LsuL1TileLinkPlugin_logic_down_d_payload_opcode_string = "???????????????";
    endcase
  end
  always @(*) begin
    case(_zz_io_ups_2_a_payload_opcode_1)
      A_PUT_FULL_DATA : _zz_io_ups_2_a_payload_opcode_1_string = "PUT_FULL_DATA   ";
      A_PUT_PARTIAL_DATA : _zz_io_ups_2_a_payload_opcode_1_string = "PUT_PARTIAL_DATA";
      A_GET : _zz_io_ups_2_a_payload_opcode_1_string = "GET             ";
      A_ACQUIRE_BLOCK : _zz_io_ups_2_a_payload_opcode_1_string = "ACQUIRE_BLOCK   ";
      A_ACQUIRE_PERM : _zz_io_ups_2_a_payload_opcode_1_string = "ACQUIRE_PERM    ";
      default : _zz_io_ups_2_a_payload_opcode_1_string = "????????????????";
    endcase
  end
  always @(*) begin
    case(_zz_LsuL1TileLinkPlugin_logic_down_d_payload_opcode_1)
      D_ACCESS_ACK : _zz_LsuL1TileLinkPlugin_logic_down_d_payload_opcode_1_string = "ACCESS_ACK     ";
      D_ACCESS_ACK_DATA : _zz_LsuL1TileLinkPlugin_logic_down_d_payload_opcode_1_string = "ACCESS_ACK_DATA";
      D_GRANT : _zz_LsuL1TileLinkPlugin_logic_down_d_payload_opcode_1_string = "GRANT          ";
      D_GRANT_DATA : _zz_LsuL1TileLinkPlugin_logic_down_d_payload_opcode_1_string = "GRANT_DATA     ";
      D_RELEASE_ACK : _zz_LsuL1TileLinkPlugin_logic_down_d_payload_opcode_1_string = "RELEASE_ACK    ";
      default : _zz_LsuL1TileLinkPlugin_logic_down_d_payload_opcode_1_string = "???????????????";
    endcase
  end
  always @(*) begin
    case(_zz_io_ups_2_a_payload_opcode_2)
      A_PUT_FULL_DATA : _zz_io_ups_2_a_payload_opcode_2_string = "PUT_FULL_DATA   ";
      A_PUT_PARTIAL_DATA : _zz_io_ups_2_a_payload_opcode_2_string = "PUT_PARTIAL_DATA";
      A_GET : _zz_io_ups_2_a_payload_opcode_2_string = "GET             ";
      A_ACQUIRE_BLOCK : _zz_io_ups_2_a_payload_opcode_2_string = "ACQUIRE_BLOCK   ";
      A_ACQUIRE_PERM : _zz_io_ups_2_a_payload_opcode_2_string = "ACQUIRE_PERM    ";
      default : _zz_io_ups_2_a_payload_opcode_2_string = "????????????????";
    endcase
  end
  always @(*) begin
    case(_zz_io_ups_2_a_payload_opcode_3)
      A_PUT_FULL_DATA : _zz_io_ups_2_a_payload_opcode_3_string = "PUT_FULL_DATA   ";
      A_PUT_PARTIAL_DATA : _zz_io_ups_2_a_payload_opcode_3_string = "PUT_PARTIAL_DATA";
      A_GET : _zz_io_ups_2_a_payload_opcode_3_string = "GET             ";
      A_ACQUIRE_BLOCK : _zz_io_ups_2_a_payload_opcode_3_string = "ACQUIRE_BLOCK   ";
      A_ACQUIRE_PERM : _zz_io_ups_2_a_payload_opcode_3_string = "ACQUIRE_PERM    ";
      default : _zz_io_ups_2_a_payload_opcode_3_string = "????????????????";
    endcase
  end
  always @(*) begin
    case(_zz_LsuL1TileLinkPlugin_logic_down_d_payload_opcode_2)
      D_ACCESS_ACK : _zz_LsuL1TileLinkPlugin_logic_down_d_payload_opcode_2_string = "ACCESS_ACK     ";
      D_ACCESS_ACK_DATA : _zz_LsuL1TileLinkPlugin_logic_down_d_payload_opcode_2_string = "ACCESS_ACK_DATA";
      D_GRANT : _zz_LsuL1TileLinkPlugin_logic_down_d_payload_opcode_2_string = "GRANT          ";
      D_GRANT_DATA : _zz_LsuL1TileLinkPlugin_logic_down_d_payload_opcode_2_string = "GRANT_DATA     ";
      D_RELEASE_ACK : _zz_LsuL1TileLinkPlugin_logic_down_d_payload_opcode_2_string = "RELEASE_ACK    ";
      default : _zz_LsuL1TileLinkPlugin_logic_down_d_payload_opcode_2_string = "???????????????";
    endcase
  end
  always @(*) begin
    case(_zz_LsuL1TileLinkPlugin_logic_down_d_payload_opcode_3)
      D_ACCESS_ACK : _zz_LsuL1TileLinkPlugin_logic_down_d_payload_opcode_3_string = "ACCESS_ACK     ";
      D_ACCESS_ACK_DATA : _zz_LsuL1TileLinkPlugin_logic_down_d_payload_opcode_3_string = "ACCESS_ACK_DATA";
      D_GRANT : _zz_LsuL1TileLinkPlugin_logic_down_d_payload_opcode_3_string = "GRANT          ";
      D_GRANT_DATA : _zz_LsuL1TileLinkPlugin_logic_down_d_payload_opcode_3_string = "GRANT_DATA     ";
      D_RELEASE_ACK : _zz_LsuL1TileLinkPlugin_logic_down_d_payload_opcode_3_string = "RELEASE_ACK    ";
      default : _zz_LsuL1TileLinkPlugin_logic_down_d_payload_opcode_3_string = "???????????????";
    endcase
  end
  always @(*) begin
    case(_zz_io_up_a_payload_opcode_4)
      A_PUT_FULL_DATA : _zz_io_up_a_payload_opcode_4_string = "PUT_FULL_DATA   ";
      A_PUT_PARTIAL_DATA : _zz_io_up_a_payload_opcode_4_string = "PUT_PARTIAL_DATA";
      A_GET : _zz_io_up_a_payload_opcode_4_string = "GET             ";
      A_ACQUIRE_BLOCK : _zz_io_up_a_payload_opcode_4_string = "ACQUIRE_BLOCK   ";
      A_ACQUIRE_PERM : _zz_io_up_a_payload_opcode_4_string = "ACQUIRE_PERM    ";
      default : _zz_io_up_a_payload_opcode_4_string = "????????????????";
    endcase
  end
  always @(*) begin
    case(_zz_io_down_d_payload_opcode)
      D_ACCESS_ACK : _zz_io_down_d_payload_opcode_string = "ACCESS_ACK     ";
      D_ACCESS_ACK_DATA : _zz_io_down_d_payload_opcode_string = "ACCESS_ACK_DATA";
      D_GRANT : _zz_io_down_d_payload_opcode_string = "GRANT          ";
      D_GRANT_DATA : _zz_io_down_d_payload_opcode_string = "GRANT_DATA     ";
      D_RELEASE_ACK : _zz_io_down_d_payload_opcode_string = "RELEASE_ACK    ";
      default : _zz_io_down_d_payload_opcode_string = "???????????????";
    endcase
  end
  always @(*) begin
    case(_zz_io_ups_0_a_payload_opcode_6)
      A_PUT_FULL_DATA : _zz_io_ups_0_a_payload_opcode_6_string = "PUT_FULL_DATA   ";
      A_PUT_PARTIAL_DATA : _zz_io_ups_0_a_payload_opcode_6_string = "PUT_PARTIAL_DATA";
      A_GET : _zz_io_ups_0_a_payload_opcode_6_string = "GET             ";
      A_ACQUIRE_BLOCK : _zz_io_ups_0_a_payload_opcode_6_string = "ACQUIRE_BLOCK   ";
      A_ACQUIRE_PERM : _zz_io_ups_0_a_payload_opcode_6_string = "ACQUIRE_PERM    ";
      default : _zz_io_ups_0_a_payload_opcode_6_string = "????????????????";
    endcase
  end
  always @(*) begin
    case(_zz_FetchL1TileLinkPlugin_logic_down_d_payload_opcode_4)
      D_ACCESS_ACK : _zz_FetchL1TileLinkPlugin_logic_down_d_payload_opcode_4_string = "ACCESS_ACK     ";
      D_ACCESS_ACK_DATA : _zz_FetchL1TileLinkPlugin_logic_down_d_payload_opcode_4_string = "ACCESS_ACK_DATA";
      D_GRANT : _zz_FetchL1TileLinkPlugin_logic_down_d_payload_opcode_4_string = "GRANT          ";
      D_GRANT_DATA : _zz_FetchL1TileLinkPlugin_logic_down_d_payload_opcode_4_string = "GRANT_DATA     ";
      D_RELEASE_ACK : _zz_FetchL1TileLinkPlugin_logic_down_d_payload_opcode_4_string = "RELEASE_ACK    ";
      default : _zz_FetchL1TileLinkPlugin_logic_down_d_payload_opcode_4_string = "???????????????";
    endcase
  end
  always @(*) begin
    case(_zz_io_ups_1_a_payload_opcode)
      A_PUT_FULL_DATA : _zz_io_ups_1_a_payload_opcode_string = "PUT_FULL_DATA   ";
      A_PUT_PARTIAL_DATA : _zz_io_ups_1_a_payload_opcode_string = "PUT_PARTIAL_DATA";
      A_GET : _zz_io_ups_1_a_payload_opcode_string = "GET             ";
      A_ACQUIRE_BLOCK : _zz_io_ups_1_a_payload_opcode_string = "ACQUIRE_BLOCK   ";
      A_ACQUIRE_PERM : _zz_io_ups_1_a_payload_opcode_string = "ACQUIRE_PERM    ";
      default : _zz_io_ups_1_a_payload_opcode_string = "????????????????";
    endcase
  end
  always @(*) begin
    case(_zz_io_down_d_payload_opcode_1)
      D_ACCESS_ACK : _zz_io_down_d_payload_opcode_1_string = "ACCESS_ACK     ";
      D_ACCESS_ACK_DATA : _zz_io_down_d_payload_opcode_1_string = "ACCESS_ACK_DATA";
      D_GRANT : _zz_io_down_d_payload_opcode_1_string = "GRANT          ";
      D_GRANT_DATA : _zz_io_down_d_payload_opcode_1_string = "GRANT_DATA     ";
      D_RELEASE_ACK : _zz_io_down_d_payload_opcode_1_string = "RELEASE_ACK    ";
      default : _zz_io_down_d_payload_opcode_1_string = "???????????????";
    endcase
  end
  always @(*) begin
    case(_zz_io_ups_2_a_payload_opcode_4)
      A_PUT_FULL_DATA : _zz_io_ups_2_a_payload_opcode_4_string = "PUT_FULL_DATA   ";
      A_PUT_PARTIAL_DATA : _zz_io_ups_2_a_payload_opcode_4_string = "PUT_PARTIAL_DATA";
      A_GET : _zz_io_ups_2_a_payload_opcode_4_string = "GET             ";
      A_ACQUIRE_BLOCK : _zz_io_ups_2_a_payload_opcode_4_string = "ACQUIRE_BLOCK   ";
      A_ACQUIRE_PERM : _zz_io_ups_2_a_payload_opcode_4_string = "ACQUIRE_PERM    ";
      default : _zz_io_ups_2_a_payload_opcode_4_string = "????????????????";
    endcase
  end
  always @(*) begin
    case(_zz_LsuL1TileLinkPlugin_logic_down_d_payload_opcode_4)
      D_ACCESS_ACK : _zz_LsuL1TileLinkPlugin_logic_down_d_payload_opcode_4_string = "ACCESS_ACK     ";
      D_ACCESS_ACK_DATA : _zz_LsuL1TileLinkPlugin_logic_down_d_payload_opcode_4_string = "ACCESS_ACK_DATA";
      D_GRANT : _zz_LsuL1TileLinkPlugin_logic_down_d_payload_opcode_4_string = "GRANT          ";
      D_GRANT_DATA : _zz_LsuL1TileLinkPlugin_logic_down_d_payload_opcode_4_string = "GRANT_DATA     ";
      D_RELEASE_ACK : _zz_LsuL1TileLinkPlugin_logic_down_d_payload_opcode_4_string = "RELEASE_ACK    ";
      default : _zz_LsuL1TileLinkPlugin_logic_down_d_payload_opcode_4_string = "???????????????";
    endcase
  end
  always @(*) begin
    case(_zz_io_up_a_payload_opcode_5)
      A_PUT_FULL_DATA : _zz_io_up_a_payload_opcode_5_string = "PUT_FULL_DATA   ";
      A_PUT_PARTIAL_DATA : _zz_io_up_a_payload_opcode_5_string = "PUT_PARTIAL_DATA";
      A_GET : _zz_io_up_a_payload_opcode_5_string = "GET             ";
      A_ACQUIRE_BLOCK : _zz_io_up_a_payload_opcode_5_string = "ACQUIRE_BLOCK   ";
      A_ACQUIRE_PERM : _zz_io_up_a_payload_opcode_5_string = "ACQUIRE_PERM    ";
      default : _zz_io_up_a_payload_opcode_5_string = "????????????????";
    endcase
  end
  always @(*) begin
    case(_zz_io_down_d_payload_opcode_2)
      D_ACCESS_ACK : _zz_io_down_d_payload_opcode_2_string = "ACCESS_ACK     ";
      D_ACCESS_ACK_DATA : _zz_io_down_d_payload_opcode_2_string = "ACCESS_ACK_DATA";
      D_GRANT : _zz_io_down_d_payload_opcode_2_string = "GRANT          ";
      D_GRANT_DATA : _zz_io_down_d_payload_opcode_2_string = "GRANT_DATA     ";
      D_RELEASE_ACK : _zz_io_down_d_payload_opcode_2_string = "RELEASE_ACK    ";
      default : _zz_io_down_d_payload_opcode_2_string = "???????????????";
    endcase
  end
  always @(*) begin
    case(_zz_io_up_a_payload_opcode_6)
      A_PUT_FULL_DATA : _zz_io_up_a_payload_opcode_6_string = "PUT_FULL_DATA   ";
      A_PUT_PARTIAL_DATA : _zz_io_up_a_payload_opcode_6_string = "PUT_PARTIAL_DATA";
      A_GET : _zz_io_up_a_payload_opcode_6_string = "GET             ";
      A_ACQUIRE_BLOCK : _zz_io_up_a_payload_opcode_6_string = "ACQUIRE_BLOCK   ";
      A_ACQUIRE_PERM : _zz_io_up_a_payload_opcode_6_string = "ACQUIRE_PERM    ";
      default : _zz_io_up_a_payload_opcode_6_string = "????????????????";
    endcase
  end
  always @(*) begin
    case(_zz_io_down_d_payload_opcode_3)
      D_ACCESS_ACK : _zz_io_down_d_payload_opcode_3_string = "ACCESS_ACK     ";
      D_ACCESS_ACK_DATA : _zz_io_down_d_payload_opcode_3_string = "ACCESS_ACK_DATA";
      D_GRANT : _zz_io_down_d_payload_opcode_3_string = "GRANT          ";
      D_GRANT_DATA : _zz_io_down_d_payload_opcode_3_string = "GRANT_DATA     ";
      D_RELEASE_ACK : _zz_io_down_d_payload_opcode_3_string = "RELEASE_ACK    ";
      default : _zz_io_down_d_payload_opcode_3_string = "???????????????";
    endcase
  end
  always @(*) begin
    case(ramBridge_up_bus_a_payload_opcode)
      A_PUT_FULL_DATA : ramBridge_up_bus_a_payload_opcode_string = "PUT_FULL_DATA   ";
      A_PUT_PARTIAL_DATA : ramBridge_up_bus_a_payload_opcode_string = "PUT_PARTIAL_DATA";
      A_GET : ramBridge_up_bus_a_payload_opcode_string = "GET             ";
      A_ACQUIRE_BLOCK : ramBridge_up_bus_a_payload_opcode_string = "ACQUIRE_BLOCK   ";
      A_ACQUIRE_PERM : ramBridge_up_bus_a_payload_opcode_string = "ACQUIRE_PERM    ";
      default : ramBridge_up_bus_a_payload_opcode_string = "????????????????";
    endcase
  end
  always @(*) begin
    case(ramBridge_up_bus_d_payload_opcode)
      D_ACCESS_ACK : ramBridge_up_bus_d_payload_opcode_string = "ACCESS_ACK     ";
      D_ACCESS_ACK_DATA : ramBridge_up_bus_d_payload_opcode_string = "ACCESS_ACK_DATA";
      D_GRANT : ramBridge_up_bus_d_payload_opcode_string = "GRANT          ";
      D_GRANT_DATA : ramBridge_up_bus_d_payload_opcode_string = "GRANT_DATA     ";
      D_RELEASE_ACK : ramBridge_up_bus_d_payload_opcode_string = "RELEASE_ACK    ";
      default : ramBridge_up_bus_d_payload_opcode_string = "???????????????";
    endcase
  end
  always @(*) begin
    case(_zz_ramBridge_up_bus_a_payload_opcode)
      A_PUT_FULL_DATA : _zz_ramBridge_up_bus_a_payload_opcode_string = "PUT_FULL_DATA   ";
      A_PUT_PARTIAL_DATA : _zz_ramBridge_up_bus_a_payload_opcode_string = "PUT_PARTIAL_DATA";
      A_GET : _zz_ramBridge_up_bus_a_payload_opcode_string = "GET             ";
      A_ACQUIRE_BLOCK : _zz_ramBridge_up_bus_a_payload_opcode_string = "ACQUIRE_BLOCK   ";
      A_ACQUIRE_PERM : _zz_ramBridge_up_bus_a_payload_opcode_string = "ACQUIRE_PERM    ";
      default : _zz_ramBridge_up_bus_a_payload_opcode_string = "????????????????";
    endcase
  end
  always @(*) begin
    case(_zz_io_downs_1_d_payload_opcode)
      D_ACCESS_ACK : _zz_io_downs_1_d_payload_opcode_string = "ACCESS_ACK     ";
      D_ACCESS_ACK_DATA : _zz_io_downs_1_d_payload_opcode_string = "ACCESS_ACK_DATA";
      D_GRANT : _zz_io_downs_1_d_payload_opcode_string = "GRANT          ";
      D_GRANT_DATA : _zz_io_downs_1_d_payload_opcode_string = "GRANT_DATA     ";
      D_RELEASE_ACK : _zz_io_downs_1_d_payload_opcode_string = "RELEASE_ACK    ";
      default : _zz_io_downs_1_d_payload_opcode_string = "???????????????";
    endcase
  end
  always @(*) begin
    case(_zz_io_ups_0_a_payload_opcode_7)
      A_PUT_FULL_DATA : _zz_io_ups_0_a_payload_opcode_7_string = "PUT_FULL_DATA   ";
      A_PUT_PARTIAL_DATA : _zz_io_ups_0_a_payload_opcode_7_string = "PUT_PARTIAL_DATA";
      A_GET : _zz_io_ups_0_a_payload_opcode_7_string = "GET             ";
      A_ACQUIRE_BLOCK : _zz_io_ups_0_a_payload_opcode_7_string = "ACQUIRE_BLOCK   ";
      A_ACQUIRE_PERM : _zz_io_ups_0_a_payload_opcode_7_string = "ACQUIRE_PERM    ";
      default : _zz_io_ups_0_a_payload_opcode_7_string = "????????????????";
    endcase
  end
  always @(*) begin
    case(_zz_FetchL1TileLinkPlugin_logic_down_d_payload_opcode_5)
      D_ACCESS_ACK : _zz_FetchL1TileLinkPlugin_logic_down_d_payload_opcode_5_string = "ACCESS_ACK     ";
      D_ACCESS_ACK_DATA : _zz_FetchL1TileLinkPlugin_logic_down_d_payload_opcode_5_string = "ACCESS_ACK_DATA";
      D_GRANT : _zz_FetchL1TileLinkPlugin_logic_down_d_payload_opcode_5_string = "GRANT          ";
      D_GRANT_DATA : _zz_FetchL1TileLinkPlugin_logic_down_d_payload_opcode_5_string = "GRANT_DATA     ";
      D_RELEASE_ACK : _zz_FetchL1TileLinkPlugin_logic_down_d_payload_opcode_5_string = "RELEASE_ACK    ";
      default : _zz_FetchL1TileLinkPlugin_logic_down_d_payload_opcode_5_string = "???????????????";
    endcase
  end
  always @(*) begin
    case(_zz_io_up_a_payload_opcode_7)
      A_PUT_FULL_DATA : _zz_io_up_a_payload_opcode_7_string = "PUT_FULL_DATA   ";
      A_PUT_PARTIAL_DATA : _zz_io_up_a_payload_opcode_7_string = "PUT_PARTIAL_DATA";
      A_GET : _zz_io_up_a_payload_opcode_7_string = "GET             ";
      A_ACQUIRE_BLOCK : _zz_io_up_a_payload_opcode_7_string = "ACQUIRE_BLOCK   ";
      A_ACQUIRE_PERM : _zz_io_up_a_payload_opcode_7_string = "ACQUIRE_PERM    ";
      default : _zz_io_up_a_payload_opcode_7_string = "????????????????";
    endcase
  end
  always @(*) begin
    case(_zz_LsuTileLinkPlugin_logic_bridge_down_d_payload_opcode_4)
      D_ACCESS_ACK : _zz_LsuTileLinkPlugin_logic_bridge_down_d_payload_opcode_4_string = "ACCESS_ACK     ";
      D_ACCESS_ACK_DATA : _zz_LsuTileLinkPlugin_logic_bridge_down_d_payload_opcode_4_string = "ACCESS_ACK_DATA";
      D_GRANT : _zz_LsuTileLinkPlugin_logic_bridge_down_d_payload_opcode_4_string = "GRANT          ";
      D_GRANT_DATA : _zz_LsuTileLinkPlugin_logic_bridge_down_d_payload_opcode_4_string = "GRANT_DATA     ";
      D_RELEASE_ACK : _zz_LsuTileLinkPlugin_logic_bridge_down_d_payload_opcode_4_string = "RELEASE_ACK    ";
      default : _zz_LsuTileLinkPlugin_logic_bridge_down_d_payload_opcode_4_string = "???????????????";
    endcase
  end
  always @(*) begin
    case(_zz_io_ups_2_a_payload_opcode_5)
      A_PUT_FULL_DATA : _zz_io_ups_2_a_payload_opcode_5_string = "PUT_FULL_DATA   ";
      A_PUT_PARTIAL_DATA : _zz_io_ups_2_a_payload_opcode_5_string = "PUT_PARTIAL_DATA";
      A_GET : _zz_io_ups_2_a_payload_opcode_5_string = "GET             ";
      A_ACQUIRE_BLOCK : _zz_io_ups_2_a_payload_opcode_5_string = "ACQUIRE_BLOCK   ";
      A_ACQUIRE_PERM : _zz_io_ups_2_a_payload_opcode_5_string = "ACQUIRE_PERM    ";
      default : _zz_io_ups_2_a_payload_opcode_5_string = "????????????????";
    endcase
  end
  always @(*) begin
    case(_zz_LsuL1TileLinkPlugin_logic_down_d_payload_opcode_5)
      D_ACCESS_ACK : _zz_LsuL1TileLinkPlugin_logic_down_d_payload_opcode_5_string = "ACCESS_ACK     ";
      D_ACCESS_ACK_DATA : _zz_LsuL1TileLinkPlugin_logic_down_d_payload_opcode_5_string = "ACCESS_ACK_DATA";
      D_GRANT : _zz_LsuL1TileLinkPlugin_logic_down_d_payload_opcode_5_string = "GRANT          ";
      D_GRANT_DATA : _zz_LsuL1TileLinkPlugin_logic_down_d_payload_opcode_5_string = "GRANT_DATA     ";
      D_RELEASE_ACK : _zz_LsuL1TileLinkPlugin_logic_down_d_payload_opcode_5_string = "RELEASE_ACK    ";
      default : _zz_LsuL1TileLinkPlugin_logic_down_d_payload_opcode_5_string = "???????????????";
    endcase
  end
  always @(*) begin
    case(toApb_up_bus_a_payload_opcode)
      A_PUT_FULL_DATA : toApb_up_bus_a_payload_opcode_string = "PUT_FULL_DATA   ";
      A_PUT_PARTIAL_DATA : toApb_up_bus_a_payload_opcode_string = "PUT_PARTIAL_DATA";
      A_GET : toApb_up_bus_a_payload_opcode_string = "GET             ";
      A_ACQUIRE_BLOCK : toApb_up_bus_a_payload_opcode_string = "ACQUIRE_BLOCK   ";
      A_ACQUIRE_PERM : toApb_up_bus_a_payload_opcode_string = "ACQUIRE_PERM    ";
      default : toApb_up_bus_a_payload_opcode_string = "????????????????";
    endcase
  end
  always @(*) begin
    case(toApb_up_bus_d_payload_opcode)
      D_ACCESS_ACK : toApb_up_bus_d_payload_opcode_string = "ACCESS_ACK     ";
      D_ACCESS_ACK_DATA : toApb_up_bus_d_payload_opcode_string = "ACCESS_ACK_DATA";
      D_GRANT : toApb_up_bus_d_payload_opcode_string = "GRANT          ";
      D_GRANT_DATA : toApb_up_bus_d_payload_opcode_string = "GRANT_DATA     ";
      D_RELEASE_ACK : toApb_up_bus_d_payload_opcode_string = "RELEASE_ACK    ";
      default : toApb_up_bus_d_payload_opcode_string = "???????????????";
    endcase
  end
  always @(*) begin
    case(_zz_toApb_up_bus_a_payload_opcode)
      A_PUT_FULL_DATA : _zz_toApb_up_bus_a_payload_opcode_string = "PUT_FULL_DATA   ";
      A_PUT_PARTIAL_DATA : _zz_toApb_up_bus_a_payload_opcode_string = "PUT_PARTIAL_DATA";
      A_GET : _zz_toApb_up_bus_a_payload_opcode_string = "GET             ";
      A_ACQUIRE_BLOCK : _zz_toApb_up_bus_a_payload_opcode_string = "ACQUIRE_BLOCK   ";
      A_ACQUIRE_PERM : _zz_toApb_up_bus_a_payload_opcode_string = "ACQUIRE_PERM    ";
      default : _zz_toApb_up_bus_a_payload_opcode_string = "????????????????";
    endcase
  end
  always @(*) begin
    case(_zz_io_downs_0_d_payload_opcode)
      D_ACCESS_ACK : _zz_io_downs_0_d_payload_opcode_string = "ACCESS_ACK     ";
      D_ACCESS_ACK_DATA : _zz_io_downs_0_d_payload_opcode_string = "ACCESS_ACK_DATA";
      D_GRANT : _zz_io_downs_0_d_payload_opcode_string = "GRANT          ";
      D_GRANT_DATA : _zz_io_downs_0_d_payload_opcode_string = "GRANT_DATA     ";
      D_RELEASE_ACK : _zz_io_downs_0_d_payload_opcode_string = "RELEASE_ACK    ";
      default : _zz_io_downs_0_d_payload_opcode_string = "???????????????";
    endcase
  end
  always @(*) begin
    case(internalRam_up_bus_a_payload_opcode)
      A_PUT_FULL_DATA : internalRam_up_bus_a_payload_opcode_string = "PUT_FULL_DATA   ";
      A_PUT_PARTIAL_DATA : internalRam_up_bus_a_payload_opcode_string = "PUT_PARTIAL_DATA";
      A_GET : internalRam_up_bus_a_payload_opcode_string = "GET             ";
      A_ACQUIRE_BLOCK : internalRam_up_bus_a_payload_opcode_string = "ACQUIRE_BLOCK   ";
      A_ACQUIRE_PERM : internalRam_up_bus_a_payload_opcode_string = "ACQUIRE_PERM    ";
      default : internalRam_up_bus_a_payload_opcode_string = "????????????????";
    endcase
  end
  always @(*) begin
    case(internalRam_up_bus_d_payload_opcode)
      D_ACCESS_ACK : internalRam_up_bus_d_payload_opcode_string = "ACCESS_ACK     ";
      D_ACCESS_ACK_DATA : internalRam_up_bus_d_payload_opcode_string = "ACCESS_ACK_DATA";
      D_GRANT : internalRam_up_bus_d_payload_opcode_string = "GRANT          ";
      D_GRANT_DATA : internalRam_up_bus_d_payload_opcode_string = "GRANT_DATA     ";
      D_RELEASE_ACK : internalRam_up_bus_d_payload_opcode_string = "RELEASE_ACK    ";
      default : internalRam_up_bus_d_payload_opcode_string = "???????????????";
    endcase
  end
  always @(*) begin
    case(_zz_internalRam_up_bus_a_payload_opcode)
      A_PUT_FULL_DATA : _zz_internalRam_up_bus_a_payload_opcode_string = "PUT_FULL_DATA   ";
      A_PUT_PARTIAL_DATA : _zz_internalRam_up_bus_a_payload_opcode_string = "PUT_PARTIAL_DATA";
      A_GET : _zz_internalRam_up_bus_a_payload_opcode_string = "GET             ";
      A_ACQUIRE_BLOCK : _zz_internalRam_up_bus_a_payload_opcode_string = "ACQUIRE_BLOCK   ";
      A_ACQUIRE_PERM : _zz_internalRam_up_bus_a_payload_opcode_string = "ACQUIRE_PERM    ";
      default : _zz_internalRam_up_bus_a_payload_opcode_string = "????????????????";
    endcase
  end
  always @(*) begin
    case(_zz_io_downs_1_d_payload_opcode_1)
      D_ACCESS_ACK : _zz_io_downs_1_d_payload_opcode_1_string = "ACCESS_ACK     ";
      D_ACCESS_ACK_DATA : _zz_io_downs_1_d_payload_opcode_1_string = "ACCESS_ACK_DATA";
      D_GRANT : _zz_io_downs_1_d_payload_opcode_1_string = "GRANT          ";
      D_GRANT_DATA : _zz_io_downs_1_d_payload_opcode_1_string = "GRANT_DATA     ";
      D_RELEASE_ACK : _zz_io_downs_1_d_payload_opcode_1_string = "RELEASE_ACK    ";
      default : _zz_io_downs_1_d_payload_opcode_1_string = "???????????????";
    endcase
  end
  always @(*) begin
    case(_zz_io_up_a_payload_opcode_8)
      A_PUT_FULL_DATA : _zz_io_up_a_payload_opcode_8_string = "PUT_FULL_DATA   ";
      A_PUT_PARTIAL_DATA : _zz_io_up_a_payload_opcode_8_string = "PUT_PARTIAL_DATA";
      A_GET : _zz_io_up_a_payload_opcode_8_string = "GET             ";
      A_ACQUIRE_BLOCK : _zz_io_up_a_payload_opcode_8_string = "ACQUIRE_BLOCK   ";
      A_ACQUIRE_PERM : _zz_io_up_a_payload_opcode_8_string = "ACQUIRE_PERM    ";
      default : _zz_io_up_a_payload_opcode_8_string = "????????????????";
    endcase
  end
  always @(*) begin
    case(_zz_io_downs_0_d_payload_opcode_1)
      D_ACCESS_ACK : _zz_io_downs_0_d_payload_opcode_1_string = "ACCESS_ACK     ";
      D_ACCESS_ACK_DATA : _zz_io_downs_0_d_payload_opcode_1_string = "ACCESS_ACK_DATA";
      D_GRANT : _zz_io_downs_0_d_payload_opcode_1_string = "GRANT          ";
      D_GRANT_DATA : _zz_io_downs_0_d_payload_opcode_1_string = "GRANT_DATA     ";
      D_RELEASE_ACK : _zz_io_downs_0_d_payload_opcode_1_string = "RELEASE_ACK    ";
      default : _zz_io_downs_0_d_payload_opcode_1_string = "???????????????";
    endcase
  end
  always @(*) begin
    case(_zz_ramBridge_up_bus_a_payload_opcode_1)
      A_PUT_FULL_DATA : _zz_ramBridge_up_bus_a_payload_opcode_1_string = "PUT_FULL_DATA   ";
      A_PUT_PARTIAL_DATA : _zz_ramBridge_up_bus_a_payload_opcode_1_string = "PUT_PARTIAL_DATA";
      A_GET : _zz_ramBridge_up_bus_a_payload_opcode_1_string = "GET             ";
      A_ACQUIRE_BLOCK : _zz_ramBridge_up_bus_a_payload_opcode_1_string = "ACQUIRE_BLOCK   ";
      A_ACQUIRE_PERM : _zz_ramBridge_up_bus_a_payload_opcode_1_string = "ACQUIRE_PERM    ";
      default : _zz_ramBridge_up_bus_a_payload_opcode_1_string = "????????????????";
    endcase
  end
  always @(*) begin
    case(_zz_io_downs_1_d_payload_opcode_2)
      D_ACCESS_ACK : _zz_io_downs_1_d_payload_opcode_2_string = "ACCESS_ACK     ";
      D_ACCESS_ACK_DATA : _zz_io_downs_1_d_payload_opcode_2_string = "ACCESS_ACK_DATA";
      D_GRANT : _zz_io_downs_1_d_payload_opcode_2_string = "GRANT          ";
      D_GRANT_DATA : _zz_io_downs_1_d_payload_opcode_2_string = "GRANT_DATA     ";
      D_RELEASE_ACK : _zz_io_downs_1_d_payload_opcode_2_string = "RELEASE_ACK    ";
      default : _zz_io_downs_1_d_payload_opcode_2_string = "???????????????";
    endcase
  end
  always @(*) begin
    case(_zz_toApb_up_bus_a_payload_opcode_1)
      A_PUT_FULL_DATA : _zz_toApb_up_bus_a_payload_opcode_1_string = "PUT_FULL_DATA   ";
      A_PUT_PARTIAL_DATA : _zz_toApb_up_bus_a_payload_opcode_1_string = "PUT_PARTIAL_DATA";
      A_GET : _zz_toApb_up_bus_a_payload_opcode_1_string = "GET             ";
      A_ACQUIRE_BLOCK : _zz_toApb_up_bus_a_payload_opcode_1_string = "ACQUIRE_BLOCK   ";
      A_ACQUIRE_PERM : _zz_toApb_up_bus_a_payload_opcode_1_string = "ACQUIRE_PERM    ";
      default : _zz_toApb_up_bus_a_payload_opcode_1_string = "????????????????";
    endcase
  end
  always @(*) begin
    case(_zz_io_downs_0_d_payload_opcode_2)
      D_ACCESS_ACK : _zz_io_downs_0_d_payload_opcode_2_string = "ACCESS_ACK     ";
      D_ACCESS_ACK_DATA : _zz_io_downs_0_d_payload_opcode_2_string = "ACCESS_ACK_DATA";
      D_GRANT : _zz_io_downs_0_d_payload_opcode_2_string = "GRANT          ";
      D_GRANT_DATA : _zz_io_downs_0_d_payload_opcode_2_string = "GRANT_DATA     ";
      D_RELEASE_ACK : _zz_io_downs_0_d_payload_opcode_2_string = "RELEASE_ACK    ";
      default : _zz_io_downs_0_d_payload_opcode_2_string = "???????????????";
    endcase
  end
  always @(*) begin
    case(_zz_internalRam_up_bus_a_payload_opcode_1)
      A_PUT_FULL_DATA : _zz_internalRam_up_bus_a_payload_opcode_1_string = "PUT_FULL_DATA   ";
      A_PUT_PARTIAL_DATA : _zz_internalRam_up_bus_a_payload_opcode_1_string = "PUT_PARTIAL_DATA";
      A_GET : _zz_internalRam_up_bus_a_payload_opcode_1_string = "GET             ";
      A_ACQUIRE_BLOCK : _zz_internalRam_up_bus_a_payload_opcode_1_string = "ACQUIRE_BLOCK   ";
      A_ACQUIRE_PERM : _zz_internalRam_up_bus_a_payload_opcode_1_string = "ACQUIRE_PERM    ";
      default : _zz_internalRam_up_bus_a_payload_opcode_1_string = "????????????????";
    endcase
  end
  always @(*) begin
    case(_zz_io_downs_1_d_payload_opcode_3)
      D_ACCESS_ACK : _zz_io_downs_1_d_payload_opcode_3_string = "ACCESS_ACK     ";
      D_ACCESS_ACK_DATA : _zz_io_downs_1_d_payload_opcode_3_string = "ACCESS_ACK_DATA";
      D_GRANT : _zz_io_downs_1_d_payload_opcode_3_string = "GRANT          ";
      D_GRANT_DATA : _zz_io_downs_1_d_payload_opcode_3_string = "GRANT_DATA     ";
      D_RELEASE_ACK : _zz_io_downs_1_d_payload_opcode_3_string = "RELEASE_ACK    ";
      default : _zz_io_downs_1_d_payload_opcode_3_string = "???????????????";
    endcase
  end
  `endif

  assign io_plla_i2c_scl = board_ctrl_plla_i2c_scl;
  assign io_pllb_i2c_scl = board_ctrl_pllb_i2c_scl;
  assign io_leds = board_ctrl_leds;
  assign io_dvi_tmds0p = video_ctrl_dvi_tmds0p;
  assign io_dvi_tmds0m = video_ctrl_dvi_tmds0m;
  assign io_dvi_tmds1p = video_ctrl_dvi_tmds1p;
  assign io_dvi_tmds1m = video_ctrl_dvi_tmds1m;
  assign io_dvi_tmds2p = video_ctrl_dvi_tmds2p;
  assign io_dvi_tmds2m = video_ctrl_dvi_tmds2m;
  assign io_dvi_tmdsCp = video_ctrl_dvi_tmdsCp;
  assign io_dvi_tmdsCm = video_ctrl_dvi_tmdsCm;
  assign io_uart_tx = peripheral_uart_ctrl_uart_tx;
  assign io_audio_shdn = peripheral_audio_ctrl_shdn;
  assign io_audio_i2c_scl = peripheral_audio_ctrl_i2c_scl;
  assign io_sdcard_clk = peripheral_sdcard_ctrl_sdcard_clk;
  assign peripheral_apb_PREADY = peripheral_apb_decoder_io_input_PREADY;
  assign peripheral_apb_PRDATA = peripheral_apb_decoder_io_input_PRDATA;
  assign peripheral_uart_ctrl_apb_PADDR = apb3Router_2_io_outputs_0_PADDR[3:0];
  assign peripheral_audio_ctrl_apb_PADDR = apb3Router_2_io_outputs_1_PADDR[2:0];
  assign peripheral_sdcard_ctrl_apb_PADDR = apb3Router_2_io_outputs_2_PADDR[4:0];
  assign peripheral_usb_ctrl_io_apb_ctrl_PADDR = apb3Router_2_io_outputs_3_PADDR[11:0];
  assign peripheral_usb_ctrl_io_apb_dma_PADDR = apb3Router_2_io_outputs_4_PADDR[11:0];
  assign peripheral_apb_PADDR = peripheral_apb_bridge_output_PADDR;
  assign peripheral_apb_PSEL = peripheral_apb_bridge_output_PSEL;
  assign peripheral_apb_PENABLE = peripheral_apb_bridge_output_PENABLE;
  assign peripheral_apb_PWRITE = peripheral_apb_bridge_output_PWRITE;
  assign peripheral_apb_PWDATA = peripheral_apb_bridge_output_PWDATA;
  assign when_PlicGateway_l21 = (! plic_gateways_0_waitCompletion);
  assign when_PlicGateway_l21_1 = (! plic_gateways_1_waitCompletion);
  assign when_PlicGateway_l21_2 = (! plic_gateways_2_waitCompletion);
  assign plic_target_requests_0_priority = 1'b0;
  assign plic_target_requests_0_id = 2'b00;
  assign plic_target_requests_0_valid = 1'b1;
  assign plic_target_requests_1_priority = plic_gateways_0_priority;
  assign plic_target_requests_1_id = 2'b01;
  assign plic_target_requests_1_valid = (plic_gateways_0_ip && plic_target_ie_0);
  assign plic_target_requests_2_priority = plic_gateways_1_priority;
  assign plic_target_requests_2_id = 2'b10;
  assign plic_target_requests_2_valid = (plic_gateways_1_ip && plic_target_ie_1);
  assign plic_target_requests_3_priority = plic_gateways_2_priority;
  assign plic_target_requests_3_id = 2'b11;
  assign plic_target_requests_3_valid = (plic_gateways_2_ip && plic_target_ie_2);
  assign _zz_plic_target_bestRequest_id = ((! plic_target_requests_1_valid) || (plic_target_requests_0_valid && (plic_target_requests_1_priority <= plic_target_requests_0_priority)));
  assign _zz_plic_target_bestRequest_priority = (_zz_plic_target_bestRequest_id ? plic_target_requests_0_priority : plic_target_requests_1_priority);
  assign _zz_plic_target_bestRequest_valid = (_zz_plic_target_bestRequest_id ? plic_target_requests_0_valid : plic_target_requests_1_valid);
  assign _zz_plic_target_bestRequest_id_1 = ((! plic_target_requests_3_valid) || (plic_target_requests_2_valid && (plic_target_requests_3_priority <= plic_target_requests_2_priority)));
  assign _zz_plic_target_bestRequest_priority_1 = (_zz_plic_target_bestRequest_id_1 ? plic_target_requests_2_priority : plic_target_requests_3_priority);
  assign _zz_plic_target_bestRequest_valid_1 = (_zz_plic_target_bestRequest_id_1 ? plic_target_requests_2_valid : plic_target_requests_3_valid);
  assign _zz_plic_target_bestRequest_priority_2 = ((! _zz_plic_target_bestRequest_valid_1) || (_zz_plic_target_bestRequest_valid && (_zz_plic_target_bestRequest_priority_1 <= _zz_plic_target_bestRequest_priority)));
  assign plic_target_iep = (plic_target_threshold < plic_target_bestRequest_priority);
  assign plic_target_claim = (plic_target_iep ? plic_target_bestRequest_id : 2'b00);
  always @(*) begin
    plic_apb_PREADY = 1'b1;
    if(when_PlicMapper_l122) begin
      plic_apb_PREADY = 1'b0;
    end
  end

  always @(*) begin
    plic_apb_PRDATA = 32'h0;
    case(plic_apb_PADDR)
      26'h0000004 : begin
        plic_apb_PRDATA[0 : 0] = plic_gateways_0_priority;
      end
      26'h0001000 : begin
        plic_apb_PRDATA[1 : 1] = plic_gateways_0_ip;
        plic_apb_PRDATA[2 : 2] = plic_gateways_1_ip;
        plic_apb_PRDATA[3 : 3] = plic_gateways_2_ip;
      end
      26'h0000008 : begin
        plic_apb_PRDATA[0 : 0] = plic_gateways_1_priority;
      end
      26'h000000c : begin
        plic_apb_PRDATA[0 : 0] = plic_gateways_2_priority;
      end
      26'h0200000 : begin
        plic_apb_PRDATA[0 : 0] = plic_target_threshold;
      end
      26'h0200004 : begin
        plic_apb_PRDATA[1 : 0] = plic_target_claim;
      end
      26'h0002000 : begin
        plic_apb_PRDATA[1 : 1] = plic_target_ie_0;
        plic_apb_PRDATA[2 : 2] = plic_target_ie_1;
        plic_apb_PRDATA[3 : 3] = plic_target_ie_2;
      end
      default : begin
      end
    endcase
  end

  assign _zz_1 = ((plic_apb_PSEL[0] && plic_apb_PENABLE) && plic_apb_PWRITE);
  assign _zz_2 = ((plic_apb_PSEL[0] && plic_apb_PENABLE) && (! plic_apb_PWRITE));
  assign _zz_3 = (((plic_apb_PSEL[0] && plic_apb_PENABLE) && plic_apb_PREADY) && plic_apb_PWRITE);
  assign _zz_4 = (((plic_apb_PSEL[0] && plic_apb_PENABLE) && plic_apb_PREADY) && (! plic_apb_PWRITE));
  assign plic_gateways_0_priority = _zz_plic_gateways_0_priority;
  assign plic_gateways_1_priority = _zz_plic_gateways_1_priority;
  assign plic_gateways_2_priority = _zz_plic_gateways_2_priority;
  always @(*) begin
    plic_claim_valid = 1'b0;
    case(plic_apb_PADDR)
      26'h0200004 : begin
        if(_zz_4) begin
          plic_claim_valid = 1'b1;
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    plic_claim_payload = 2'bxx;
    case(plic_apb_PADDR)
      26'h0200004 : begin
        if(_zz_4) begin
          plic_claim_payload = plic_target_claim;
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    plic_completion_valid = 1'b0;
    if(plic_targetMapping_0_targetCompletion_valid) begin
      plic_completion_valid = 1'b1;
    end
  end

  always @(*) begin
    plic_completion_payload = 2'bxx;
    if(plic_targetMapping_0_targetCompletion_valid) begin
      plic_completion_payload = plic_targetMapping_0_targetCompletion_payload;
    end
  end

  always @(*) begin
    plic_coherencyStall_willIncrement = 1'b0;
    if(when_PlicMapper_l122) begin
      plic_coherencyStall_willIncrement = 1'b1;
    end
    if(when_Apb3SlaveFactory_l81) begin
      if(_zz_1) begin
        plic_coherencyStall_willIncrement = 1'b1;
      end
      if(_zz_2) begin
        plic_coherencyStall_willIncrement = 1'b1;
      end
    end
  end

  assign plic_coherencyStall_willClear = 1'b0;
  assign plic_coherencyStall_willOverflowIfInc = (plic_coherencyStall_value == 1'b1);
  assign plic_coherencyStall_willOverflow = (plic_coherencyStall_willOverflowIfInc && plic_coherencyStall_willIncrement);
  always @(*) begin
    plic_coherencyStall_valueNext = (plic_coherencyStall_value + plic_coherencyStall_willIncrement);
    if(plic_coherencyStall_willClear) begin
      plic_coherencyStall_valueNext = 1'b0;
    end
  end

  assign when_PlicMapper_l122 = (plic_coherencyStall_value != 1'b0);
  assign plic_target_threshold = _zz_plic_target_threshold;
  always @(*) begin
    plic_targetMapping_0_targetCompletion_valid = 1'b0;
    case(plic_apb_PADDR)
      26'h0200004 : begin
        if(_zz_3) begin
          plic_targetMapping_0_targetCompletion_valid = 1'b1;
        end
      end
      default : begin
      end
    endcase
  end

  assign plic_target_ie_0 = _zz_plic_target_ie_0;
  assign plic_target_ie_1 = _zz_plic_target_ie_1;
  assign plic_target_ie_2 = _zz_plic_target_ie_2;
  assign plic_targetMapping_0_targetCompletion_payload = plic_apb_PWDATA[1 : 0];
  assign when_Apb3SlaveFactory_l81 = 1'b1;
  assign _zz_FetchL1TileLinkPlugin_logic_down_a_ready = (! _zz_FetchL1TileLinkPlugin_logic_down_a_ready_1);
  assign _zz_5 = _zz_FetchL1TileLinkPlugin_logic_down_a_ready_1;
  assign _zz_io_ups_0_a_payload_opcode_2 = _zz_io_ups_0_a_payload_opcode_3;
  assign _zz_6 = (! _zz_io_ups_0_a_valid_1);
  assign _zz_io_ups_0_a_valid = _zz_io_ups_0_a_valid_1;
  assign _zz_io_ups_0_a_payload_opcode_4 = _zz_io_ups_0_a_payload_opcode_5;
  assign _zz_io_ups_0_a_payload_opcode_1 = _zz_io_ups_0_a_payload_opcode_4;
  always @(*) begin
    _zz_io_ups_0_d_ready = vexiiRiscv_1_FetchL1TileLinkPlugin_logic_down_d_ready;
    if(when_Stream_l393) begin
      _zz_io_ups_0_d_ready = 1'b1;
    end
  end

  assign when_Stream_l393 = (! _zz_when_Stream_l393);
  assign _zz_when_Stream_l393 = _zz_when_Stream_l393_1;
  assign _zz_FetchL1TileLinkPlugin_logic_down_d_payload_opcode_2 = _zz_FetchL1TileLinkPlugin_logic_down_d_payload_opcode_3;
  assign _zz_FetchL1TileLinkPlugin_logic_down_d_payload_opcode = _zz_FetchL1TileLinkPlugin_logic_down_d_payload_opcode_2;
  assign _zz_LsuTileLinkPlugin_logic_bridge_down_a_ready = (! _zz_LsuTileLinkPlugin_logic_bridge_down_a_ready_1);
  assign _zz_io_up_a_valid = _zz_LsuTileLinkPlugin_logic_bridge_down_a_ready_1;
  assign _zz_io_up_a_payload_opcode_2 = _zz_io_up_a_payload_opcode_3;
  assign _zz_io_up_a_payload_opcode_1 = _zz_io_up_a_payload_opcode_2;
  always @(*) begin
    _zz_io_up_d_ready = vexiiRiscv_1_LsuTileLinkPlugin_logic_bridge_down_d_ready;
    if(when_Stream_l393_1) begin
      _zz_io_up_d_ready = 1'b1;
    end
  end

  assign when_Stream_l393_1 = (! _zz_when_Stream_l393_2);
  assign _zz_when_Stream_l393_2 = _zz_when_Stream_l393_3;
  assign _zz_LsuTileLinkPlugin_logic_bridge_down_d_payload_opcode_2 = _zz_LsuTileLinkPlugin_logic_bridge_down_d_payload_opcode_3;
  assign _zz_LsuTileLinkPlugin_logic_bridge_down_d_payload_opcode = _zz_LsuTileLinkPlugin_logic_bridge_down_d_payload_opcode_2;
  assign _zz_LsuL1TileLinkPlugin_logic_down_a_ready = (! _zz_LsuL1TileLinkPlugin_logic_down_a_ready_1);
  assign _zz_io_ups_2_a_valid = _zz_LsuL1TileLinkPlugin_logic_down_a_ready_1;
  assign _zz_io_ups_2_a_payload_opcode_2 = _zz_io_ups_2_a_payload_opcode_3;
  assign _zz_io_ups_2_a_payload_opcode_1 = _zz_io_ups_2_a_payload_opcode_2;
  always @(*) begin
    _zz_io_ups_2_d_ready = vexiiRiscv_1_LsuL1TileLinkPlugin_logic_down_d_ready;
    if(when_Stream_l393_2) begin
      _zz_io_ups_2_d_ready = 1'b1;
    end
  end

  assign when_Stream_l393_2 = (! _zz_when_Stream_l393_4);
  assign _zz_when_Stream_l393_4 = _zz_when_Stream_l393_5;
  assign _zz_LsuL1TileLinkPlugin_logic_down_d_payload_opcode_2 = _zz_LsuL1TileLinkPlugin_logic_down_d_payload_opcode_3;
  assign _zz_LsuL1TileLinkPlugin_logic_down_d_payload_opcode = _zz_LsuL1TileLinkPlugin_logic_down_d_payload_opcode_2;
  assign _zz_io_ups_0_a_payload_opcode = vexiiRiscv_1_FetchL1TileLinkPlugin_logic_down_a_payload_opcode;
  assign _zz_FetchL1TileLinkPlugin_logic_down_d_payload_opcode_4 = arbiter_1_io_ups_0_d_payload_opcode;
  assign _zz_io_down_d_payload_opcode_1 = arbiter_1_io_ups_1_d_payload_opcode;
  assign _zz_LsuL1TileLinkPlugin_logic_down_d_payload_opcode_4 = arbiter_1_io_ups_2_d_payload_opcode;
  assign _zz_io_up_a_payload_opcode_4 = arbiter_1_io_down_a_payload_opcode;
  assign _zz_io_ups_2_a_payload_opcode = vexiiRiscv_1_LsuL1TileLinkPlugin_logic_down_a_payload_opcode;
  assign _zz_io_up_a_payload_opcode_5 = _zz_io_up_a_payload_opcode_6;
  assign _zz_io_down_d_payload_opcode_3 = _zz_io_down_d_payload_opcode_2;
  assign ramBridge_up_bus_a_valid = decoder_2_io_downs_1_a_valid;
  assign ramBridge_up_bus_a_payload_opcode = _zz_ramBridge_up_bus_a_payload_opcode;
  assign ramBridge_up_bus_a_payload_param = decoder_2_io_downs_1_a_payload_param;
  assign ramBridge_up_bus_a_payload_source = decoder_2_io_downs_1_a_payload_source;
  assign ramBridge_up_bus_a_payload_address = decoder_2_io_downs_1_a_payload_address;
  assign ramBridge_up_bus_a_payload_size = decoder_2_io_downs_1_a_payload_size;
  assign ramBridge_up_bus_a_payload_mask = decoder_2_io_downs_1_a_payload_mask;
  assign ramBridge_up_bus_a_payload_data = decoder_2_io_downs_1_a_payload_data;
  assign ramBridge_up_bus_a_payload_corrupt = decoder_2_io_downs_1_a_payload_corrupt;
  assign ramBridge_up_bus_d_ready = decoder_2_io_downs_1_d_ready;
  assign _zz_io_downs_1_d_payload_opcode = ramBridge_up_bus_d_payload_opcode;
  assign _zz_io_ups_0_a_payload_opcode_7 = _zz_io_ups_0_a_payload_opcode_1;
  assign _zz_FetchL1TileLinkPlugin_logic_down_d_payload_opcode_1 = _zz_FetchL1TileLinkPlugin_logic_down_d_payload_opcode_5;
  assign _zz_io_up_a_payload_opcode_7 = _zz_io_up_a_payload_opcode_1;
  assign _zz_LsuTileLinkPlugin_logic_bridge_down_d_payload_opcode_1 = _zz_LsuTileLinkPlugin_logic_bridge_down_d_payload_opcode_4;
  assign _zz_io_ups_2_a_payload_opcode_5 = _zz_io_ups_2_a_payload_opcode_1;
  assign _zz_LsuL1TileLinkPlugin_logic_down_d_payload_opcode_1 = _zz_LsuL1TileLinkPlugin_logic_down_d_payload_opcode_5;
  assign _zz_io_up_a_payload_opcode = vexiiRiscv_1_LsuTileLinkPlugin_logic_bridge_down_a_payload_opcode;
  assign ramBridge_up_bus_a_ready = ramBridge_logic_bridge_io_up_a_ready;
  assign ramBridge_up_bus_d_valid = ramBridge_logic_bridge_io_up_d_valid;
  assign ramBridge_up_bus_d_payload_opcode = ramBridge_logic_bridge_io_up_d_payload_opcode;
  assign ramBridge_up_bus_d_payload_param = ramBridge_logic_bridge_io_up_d_payload_param;
  assign ramBridge_up_bus_d_payload_source = ramBridge_logic_bridge_io_up_d_payload_source;
  assign ramBridge_up_bus_d_payload_size = ramBridge_logic_bridge_io_up_d_payload_size;
  assign ramBridge_up_bus_d_payload_denied = ramBridge_logic_bridge_io_up_d_payload_denied;
  assign ramBridge_up_bus_d_payload_data = ramBridge_logic_bridge_io_up_d_payload_data;
  assign ramBridge_up_bus_d_payload_corrupt = ramBridge_logic_bridge_io_up_d_payload_corrupt;
  assign ramBridge_down_ar_valid = ramBridge_logic_bridge_io_down_ar_valid;
  assign ramBridge_down_ar_payload_addr = ramBridge_logic_bridge_io_down_ar_payload_addr;
  assign ramBridge_down_ar_payload_id = ramBridge_logic_bridge_io_down_ar_payload_id;
  assign ramBridge_down_ar_payload_len = ramBridge_logic_bridge_io_down_ar_payload_len;
  assign ramBridge_down_ar_payload_size = ramBridge_logic_bridge_io_down_ar_payload_size;
  assign ramBridge_down_ar_payload_burst = ramBridge_logic_bridge_io_down_ar_payload_burst;
  assign ramBridge_down_aw_valid = ramBridge_logic_bridge_io_down_aw_valid;
  assign ramBridge_down_aw_payload_addr = ramBridge_logic_bridge_io_down_aw_payload_addr;
  assign ramBridge_down_aw_payload_id = ramBridge_logic_bridge_io_down_aw_payload_id;
  assign ramBridge_down_aw_payload_len = ramBridge_logic_bridge_io_down_aw_payload_len;
  assign ramBridge_down_aw_payload_size = ramBridge_logic_bridge_io_down_aw_payload_size;
  assign ramBridge_down_aw_payload_burst = ramBridge_logic_bridge_io_down_aw_payload_burst;
  assign ramBridge_down_aw_payload_allStrb = ramBridge_logic_bridge_io_down_aw_payload_allStrb;
  assign ramBridge_down_w_valid = ramBridge_logic_bridge_io_down_w_valid;
  assign ramBridge_down_w_payload_data = ramBridge_logic_bridge_io_down_w_payload_data;
  assign ramBridge_down_w_payload_strb = ramBridge_logic_bridge_io_down_w_payload_strb;
  assign ramBridge_down_w_payload_last = ramBridge_logic_bridge_io_down_w_payload_last;
  assign ramBridge_down_r_ready = ramBridge_logic_bridge_io_down_r_ready;
  assign ramBridge_down_b_ready = ramBridge_logic_bridge_io_down_b_ready;
  assign _zz_io_ups_0_a_payload_opcode_6 = _zz_io_ups_0_a_payload_opcode_7;
  assign _zz_FetchL1TileLinkPlugin_logic_down_d_payload_opcode_5 = _zz_FetchL1TileLinkPlugin_logic_down_d_payload_opcode_4;
  assign _zz_LsuTileLinkPlugin_logic_bridge_down_d_payload_opcode_4 = widthAdapter_2_io_up_d_payload_opcode;
  assign _zz_io_ups_1_a_payload_opcode = widthAdapter_2_io_down_a_payload_opcode;
  assign _zz_io_ups_2_a_payload_opcode_4 = _zz_io_ups_2_a_payload_opcode_5;
  assign _zz_LsuL1TileLinkPlugin_logic_down_d_payload_opcode_5 = _zz_LsuL1TileLinkPlugin_logic_down_d_payload_opcode_4;
  assign toApb_up_bus_a_valid = decoder_3_io_downs_0_a_valid;
  assign toApb_up_bus_a_payload_opcode = _zz_toApb_up_bus_a_payload_opcode;
  assign toApb_up_bus_a_payload_param = decoder_3_io_downs_0_a_payload_param;
  assign toApb_up_bus_a_payload_source = decoder_3_io_downs_0_a_payload_source;
  assign toApb_up_bus_a_payload_address = decoder_3_io_downs_0_a_payload_address;
  assign toApb_up_bus_a_payload_size = decoder_3_io_downs_0_a_payload_size;
  assign toApb_up_bus_a_payload_mask = decoder_3_io_downs_0_a_payload_mask;
  assign toApb_up_bus_a_payload_data = decoder_3_io_downs_0_a_payload_data;
  assign toApb_up_bus_a_payload_corrupt = decoder_3_io_downs_0_a_payload_corrupt;
  assign toApb_up_bus_d_ready = decoder_3_io_downs_0_d_ready;
  assign _zz_io_downs_0_d_payload_opcode = toApb_up_bus_d_payload_opcode;
  assign internalRam_up_bus_a_valid = decoder_3_io_downs_1_a_valid;
  assign internalRam_up_bus_a_payload_opcode = _zz_internalRam_up_bus_a_payload_opcode;
  assign internalRam_up_bus_a_payload_param = decoder_3_io_downs_1_a_payload_param;
  assign internalRam_up_bus_a_payload_source = decoder_3_io_downs_1_a_payload_source;
  assign internalRam_up_bus_a_payload_address = decoder_3_io_downs_1_a_payload_address;
  assign internalRam_up_bus_a_payload_size = decoder_3_io_downs_1_a_payload_size;
  assign internalRam_up_bus_a_payload_mask = decoder_3_io_downs_1_a_payload_mask;
  assign internalRam_up_bus_a_payload_data = decoder_3_io_downs_1_a_payload_data;
  assign internalRam_up_bus_a_payload_corrupt = decoder_3_io_downs_1_a_payload_corrupt;
  assign internalRam_up_bus_d_ready = decoder_3_io_downs_1_d_ready;
  assign _zz_io_downs_1_d_payload_opcode_1 = internalRam_up_bus_d_payload_opcode;
  assign ramBridge_down_ar_ready = streamArbiter_10_io_inputs_0_ready;
  assign ramBridge_down_aw_ready = streamArbiter_10_io_inputs_1_ready;
  assign ram_axi_arw_valid = streamArbiter_10_io_output_valid;
  assign ram_axi_arw_payload_addr = streamArbiter_10_io_output_payload_addr;
  assign ram_axi_arw_payload_id = streamArbiter_10_io_output_payload_id;
  assign ram_axi_arw_payload_len = streamArbiter_10_io_output_payload_len;
  assign ram_axi_arw_payload_size = streamArbiter_10_io_output_payload_size;
  assign ram_axi_arw_payload_burst = streamArbiter_10_io_output_payload_burst;
  assign ram_axi_arw_payload_allStrb = streamArbiter_10_io_output_payload_allStrb;
  assign ram_axi_arw_payload_write = streamArbiter_10_io_chosenOH[1];
  assign ram_axi_w_valid = ramBridge_down_w_valid;
  assign ramBridge_down_w_ready = ram_axi_w_ready;
  assign ram_axi_w_payload_data = ramBridge_down_w_payload_data;
  assign ram_axi_w_payload_strb = ramBridge_down_w_payload_strb;
  assign ram_axi_w_payload_last = ramBridge_down_w_payload_last;
  assign ramBridge_down_b_valid = ram_axi_b_valid;
  assign ram_axi_b_ready = ramBridge_down_b_ready;
  assign ramBridge_down_b_payload_id = ram_axi_b_payload_id;
  assign ramBridge_down_b_payload_resp = ram_axi_b_payload_resp;
  assign ramBridge_down_r_valid = ram_axi_r_valid;
  assign ram_axi_r_ready = ramBridge_down_r_ready;
  assign ramBridge_down_r_payload_data = ram_axi_r_payload_data;
  assign ramBridge_down_r_payload_id = ram_axi_r_payload_id;
  assign ramBridge_down_r_payload_resp = ram_axi_r_payload_resp;
  assign ramBridge_down_r_payload_last = ram_axi_r_payload_last;
  assign io_ddr_sdram_ck_p = ram_ddr_ctrl_ddr_ck_p;
  assign io_ddr_sdram_ck_n = ram_ddr_ctrl_ddr_ck_n;
  assign io_ddr_sdram_cke = ram_ddr_ctrl_ddr_cke;
  assign io_ddr_sdram_ras_n = ram_ddr_ctrl_ddr_ras_n;
  assign io_ddr_sdram_cas_n = ram_ddr_ctrl_ddr_cas_n;
  assign io_ddr_sdram_we_n = ram_ddr_ctrl_ddr_we_n;
  assign io_ddr_sdram_ba = ram_ddr_ctrl_ddr_ba;
  assign io_ddr_sdram_a = ram_ddr_ctrl_ddr_a;
  assign io_ddr_sdram_dm = ram_ddr_ctrl_ddr_dm;
  assign ram_axi_arw_ready = ram_axi_cc_io_input_arw_ready;
  assign ram_axi_w_ready = ram_axi_cc_io_input_w_ready;
  assign ram_axi_b_valid = ram_axi_cc_io_input_b_valid;
  assign ram_axi_b_payload_id = ram_axi_cc_io_input_b_payload_id;
  assign ram_axi_b_payload_resp = ram_axi_cc_io_input_b_payload_resp;
  assign ram_axi_r_valid = ram_axi_cc_io_input_r_valid;
  assign ram_axi_r_payload_data = ram_axi_cc_io_input_r_payload_data;
  assign ram_axi_r_payload_id = ram_axi_cc_io_input_r_payload_id;
  assign ram_axi_r_payload_resp = ram_axi_cc_io_input_r_payload_resp;
  assign ram_axi_r_payload_last = ram_axi_cc_io_input_r_payload_last;
  assign vexiiRiscv_1_PrivilegedPlugin_logic_harts_0_int_m_timer = (|1'b0);
  assign vexiiRiscv_1_PrivilegedPlugin_logic_harts_0_int_m_software = (|1'b0);
  assign vexiiRiscv_1_PrivilegedPlugin_logic_harts_0_int_m_external = (|1'b0);
  assign vexiiRiscv_1_PrivilegedPlugin_logic_harts_0_int_s_external = (|1'b0);
  assign _zz_io_up_a_payload_opcode_8 = decoder_2_io_downs_0_a_payload_opcode;
  assign _zz_ramBridge_up_bus_a_payload_opcode_1 = decoder_2_io_downs_1_a_payload_opcode;
  assign _zz_io_down_d_payload_opcode = decoder_2_io_up_d_payload_opcode;
  assign toApb_up_bus_a_ready = toApb_logic_bridge_io_up_a_ready;
  assign toApb_up_bus_d_valid = toApb_logic_bridge_io_up_d_valid;
  assign toApb_up_bus_d_payload_opcode = toApb_logic_bridge_io_up_d_payload_opcode;
  assign toApb_up_bus_d_payload_param = toApb_logic_bridge_io_up_d_payload_param;
  assign toApb_up_bus_d_payload_source = toApb_logic_bridge_io_up_d_payload_source;
  assign toApb_up_bus_d_payload_size = toApb_logic_bridge_io_up_d_payload_size;
  assign toApb_up_bus_d_payload_denied = toApb_logic_bridge_io_up_d_payload_denied;
  assign toApb_up_bus_d_payload_data = toApb_logic_bridge_io_up_d_payload_data;
  assign toApb_up_bus_d_payload_corrupt = toApb_logic_bridge_io_up_d_payload_corrupt;
  assign toApb_down_PADDR = toApb_logic_bridge_io_down_PADDR;
  assign toApb_down_PSEL = toApb_logic_bridge_io_down_PSEL;
  assign toApb_down_PENABLE = toApb_logic_bridge_io_down_PENABLE;
  assign toApb_down_PWRITE = toApb_logic_bridge_io_down_PWRITE;
  assign toApb_down_PWDATA = toApb_logic_bridge_io_down_PWDATA;
  assign internalRam_up_bus_a_ready = internalRam_thread_logic_io_up_a_ready;
  assign internalRam_up_bus_d_valid = internalRam_thread_logic_io_up_d_valid;
  assign internalRam_up_bus_d_payload_opcode = internalRam_thread_logic_io_up_d_payload_opcode;
  assign internalRam_up_bus_d_payload_param = internalRam_thread_logic_io_up_d_payload_param;
  assign internalRam_up_bus_d_payload_source = internalRam_thread_logic_io_up_d_payload_source;
  assign internalRam_up_bus_d_payload_size = internalRam_thread_logic_io_up_d_payload_size;
  assign internalRam_up_bus_d_payload_denied = internalRam_thread_logic_io_up_d_payload_denied;
  assign internalRam_up_bus_d_payload_data = internalRam_thread_logic_io_up_d_payload_data;
  assign internalRam_up_bus_d_payload_corrupt = internalRam_thread_logic_io_up_d_payload_corrupt;
  assign _zz_io_downs_0_d_payload_opcode_1 = widthAdapter_3_io_up_d_payload_opcode;
  assign _zz_io_up_a_payload_opcode_6 = widthAdapter_3_io_down_a_payload_opcode;
  assign _zz_ramBridge_up_bus_a_payload_opcode = _zz_ramBridge_up_bus_a_payload_opcode_1;
  assign _zz_io_downs_1_d_payload_opcode_2 = _zz_io_downs_1_d_payload_opcode;
  assign _zz_toApb_up_bus_a_payload_opcode_1 = decoder_3_io_downs_0_a_payload_opcode;
  assign _zz_internalRam_up_bus_a_payload_opcode_1 = decoder_3_io_downs_1_a_payload_opcode;
  assign _zz_io_down_d_payload_opcode_2 = decoder_3_io_up_d_payload_opcode;
  assign toApb_down_PREADY = toApb_down_decoder_io_input_PREADY;
  assign toApb_down_PRDATA = toApb_down_decoder_io_input_PRDATA;
  assign toApb_down_PSLVERROR = toApb_down_decoder_io_input_PSLVERROR;
  assign peripheral_apb_bridge_input_PADDR = apb3Router_3_io_outputs_0_PADDR[18:0];
  assign board_ctrl_apb_PADDR = apb3Router_3_io_outputs_1_PADDR[4:0];
  assign video_ctrl_apb_PADDR = apb3Router_3_io_outputs_2_PADDR[4:0];
  assign plic_apb_PADDR = apb3Router_3_io_outputs_3_PADDR[25:0];
  assign plic_apb_PSEL = apb3Router_3_io_outputs_3_PSEL;
  assign plic_apb_PENABLE = apb3Router_3_io_outputs_3_PENABLE;
  assign plic_apb_PWRITE = apb3Router_3_io_outputs_3_PWRITE;
  assign plic_apb_PWDATA = apb3Router_3_io_outputs_3_PWDATA;
  assign _zz_toApb_up_bus_a_payload_opcode = _zz_toApb_up_bus_a_payload_opcode_1;
  assign _zz_io_downs_0_d_payload_opcode_2 = _zz_io_downs_0_d_payload_opcode;
  assign _zz_internalRam_up_bus_a_payload_opcode = _zz_internalRam_up_bus_a_payload_opcode_1;
  assign _zz_io_downs_1_d_payload_opcode_3 = _zz_io_downs_1_d_payload_opcode_1;
  always @(posedge board_ctrl_clk_cpu) begin
    usb_interrupt <= peripheral_usb_ctrl_io_interrupt;
    plic_target_bestRequest_priority <= (_zz_plic_target_bestRequest_priority_2 ? _zz_plic_target_bestRequest_priority : _zz_plic_target_bestRequest_priority_1);
    plic_target_bestRequest_id <= (_zz_plic_target_bestRequest_priority_2 ? (_zz_plic_target_bestRequest_id ? plic_target_requests_0_id : plic_target_requests_1_id) : (_zz_plic_target_bestRequest_id_1 ? plic_target_requests_2_id : plic_target_requests_3_id));
    plic_target_bestRequest_valid <= (_zz_plic_target_bestRequest_priority_2 ? _zz_plic_target_bestRequest_valid : _zz_plic_target_bestRequest_valid_1);
    if(_zz_FetchL1TileLinkPlugin_logic_down_a_ready) begin
      _zz_io_ups_0_a_payload_opcode_3 <= _zz_io_ups_0_a_payload_opcode;
      _zz_io_ups_0_a_payload_param <= vexiiRiscv_1_FetchL1TileLinkPlugin_logic_down_a_payload_param;
      _zz_io_ups_0_a_payload_address <= vexiiRiscv_1_FetchL1TileLinkPlugin_logic_down_a_payload_address;
      _zz_io_ups_0_a_payload_size <= vexiiRiscv_1_FetchL1TileLinkPlugin_logic_down_a_payload_size;
    end
    if(_zz_6) begin
      _zz_io_ups_0_a_payload_opcode_5 <= _zz_io_ups_0_a_payload_opcode_2;
      _zz_io_ups_0_a_payload_param_1 <= _zz_io_ups_0_a_payload_param;
      _zz_io_ups_0_a_payload_address_1 <= _zz_io_ups_0_a_payload_address;
      _zz_io_ups_0_a_payload_size_1 <= _zz_io_ups_0_a_payload_size;
    end
    if(_zz_io_ups_0_d_ready) begin
      _zz_FetchL1TileLinkPlugin_logic_down_d_payload_opcode_3 <= _zz_FetchL1TileLinkPlugin_logic_down_d_payload_opcode_1;
      _zz_FetchL1TileLinkPlugin_logic_down_d_payload_param <= arbiter_1_io_ups_0_d_payload_param;
      _zz_FetchL1TileLinkPlugin_logic_down_d_payload_size <= arbiter_1_io_ups_0_d_payload_size;
      _zz_FetchL1TileLinkPlugin_logic_down_d_payload_denied <= arbiter_1_io_ups_0_d_payload_denied;
      _zz_FetchL1TileLinkPlugin_logic_down_d_payload_data <= arbiter_1_io_ups_0_d_payload_data;
      _zz_FetchL1TileLinkPlugin_logic_down_d_payload_corrupt <= arbiter_1_io_ups_0_d_payload_corrupt;
    end
    if(_zz_LsuTileLinkPlugin_logic_bridge_down_a_ready) begin
      _zz_io_up_a_payload_opcode_3 <= _zz_io_up_a_payload_opcode;
      _zz_io_up_a_payload_param <= vexiiRiscv_1_LsuTileLinkPlugin_logic_bridge_down_a_payload_param;
      _zz_io_up_a_payload_address <= vexiiRiscv_1_LsuTileLinkPlugin_logic_bridge_down_a_payload_address;
      _zz_io_up_a_payload_size <= vexiiRiscv_1_LsuTileLinkPlugin_logic_bridge_down_a_payload_size;
      _zz_io_up_a_payload_mask <= vexiiRiscv_1_LsuTileLinkPlugin_logic_bridge_down_a_payload_mask;
      _zz_io_up_a_payload_data <= vexiiRiscv_1_LsuTileLinkPlugin_logic_bridge_down_a_payload_data;
      _zz_io_up_a_payload_corrupt <= vexiiRiscv_1_LsuTileLinkPlugin_logic_bridge_down_a_payload_corrupt;
    end
    if(_zz_io_up_d_ready) begin
      _zz_LsuTileLinkPlugin_logic_bridge_down_d_payload_opcode_3 <= _zz_LsuTileLinkPlugin_logic_bridge_down_d_payload_opcode_1;
      _zz_LsuTileLinkPlugin_logic_bridge_down_d_payload_param <= widthAdapter_2_io_up_d_payload_param;
      _zz_LsuTileLinkPlugin_logic_bridge_down_d_payload_size <= widthAdapter_2_io_up_d_payload_size;
      _zz_LsuTileLinkPlugin_logic_bridge_down_d_payload_denied <= widthAdapter_2_io_up_d_payload_denied;
      _zz_LsuTileLinkPlugin_logic_bridge_down_d_payload_data <= widthAdapter_2_io_up_d_payload_data;
      _zz_LsuTileLinkPlugin_logic_bridge_down_d_payload_corrupt <= widthAdapter_2_io_up_d_payload_corrupt;
    end
    if(_zz_LsuL1TileLinkPlugin_logic_down_a_ready) begin
      _zz_io_ups_2_a_payload_opcode_3 <= _zz_io_ups_2_a_payload_opcode;
      _zz_io_ups_2_a_payload_param <= vexiiRiscv_1_LsuL1TileLinkPlugin_logic_down_a_payload_param;
      _zz_io_ups_2_a_payload_source <= vexiiRiscv_1_LsuL1TileLinkPlugin_logic_down_a_payload_source;
      _zz_io_ups_2_a_payload_address <= vexiiRiscv_1_LsuL1TileLinkPlugin_logic_down_a_payload_address;
      _zz_io_ups_2_a_payload_size <= vexiiRiscv_1_LsuL1TileLinkPlugin_logic_down_a_payload_size;
      _zz_io_ups_2_a_payload_mask <= vexiiRiscv_1_LsuL1TileLinkPlugin_logic_down_a_payload_mask;
      _zz_io_ups_2_a_payload_data <= vexiiRiscv_1_LsuL1TileLinkPlugin_logic_down_a_payload_data;
      _zz_io_ups_2_a_payload_corrupt <= vexiiRiscv_1_LsuL1TileLinkPlugin_logic_down_a_payload_corrupt;
    end
    if(_zz_io_ups_2_d_ready) begin
      _zz_LsuL1TileLinkPlugin_logic_down_d_payload_opcode_3 <= _zz_LsuL1TileLinkPlugin_logic_down_d_payload_opcode_1;
      _zz_LsuL1TileLinkPlugin_logic_down_d_payload_param <= arbiter_1_io_ups_2_d_payload_param;
      _zz_LsuL1TileLinkPlugin_logic_down_d_payload_source <= arbiter_1_io_ups_2_d_payload_source;
      _zz_LsuL1TileLinkPlugin_logic_down_d_payload_size <= arbiter_1_io_ups_2_d_payload_size;
      _zz_LsuL1TileLinkPlugin_logic_down_d_payload_denied <= arbiter_1_io_ups_2_d_payload_denied;
      _zz_LsuL1TileLinkPlugin_logic_down_d_payload_data <= arbiter_1_io_ups_2_d_payload_data;
      _zz_LsuL1TileLinkPlugin_logic_down_d_payload_corrupt <= arbiter_1_io_ups_2_d_payload_corrupt;
    end
  end

  always @(posedge board_ctrl_clk_cpu or posedge board_ctrl_reset_cpu) begin
    if(board_ctrl_reset_cpu) begin
      plic_gateways_0_ip <= 1'b0;
      plic_gateways_0_waitCompletion <= 1'b0;
      plic_gateways_1_ip <= 1'b0;
      plic_gateways_1_waitCompletion <= 1'b0;
      plic_gateways_2_ip <= 1'b0;
      plic_gateways_2_waitCompletion <= 1'b0;
      _zz_plic_gateways_0_priority <= 1'b0;
      _zz_plic_gateways_1_priority <= 1'b0;
      _zz_plic_gateways_2_priority <= 1'b0;
      plic_coherencyStall_value <= 1'b0;
      _zz_plic_target_threshold <= 1'b0;
      _zz_plic_target_ie_0 <= 1'b0;
      _zz_plic_target_ie_1 <= 1'b0;
      _zz_plic_target_ie_2 <= 1'b0;
      _zz_FetchL1TileLinkPlugin_logic_down_a_ready_1 <= 1'b0;
      _zz_io_ups_0_a_valid_1 <= 1'b0;
      _zz_when_Stream_l393_1 <= 1'b0;
      _zz_LsuTileLinkPlugin_logic_bridge_down_a_ready_1 <= 1'b0;
      _zz_when_Stream_l393_3 <= 1'b0;
      _zz_LsuL1TileLinkPlugin_logic_down_a_ready_1 <= 1'b0;
      _zz_when_Stream_l393_5 <= 1'b0;
    end else begin
      if(when_PlicGateway_l21) begin
        plic_gateways_0_ip <= peripheral_uart_ctrl_interrupt;
        plic_gateways_0_waitCompletion <= peripheral_uart_ctrl_interrupt;
      end
      if(when_PlicGateway_l21_1) begin
        plic_gateways_1_ip <= peripheral_sdcard_ctrl_interrupt;
        plic_gateways_1_waitCompletion <= peripheral_sdcard_ctrl_interrupt;
      end
      if(when_PlicGateway_l21_2) begin
        plic_gateways_2_ip <= usb_interrupt;
        plic_gateways_2_waitCompletion <= usb_interrupt;
      end
      if(plic_claim_valid) begin
        case(plic_claim_payload)
          2'b01 : begin
            plic_gateways_0_ip <= 1'b0;
          end
          2'b10 : begin
            plic_gateways_1_ip <= 1'b0;
          end
          2'b11 : begin
            plic_gateways_2_ip <= 1'b0;
          end
          default : begin
          end
        endcase
      end
      if(plic_completion_valid) begin
        case(plic_completion_payload)
          2'b01 : begin
            plic_gateways_0_waitCompletion <= 1'b0;
          end
          2'b10 : begin
            plic_gateways_1_waitCompletion <= 1'b0;
          end
          2'b11 : begin
            plic_gateways_2_waitCompletion <= 1'b0;
          end
          default : begin
          end
        endcase
      end
      plic_coherencyStall_value <= plic_coherencyStall_valueNext;
      case(plic_apb_PADDR)
        26'h0000004 : begin
          if(_zz_3) begin
            _zz_plic_gateways_0_priority <= plic_apb_PWDATA[0 : 0];
          end
        end
        26'h0000008 : begin
          if(_zz_3) begin
            _zz_plic_gateways_1_priority <= plic_apb_PWDATA[0 : 0];
          end
        end
        26'h000000c : begin
          if(_zz_3) begin
            _zz_plic_gateways_2_priority <= plic_apb_PWDATA[0 : 0];
          end
        end
        26'h0200000 : begin
          if(_zz_3) begin
            _zz_plic_target_threshold <= plic_apb_PWDATA[0 : 0];
          end
        end
        26'h0002000 : begin
          if(_zz_3) begin
            _zz_plic_target_ie_0 <= plic_apb_PWDATA[1];
            _zz_plic_target_ie_1 <= plic_apb_PWDATA[2];
            _zz_plic_target_ie_2 <= plic_apb_PWDATA[3];
          end
        end
        default : begin
        end
      endcase
      if(vexiiRiscv_1_FetchL1TileLinkPlugin_logic_down_a_valid) begin
        _zz_FetchL1TileLinkPlugin_logic_down_a_ready_1 <= 1'b1;
      end
      if((_zz_5 && _zz_6)) begin
        _zz_FetchL1TileLinkPlugin_logic_down_a_ready_1 <= 1'b0;
      end
      if(_zz_5) begin
        _zz_io_ups_0_a_valid_1 <= 1'b1;
      end
      if((_zz_io_ups_0_a_valid && arbiter_1_io_ups_0_a_ready)) begin
        _zz_io_ups_0_a_valid_1 <= 1'b0;
      end
      if(_zz_io_ups_0_d_ready) begin
        _zz_when_Stream_l393_1 <= arbiter_1_io_ups_0_d_valid;
      end
      if(vexiiRiscv_1_LsuTileLinkPlugin_logic_bridge_down_a_valid) begin
        _zz_LsuTileLinkPlugin_logic_bridge_down_a_ready_1 <= 1'b1;
      end
      if((_zz_io_up_a_valid && widthAdapter_2_io_up_a_ready)) begin
        _zz_LsuTileLinkPlugin_logic_bridge_down_a_ready_1 <= 1'b0;
      end
      if(_zz_io_up_d_ready) begin
        _zz_when_Stream_l393_3 <= widthAdapter_2_io_up_d_valid;
      end
      if(vexiiRiscv_1_LsuL1TileLinkPlugin_logic_down_a_valid) begin
        _zz_LsuL1TileLinkPlugin_logic_down_a_ready_1 <= 1'b1;
      end
      if((_zz_io_ups_2_a_valid && arbiter_1_io_ups_2_a_ready)) begin
        _zz_LsuL1TileLinkPlugin_logic_down_a_ready_1 <= 1'b0;
      end
      if(_zz_io_ups_2_d_ready) begin
        _zz_when_Stream_l393_5 <= arbiter_1_io_ups_2_d_valid;
      end
    end
  end


endmodule

module Apb3Router_1 (
  input  wire [26:0]   io_input_PADDR,
  input  wire [3:0]    io_input_PSEL,
  input  wire          io_input_PENABLE,
  output wire          io_input_PREADY,
  input  wire          io_input_PWRITE,
  input  wire [31:0]   io_input_PWDATA,
  output wire [31:0]   io_input_PRDATA,
  output wire          io_input_PSLVERROR,
  output wire [26:0]   io_outputs_0_PADDR,
  output wire [0:0]    io_outputs_0_PSEL,
  output wire          io_outputs_0_PENABLE,
  input  wire          io_outputs_0_PREADY,
  output wire          io_outputs_0_PWRITE,
  output wire [31:0]   io_outputs_0_PWDATA,
  input  wire [31:0]   io_outputs_0_PRDATA,
  input  wire          io_outputs_0_PSLVERROR,
  output wire [26:0]   io_outputs_1_PADDR,
  output wire [0:0]    io_outputs_1_PSEL,
  output wire          io_outputs_1_PENABLE,
  input  wire          io_outputs_1_PREADY,
  output wire          io_outputs_1_PWRITE,
  output wire [31:0]   io_outputs_1_PWDATA,
  input  wire [31:0]   io_outputs_1_PRDATA,
  input  wire          io_outputs_1_PSLVERROR,
  output wire [26:0]   io_outputs_2_PADDR,
  output wire [0:0]    io_outputs_2_PSEL,
  output wire          io_outputs_2_PENABLE,
  input  wire          io_outputs_2_PREADY,
  output wire          io_outputs_2_PWRITE,
  output wire [31:0]   io_outputs_2_PWDATA,
  input  wire [31:0]   io_outputs_2_PRDATA,
  input  wire          io_outputs_2_PSLVERROR,
  output wire [26:0]   io_outputs_3_PADDR,
  output wire [0:0]    io_outputs_3_PSEL,
  output wire          io_outputs_3_PENABLE,
  input  wire          io_outputs_3_PREADY,
  output wire          io_outputs_3_PWRITE,
  output wire [31:0]   io_outputs_3_PWDATA,
  input  wire [31:0]   io_outputs_3_PRDATA,
  input  wire          io_outputs_3_PSLVERROR,
  input  wire          clk_cpu,
  input  wire          reset_cpu
);

  reg                 _zz_io_input_PREADY;
  reg        [31:0]   _zz_io_input_PRDATA;
  reg                 _zz_io_input_PSLVERROR;
  wire                _zz_selIndex;
  wire                _zz_selIndex_1;
  wire                _zz_selIndex_2;
  reg        [1:0]    selIndex;

  always @(*) begin
    case(selIndex)
      2'b00 : begin
        _zz_io_input_PREADY = io_outputs_0_PREADY;
        _zz_io_input_PRDATA = io_outputs_0_PRDATA;
        _zz_io_input_PSLVERROR = io_outputs_0_PSLVERROR;
      end
      2'b01 : begin
        _zz_io_input_PREADY = io_outputs_1_PREADY;
        _zz_io_input_PRDATA = io_outputs_1_PRDATA;
        _zz_io_input_PSLVERROR = io_outputs_1_PSLVERROR;
      end
      2'b10 : begin
        _zz_io_input_PREADY = io_outputs_2_PREADY;
        _zz_io_input_PRDATA = io_outputs_2_PRDATA;
        _zz_io_input_PSLVERROR = io_outputs_2_PSLVERROR;
      end
      default : begin
        _zz_io_input_PREADY = io_outputs_3_PREADY;
        _zz_io_input_PRDATA = io_outputs_3_PRDATA;
        _zz_io_input_PSLVERROR = io_outputs_3_PSLVERROR;
      end
    endcase
  end

  assign io_outputs_0_PADDR = io_input_PADDR;
  assign io_outputs_0_PENABLE = io_input_PENABLE;
  assign io_outputs_0_PSEL[0] = io_input_PSEL[0];
  assign io_outputs_0_PWRITE = io_input_PWRITE;
  assign io_outputs_0_PWDATA = io_input_PWDATA;
  assign io_outputs_1_PADDR = io_input_PADDR;
  assign io_outputs_1_PENABLE = io_input_PENABLE;
  assign io_outputs_1_PSEL[0] = io_input_PSEL[1];
  assign io_outputs_1_PWRITE = io_input_PWRITE;
  assign io_outputs_1_PWDATA = io_input_PWDATA;
  assign io_outputs_2_PADDR = io_input_PADDR;
  assign io_outputs_2_PENABLE = io_input_PENABLE;
  assign io_outputs_2_PSEL[0] = io_input_PSEL[2];
  assign io_outputs_2_PWRITE = io_input_PWRITE;
  assign io_outputs_2_PWDATA = io_input_PWDATA;
  assign io_outputs_3_PADDR = io_input_PADDR;
  assign io_outputs_3_PENABLE = io_input_PENABLE;
  assign io_outputs_3_PSEL[0] = io_input_PSEL[3];
  assign io_outputs_3_PWRITE = io_input_PWRITE;
  assign io_outputs_3_PWDATA = io_input_PWDATA;
  assign _zz_selIndex = io_input_PSEL[3];
  assign _zz_selIndex_1 = (io_input_PSEL[1] || _zz_selIndex);
  assign _zz_selIndex_2 = (io_input_PSEL[2] || _zz_selIndex);
  assign io_input_PREADY = _zz_io_input_PREADY;
  assign io_input_PRDATA = _zz_io_input_PRDATA;
  assign io_input_PSLVERROR = _zz_io_input_PSLVERROR;
  always @(posedge clk_cpu) begin
    selIndex <= {_zz_selIndex_2,_zz_selIndex_1};
  end


endmodule

module Apb3Decoder_1 (
  input  wire [26:0]   io_input_PADDR,
  input  wire [0:0]    io_input_PSEL,
  input  wire          io_input_PENABLE,
  output reg           io_input_PREADY,
  input  wire          io_input_PWRITE,
  input  wire [31:0]   io_input_PWDATA,
  output wire [31:0]   io_input_PRDATA,
  output reg           io_input_PSLVERROR,
  output wire [26:0]   io_output_PADDR,
  output reg  [3:0]    io_output_PSEL,
  output wire          io_output_PENABLE,
  input  wire          io_output_PREADY,
  output wire          io_output_PWRITE,
  output wire [31:0]   io_output_PWDATA,
  input  wire [31:0]   io_output_PRDATA,
  input  wire          io_output_PSLVERROR
);

  wire                when_Apb3Decoder_l88;

  assign io_output_PADDR = io_input_PADDR;
  assign io_output_PENABLE = io_input_PENABLE;
  assign io_output_PWRITE = io_input_PWRITE;
  assign io_output_PWDATA = io_input_PWDATA;
  always @(*) begin
    io_output_PSEL[0] = (((io_input_PADDR & (~ 27'h007ffff)) == 27'h0) && io_input_PSEL[0]);
    io_output_PSEL[1] = (((io_input_PADDR & (~ 27'h000001f)) == 27'h0080000) && io_input_PSEL[0]);
    io_output_PSEL[2] = (((io_input_PADDR & (~ 27'h000001f)) == 27'h0090000) && io_input_PSEL[0]);
    io_output_PSEL[3] = (((io_input_PADDR & (~ 27'h3ffffff)) == 27'h4000000) && io_input_PSEL[0]);
  end

  always @(*) begin
    io_input_PREADY = io_output_PREADY;
    if(when_Apb3Decoder_l88) begin
      io_input_PREADY = 1'b1;
    end
  end

  assign io_input_PRDATA = io_output_PRDATA;
  always @(*) begin
    io_input_PSLVERROR = io_output_PSLVERROR;
    if(when_Apb3Decoder_l88) begin
      io_input_PSLVERROR = 1'b1;
    end
  end

  assign when_Apb3Decoder_l88 = (io_input_PSEL[0] && (io_output_PSEL == 4'b0000));

endmodule

module Decoder_1 (
  input  wire          io_up_a_valid,
  output wire          io_up_a_ready,
  input  wire [2:0]    io_up_a_payload_opcode,
  input  wire [2:0]    io_up_a_payload_param,
  input  wire [2:0]    io_up_a_payload_source,
  input  wire [30:0]   io_up_a_payload_address,
  input  wire [2:0]    io_up_a_payload_size,
  input  wire [3:0]    io_up_a_payload_mask,
  input  wire [31:0]   io_up_a_payload_data,
  input  wire          io_up_a_payload_corrupt,
  output wire          io_up_d_valid,
  input  wire          io_up_d_ready,
  output wire [2:0]    io_up_d_payload_opcode,
  output wire [2:0]    io_up_d_payload_param,
  output wire [2:0]    io_up_d_payload_source,
  output wire [2:0]    io_up_d_payload_size,
  output wire          io_up_d_payload_denied,
  output wire [31:0]   io_up_d_payload_data,
  output wire          io_up_d_payload_corrupt,
  output wire          io_downs_0_a_valid,
  input  wire          io_downs_0_a_ready,
  output wire [2:0]    io_downs_0_a_payload_opcode,
  output wire [2:0]    io_downs_0_a_payload_param,
  output wire [2:0]    io_downs_0_a_payload_source,
  output wire [26:0]   io_downs_0_a_payload_address,
  output wire [2:0]    io_downs_0_a_payload_size,
  output wire [3:0]    io_downs_0_a_payload_mask,
  output wire [31:0]   io_downs_0_a_payload_data,
  output wire          io_downs_0_a_payload_corrupt,
  input  wire          io_downs_0_d_valid,
  output wire          io_downs_0_d_ready,
  input  wire [2:0]    io_downs_0_d_payload_opcode,
  input  wire [2:0]    io_downs_0_d_payload_param,
  input  wire [2:0]    io_downs_0_d_payload_source,
  input  wire [2:0]    io_downs_0_d_payload_size,
  input  wire          io_downs_0_d_payload_denied,
  input  wire [31:0]   io_downs_0_d_payload_data,
  input  wire          io_downs_0_d_payload_corrupt,
  output wire          io_downs_1_a_valid,
  input  wire          io_downs_1_a_ready,
  output wire [2:0]    io_downs_1_a_payload_opcode,
  output wire [2:0]    io_downs_1_a_payload_param,
  output wire [2:0]    io_downs_1_a_payload_source,
  output wire [13:0]   io_downs_1_a_payload_address,
  output wire [2:0]    io_downs_1_a_payload_size,
  output wire [3:0]    io_downs_1_a_payload_mask,
  output wire [31:0]   io_downs_1_a_payload_data,
  output wire          io_downs_1_a_payload_corrupt,
  input  wire          io_downs_1_d_valid,
  output wire          io_downs_1_d_ready,
  input  wire [2:0]    io_downs_1_d_payload_opcode,
  input  wire [2:0]    io_downs_1_d_payload_param,
  input  wire [2:0]    io_downs_1_d_payload_source,
  input  wire [2:0]    io_downs_1_d_payload_size,
  input  wire          io_downs_1_d_payload_denied,
  input  wire [31:0]   io_downs_1_d_payload_data,
  input  wire          io_downs_1_d_payload_corrupt,
  input  wire          clk_cpu,
  input  wire          reset_cpu
);
  localparam A_PUT_FULL_DATA = 3'd0;
  localparam A_PUT_PARTIAL_DATA = 3'd1;
  localparam A_GET = 3'd4;
  localparam A_ACQUIRE_BLOCK = 3'd6;
  localparam A_ACQUIRE_PERM = 3'd7;
  localparam D_ACCESS_ACK = 3'd0;
  localparam D_ACCESS_ACK_DATA = 3'd1;
  localparam D_GRANT = 3'd4;
  localparam D_GRANT_DATA = 3'd5;
  localparam D_RELEASE_ACK = 3'd6;

  wire                d_arbiter_io_inputs_0_ready;
  wire                d_arbiter_io_inputs_1_ready;
  wire                d_arbiter_io_output_valid;
  wire       [2:0]    d_arbiter_io_output_payload_opcode;
  wire       [2:0]    d_arbiter_io_output_payload_param;
  wire       [2:0]    d_arbiter_io_output_payload_source;
  wire       [2:0]    d_arbiter_io_output_payload_size;
  wire                d_arbiter_io_output_payload_denied;
  wire       [31:0]   d_arbiter_io_output_payload_data;
  wire                d_arbiter_io_output_payload_corrupt;
  wire       [0:0]    d_arbiter_io_chosen;
  wire       [1:0]    d_arbiter_io_chosenOH;
  wire       [0:0]    _zz_a_logic_0_hit;
  wire       [30:0]   _zz_downs_0_a_payload_address;
  wire       [0:0]    _zz_a_logic_1_hit;
  wire       [30:0]   _zz_downs_1_a_payload_address;
  reg        [1:0]    _zz_1;
  wire       [1:0]    _zz_2;
  wire                downs_0_a_valid;
  wire                downs_0_a_ready;
  wire       [2:0]    downs_0_a_payload_opcode;
  wire       [2:0]    downs_0_a_payload_param;
  wire       [2:0]    downs_0_a_payload_source;
  wire       [26:0]   downs_0_a_payload_address;
  wire       [2:0]    downs_0_a_payload_size;
  wire       [3:0]    downs_0_a_payload_mask;
  wire       [31:0]   downs_0_a_payload_data;
  wire                downs_0_a_payload_corrupt;
  wire                downs_0_d_valid;
  wire                downs_0_d_ready;
  wire       [2:0]    downs_0_d_payload_opcode;
  wire       [2:0]    downs_0_d_payload_param;
  wire       [2:0]    downs_0_d_payload_source;
  wire       [2:0]    downs_0_d_payload_size;
  wire                downs_0_d_payload_denied;
  wire       [31:0]   downs_0_d_payload_data;
  wire                downs_0_d_payload_corrupt;
  wire                downs_1_a_valid;
  wire                downs_1_a_ready;
  wire       [2:0]    downs_1_a_payload_opcode;
  wire       [2:0]    downs_1_a_payload_param;
  wire       [2:0]    downs_1_a_payload_source;
  wire       [13:0]   downs_1_a_payload_address;
  wire       [2:0]    downs_1_a_payload_size;
  wire       [3:0]    downs_1_a_payload_mask;
  wire       [31:0]   downs_1_a_payload_data;
  wire                downs_1_a_payload_corrupt;
  wire                downs_1_d_valid;
  wire                downs_1_d_ready;
  wire       [2:0]    downs_1_d_payload_opcode;
  wire       [2:0]    downs_1_d_payload_param;
  wire       [2:0]    downs_1_d_payload_source;
  wire       [2:0]    downs_1_d_payload_size;
  wire                downs_1_d_payload_denied;
  wire       [31:0]   downs_1_d_payload_data;
  wire                downs_1_d_payload_corrupt;
  wire       [33:0]   a_key;
  wire                a_logic_0_hit;
  wire                a_logic_1_hit;
  wire                a_miss;
  `ifndef SYNTHESIS
  reg [127:0] io_up_a_payload_opcode_string;
  reg [119:0] io_up_d_payload_opcode_string;
  reg [127:0] io_downs_0_a_payload_opcode_string;
  reg [119:0] io_downs_0_d_payload_opcode_string;
  reg [127:0] io_downs_1_a_payload_opcode_string;
  reg [119:0] io_downs_1_d_payload_opcode_string;
  reg [127:0] downs_0_a_payload_opcode_string;
  reg [119:0] downs_0_d_payload_opcode_string;
  reg [127:0] downs_1_a_payload_opcode_string;
  reg [119:0] downs_1_d_payload_opcode_string;
  `endif


  assign _zz_a_logic_0_hit = (|((a_key & 34'h040000000) == 34'h0));
  assign _zz_downs_0_a_payload_address = (io_up_a_payload_address - 31'h0);
  assign _zz_a_logic_1_hit = (|((a_key & 34'h040000000) == 34'h040000000));
  assign _zz_downs_1_a_payload_address = (io_up_a_payload_address - 31'h40000000);
  assign _zz_2 = {io_downs_1_a_valid,io_downs_0_a_valid};
  StreamArbiter_8 d_arbiter (
    .io_inputs_0_valid           (downs_0_d_valid                        ), //i
    .io_inputs_0_ready           (d_arbiter_io_inputs_0_ready            ), //o
    .io_inputs_0_payload_opcode  (downs_0_d_payload_opcode[2:0]          ), //i
    .io_inputs_0_payload_param   (downs_0_d_payload_param[2:0]           ), //i
    .io_inputs_0_payload_source  (downs_0_d_payload_source[2:0]          ), //i
    .io_inputs_0_payload_size    (downs_0_d_payload_size[2:0]            ), //i
    .io_inputs_0_payload_denied  (downs_0_d_payload_denied               ), //i
    .io_inputs_0_payload_data    (downs_0_d_payload_data[31:0]           ), //i
    .io_inputs_0_payload_corrupt (downs_0_d_payload_corrupt              ), //i
    .io_inputs_1_valid           (downs_1_d_valid                        ), //i
    .io_inputs_1_ready           (d_arbiter_io_inputs_1_ready            ), //o
    .io_inputs_1_payload_opcode  (downs_1_d_payload_opcode[2:0]          ), //i
    .io_inputs_1_payload_param   (downs_1_d_payload_param[2:0]           ), //i
    .io_inputs_1_payload_source  (downs_1_d_payload_source[2:0]          ), //i
    .io_inputs_1_payload_size    (downs_1_d_payload_size[2:0]            ), //i
    .io_inputs_1_payload_denied  (downs_1_d_payload_denied               ), //i
    .io_inputs_1_payload_data    (downs_1_d_payload_data[31:0]           ), //i
    .io_inputs_1_payload_corrupt (downs_1_d_payload_corrupt              ), //i
    .io_output_valid             (d_arbiter_io_output_valid              ), //o
    .io_output_ready             (io_up_d_ready                          ), //i
    .io_output_payload_opcode    (d_arbiter_io_output_payload_opcode[2:0]), //o
    .io_output_payload_param     (d_arbiter_io_output_payload_param[2:0] ), //o
    .io_output_payload_source    (d_arbiter_io_output_payload_source[2:0]), //o
    .io_output_payload_size      (d_arbiter_io_output_payload_size[2:0]  ), //o
    .io_output_payload_denied    (d_arbiter_io_output_payload_denied     ), //o
    .io_output_payload_data      (d_arbiter_io_output_payload_data[31:0] ), //o
    .io_output_payload_corrupt   (d_arbiter_io_output_payload_corrupt    ), //o
    .io_chosen                   (d_arbiter_io_chosen                    ), //o
    .io_chosenOH                 (d_arbiter_io_chosenOH[1:0]             ), //o
    .clk_cpu                     (clk_cpu                                ), //i
    .reset_cpu                   (reset_cpu                              )  //i
  );
  always @(*) begin
    case(_zz_2)
      2'b00 : _zz_1 = 2'b00;
      2'b01 : _zz_1 = 2'b01;
      2'b10 : _zz_1 = 2'b01;
      default : _zz_1 = 2'b10;
    endcase
  end

  `ifndef SYNTHESIS
  always @(*) begin
    case(io_up_a_payload_opcode)
      A_PUT_FULL_DATA : io_up_a_payload_opcode_string = "PUT_FULL_DATA   ";
      A_PUT_PARTIAL_DATA : io_up_a_payload_opcode_string = "PUT_PARTIAL_DATA";
      A_GET : io_up_a_payload_opcode_string = "GET             ";
      A_ACQUIRE_BLOCK : io_up_a_payload_opcode_string = "ACQUIRE_BLOCK   ";
      A_ACQUIRE_PERM : io_up_a_payload_opcode_string = "ACQUIRE_PERM    ";
      default : io_up_a_payload_opcode_string = "????????????????";
    endcase
  end
  always @(*) begin
    case(io_up_d_payload_opcode)
      D_ACCESS_ACK : io_up_d_payload_opcode_string = "ACCESS_ACK     ";
      D_ACCESS_ACK_DATA : io_up_d_payload_opcode_string = "ACCESS_ACK_DATA";
      D_GRANT : io_up_d_payload_opcode_string = "GRANT          ";
      D_GRANT_DATA : io_up_d_payload_opcode_string = "GRANT_DATA     ";
      D_RELEASE_ACK : io_up_d_payload_opcode_string = "RELEASE_ACK    ";
      default : io_up_d_payload_opcode_string = "???????????????";
    endcase
  end
  always @(*) begin
    case(io_downs_0_a_payload_opcode)
      A_PUT_FULL_DATA : io_downs_0_a_payload_opcode_string = "PUT_FULL_DATA   ";
      A_PUT_PARTIAL_DATA : io_downs_0_a_payload_opcode_string = "PUT_PARTIAL_DATA";
      A_GET : io_downs_0_a_payload_opcode_string = "GET             ";
      A_ACQUIRE_BLOCK : io_downs_0_a_payload_opcode_string = "ACQUIRE_BLOCK   ";
      A_ACQUIRE_PERM : io_downs_0_a_payload_opcode_string = "ACQUIRE_PERM    ";
      default : io_downs_0_a_payload_opcode_string = "????????????????";
    endcase
  end
  always @(*) begin
    case(io_downs_0_d_payload_opcode)
      D_ACCESS_ACK : io_downs_0_d_payload_opcode_string = "ACCESS_ACK     ";
      D_ACCESS_ACK_DATA : io_downs_0_d_payload_opcode_string = "ACCESS_ACK_DATA";
      D_GRANT : io_downs_0_d_payload_opcode_string = "GRANT          ";
      D_GRANT_DATA : io_downs_0_d_payload_opcode_string = "GRANT_DATA     ";
      D_RELEASE_ACK : io_downs_0_d_payload_opcode_string = "RELEASE_ACK    ";
      default : io_downs_0_d_payload_opcode_string = "???????????????";
    endcase
  end
  always @(*) begin
    case(io_downs_1_a_payload_opcode)
      A_PUT_FULL_DATA : io_downs_1_a_payload_opcode_string = "PUT_FULL_DATA   ";
      A_PUT_PARTIAL_DATA : io_downs_1_a_payload_opcode_string = "PUT_PARTIAL_DATA";
      A_GET : io_downs_1_a_payload_opcode_string = "GET             ";
      A_ACQUIRE_BLOCK : io_downs_1_a_payload_opcode_string = "ACQUIRE_BLOCK   ";
      A_ACQUIRE_PERM : io_downs_1_a_payload_opcode_string = "ACQUIRE_PERM    ";
      default : io_downs_1_a_payload_opcode_string = "????????????????";
    endcase
  end
  always @(*) begin
    case(io_downs_1_d_payload_opcode)
      D_ACCESS_ACK : io_downs_1_d_payload_opcode_string = "ACCESS_ACK     ";
      D_ACCESS_ACK_DATA : io_downs_1_d_payload_opcode_string = "ACCESS_ACK_DATA";
      D_GRANT : io_downs_1_d_payload_opcode_string = "GRANT          ";
      D_GRANT_DATA : io_downs_1_d_payload_opcode_string = "GRANT_DATA     ";
      D_RELEASE_ACK : io_downs_1_d_payload_opcode_string = "RELEASE_ACK    ";
      default : io_downs_1_d_payload_opcode_string = "???????????????";
    endcase
  end
  always @(*) begin
    case(downs_0_a_payload_opcode)
      A_PUT_FULL_DATA : downs_0_a_payload_opcode_string = "PUT_FULL_DATA   ";
      A_PUT_PARTIAL_DATA : downs_0_a_payload_opcode_string = "PUT_PARTIAL_DATA";
      A_GET : downs_0_a_payload_opcode_string = "GET             ";
      A_ACQUIRE_BLOCK : downs_0_a_payload_opcode_string = "ACQUIRE_BLOCK   ";
      A_ACQUIRE_PERM : downs_0_a_payload_opcode_string = "ACQUIRE_PERM    ";
      default : downs_0_a_payload_opcode_string = "????????????????";
    endcase
  end
  always @(*) begin
    case(downs_0_d_payload_opcode)
      D_ACCESS_ACK : downs_0_d_payload_opcode_string = "ACCESS_ACK     ";
      D_ACCESS_ACK_DATA : downs_0_d_payload_opcode_string = "ACCESS_ACK_DATA";
      D_GRANT : downs_0_d_payload_opcode_string = "GRANT          ";
      D_GRANT_DATA : downs_0_d_payload_opcode_string = "GRANT_DATA     ";
      D_RELEASE_ACK : downs_0_d_payload_opcode_string = "RELEASE_ACK    ";
      default : downs_0_d_payload_opcode_string = "???????????????";
    endcase
  end
  always @(*) begin
    case(downs_1_a_payload_opcode)
      A_PUT_FULL_DATA : downs_1_a_payload_opcode_string = "PUT_FULL_DATA   ";
      A_PUT_PARTIAL_DATA : downs_1_a_payload_opcode_string = "PUT_PARTIAL_DATA";
      A_GET : downs_1_a_payload_opcode_string = "GET             ";
      A_ACQUIRE_BLOCK : downs_1_a_payload_opcode_string = "ACQUIRE_BLOCK   ";
      A_ACQUIRE_PERM : downs_1_a_payload_opcode_string = "ACQUIRE_PERM    ";
      default : downs_1_a_payload_opcode_string = "????????????????";
    endcase
  end
  always @(*) begin
    case(downs_1_d_payload_opcode)
      D_ACCESS_ACK : downs_1_d_payload_opcode_string = "ACCESS_ACK     ";
      D_ACCESS_ACK_DATA : downs_1_d_payload_opcode_string = "ACCESS_ACK_DATA";
      D_GRANT : downs_1_d_payload_opcode_string = "GRANT          ";
      D_GRANT_DATA : downs_1_d_payload_opcode_string = "GRANT_DATA     ";
      D_RELEASE_ACK : downs_1_d_payload_opcode_string = "RELEASE_ACK    ";
      default : downs_1_d_payload_opcode_string = "???????????????";
    endcase
  end
  `endif

  assign io_downs_0_a_valid = downs_0_a_valid;
  assign downs_0_a_ready = io_downs_0_a_ready;
  assign io_downs_0_a_payload_opcode = downs_0_a_payload_opcode;
  assign io_downs_0_a_payload_param = downs_0_a_payload_param;
  assign io_downs_0_a_payload_source = downs_0_a_payload_source;
  assign io_downs_0_a_payload_address = downs_0_a_payload_address;
  assign io_downs_0_a_payload_size = downs_0_a_payload_size;
  assign io_downs_0_a_payload_mask = downs_0_a_payload_mask;
  assign io_downs_0_a_payload_data = downs_0_a_payload_data;
  assign io_downs_0_a_payload_corrupt = downs_0_a_payload_corrupt;
  assign downs_0_d_valid = io_downs_0_d_valid;
  assign io_downs_0_d_ready = downs_0_d_ready;
  assign downs_0_d_payload_opcode = io_downs_0_d_payload_opcode;
  assign downs_0_d_payload_param = io_downs_0_d_payload_param;
  assign downs_0_d_payload_source = io_downs_0_d_payload_source;
  assign downs_0_d_payload_size = io_downs_0_d_payload_size;
  assign downs_0_d_payload_denied = io_downs_0_d_payload_denied;
  assign downs_0_d_payload_data = io_downs_0_d_payload_data;
  assign downs_0_d_payload_corrupt = io_downs_0_d_payload_corrupt;
  assign io_downs_1_a_valid = downs_1_a_valid;
  assign downs_1_a_ready = io_downs_1_a_ready;
  assign io_downs_1_a_payload_opcode = downs_1_a_payload_opcode;
  assign io_downs_1_a_payload_param = downs_1_a_payload_param;
  assign io_downs_1_a_payload_source = downs_1_a_payload_source;
  assign io_downs_1_a_payload_address = downs_1_a_payload_address;
  assign io_downs_1_a_payload_size = downs_1_a_payload_size;
  assign io_downs_1_a_payload_mask = downs_1_a_payload_mask;
  assign io_downs_1_a_payload_data = downs_1_a_payload_data;
  assign io_downs_1_a_payload_corrupt = downs_1_a_payload_corrupt;
  assign downs_1_d_valid = io_downs_1_d_valid;
  assign io_downs_1_d_ready = downs_1_d_ready;
  assign downs_1_d_payload_opcode = io_downs_1_d_payload_opcode;
  assign downs_1_d_payload_param = io_downs_1_d_payload_param;
  assign downs_1_d_payload_source = io_downs_1_d_payload_source;
  assign downs_1_d_payload_size = io_downs_1_d_payload_size;
  assign downs_1_d_payload_denied = io_downs_1_d_payload_denied;
  assign downs_1_d_payload_data = io_downs_1_d_payload_data;
  assign downs_1_d_payload_corrupt = io_downs_1_d_payload_corrupt;
  assign a_key = {io_up_a_payload_opcode,io_up_a_payload_address};
  assign a_logic_0_hit = _zz_a_logic_0_hit[0];
  assign downs_0_a_valid = (io_up_a_valid && a_logic_0_hit);
  assign downs_0_a_payload_opcode = io_up_a_payload_opcode;
  assign downs_0_a_payload_param = io_up_a_payload_param;
  assign downs_0_a_payload_source = io_up_a_payload_source;
  assign downs_0_a_payload_mask = io_up_a_payload_mask;
  assign downs_0_a_payload_data = io_up_a_payload_data;
  assign downs_0_a_payload_corrupt = io_up_a_payload_corrupt;
  assign downs_0_a_payload_address = _zz_downs_0_a_payload_address[26:0];
  assign downs_0_a_payload_size = io_up_a_payload_size;
  assign a_logic_1_hit = _zz_a_logic_1_hit[0];
  assign downs_1_a_valid = (io_up_a_valid && a_logic_1_hit);
  assign downs_1_a_payload_opcode = io_up_a_payload_opcode;
  assign downs_1_a_payload_param = io_up_a_payload_param;
  assign downs_1_a_payload_source = io_up_a_payload_source;
  assign downs_1_a_payload_mask = io_up_a_payload_mask;
  assign downs_1_a_payload_data = io_up_a_payload_data;
  assign downs_1_a_payload_corrupt = io_up_a_payload_corrupt;
  assign downs_1_a_payload_address = _zz_downs_1_a_payload_address[13:0];
  assign downs_1_a_payload_size = io_up_a_payload_size;
  assign io_up_a_ready = (|{(downs_1_a_ready && a_logic_1_hit),(downs_0_a_ready && a_logic_0_hit)});
  assign a_miss = (! (|{a_logic_1_hit,a_logic_0_hit}));
  assign downs_0_d_ready = d_arbiter_io_inputs_0_ready;
  assign downs_1_d_ready = d_arbiter_io_inputs_1_ready;
  assign io_up_d_valid = d_arbiter_io_output_valid;
  assign io_up_d_payload_opcode = d_arbiter_io_output_payload_opcode;
  assign io_up_d_payload_param = d_arbiter_io_output_payload_param;
  assign io_up_d_payload_source = d_arbiter_io_output_payload_source;
  assign io_up_d_payload_size = d_arbiter_io_output_payload_size;
  assign io_up_d_payload_denied = d_arbiter_io_output_payload_denied;
  assign io_up_d_payload_data = d_arbiter_io_output_payload_data;
  assign io_up_d_payload_corrupt = d_arbiter_io_output_payload_corrupt;
  always @(posedge clk_cpu or posedge reset_cpu) begin
    if(reset_cpu) begin
    end else begin
      `ifndef SYNTHESIS
        `ifdef FORMAL
          assert((! (io_up_a_valid && a_miss))); // Decoder.scala:L106
        `else
          if(!(! (io_up_a_valid && a_miss))) begin
            $display("FAILURE Tilelink decoder miss ???"); // Decoder.scala:L106
            $finish;
          end
        `endif
      `endif
      `ifndef SYNTHESIS
        `ifdef FORMAL
          assert((! (io_up_a_valid && (_zz_1 != 2'b01)))); // Decoder.scala:L107
        `else
          if(!(! (io_up_a_valid && (_zz_1 != 2'b01)))) begin
            $display("FAILURE Tilelink decoder miss ???"); // Decoder.scala:L107
            $finish;
          end
        `endif
      `endif
    end
  end


endmodule

module WidthAdapter_1 (
  input  wire          io_up_a_valid,
  output wire          io_up_a_ready,
  input  wire [2:0]    io_up_a_payload_opcode,
  input  wire [2:0]    io_up_a_payload_param,
  input  wire [2:0]    io_up_a_payload_source,
  input  wire [30:0]   io_up_a_payload_address,
  input  wire [2:0]    io_up_a_payload_size,
  input  wire [7:0]    io_up_a_payload_mask,
  input  wire [63:0]   io_up_a_payload_data,
  input  wire          io_up_a_payload_corrupt,
  output wire          io_up_d_valid,
  input  wire          io_up_d_ready,
  output wire [2:0]    io_up_d_payload_opcode,
  output wire [2:0]    io_up_d_payload_param,
  output wire [2:0]    io_up_d_payload_source,
  output wire [2:0]    io_up_d_payload_size,
  output wire          io_up_d_payload_denied,
  output wire [63:0]   io_up_d_payload_data,
  output wire          io_up_d_payload_corrupt,
  output wire          io_down_a_valid,
  input  wire          io_down_a_ready,
  output wire [2:0]    io_down_a_payload_opcode,
  output wire [2:0]    io_down_a_payload_param,
  output wire [2:0]    io_down_a_payload_source,
  output reg  [30:0]   io_down_a_payload_address,
  output wire [2:0]    io_down_a_payload_size,
  output wire [3:0]    io_down_a_payload_mask,
  output wire [31:0]   io_down_a_payload_data,
  output wire          io_down_a_payload_corrupt,
  input  wire          io_down_d_valid,
  output wire          io_down_d_ready,
  input  wire [2:0]    io_down_d_payload_opcode,
  input  wire [2:0]    io_down_d_payload_param,
  input  wire [2:0]    io_down_d_payload_source,
  input  wire [2:0]    io_down_d_payload_size,
  input  wire          io_down_d_payload_denied,
  input  wire [31:0]   io_down_d_payload_data,
  input  wire          io_down_d_payload_corrupt,
  input  wire          clk_cpu,
  input  wire          reset_cpu
);
  localparam A_PUT_FULL_DATA = 3'd0;
  localparam A_PUT_PARTIAL_DATA = 3'd1;
  localparam A_GET = 3'd4;
  localparam A_ACQUIRE_BLOCK = 3'd6;
  localparam A_ACQUIRE_PERM = 3'd7;
  localparam D_ACCESS_ACK = 3'd0;
  localparam D_ACCESS_ACK_DATA = 3'd1;
  localparam D_GRANT = 3'd4;
  localparam D_GRANT_DATA = 3'd5;
  localparam D_RELEASE_ACK = 3'd6;

  reg        [3:0]    _zz_downsize_a_ctrl_burstLast;
  reg        [31:0]   _zz_io_down_a_payload_data;
  reg        [3:0]    _zz_io_down_a_payload_mask;
  reg        [3:0]    _zz_downsize_d_ctrl_burstLast;
  reg        [0:0]    downsize_a_ctrl_counter;
  wire       [0:0]    downsize_a_ctrl_sel;
  reg        [3:0]    io_down_a_tracker_beat;
  wire                downsize_a_ctrl_burstLast;
  wire                io_down_a_fire;
  reg        [3:0]    io_down_d_tracker_beat;
  wire                downsize_d_ctrl_burstLast;
  wire                io_down_d_fire;
  wire       [0:0]    downsize_d_sel;
  wire                downsize_d_ctrl_wordLast;
  reg                 downsize_d_ctrl_buffer_valid;
  reg                 downsize_d_ctrl_buffer_first;
  reg        [2:0]    downsize_d_ctrl_buffer_args_opcode;
  reg        [2:0]    downsize_d_ctrl_buffer_args_param;
  reg        [2:0]    downsize_d_ctrl_buffer_args_source;
  reg        [30:0]   downsize_d_ctrl_buffer_args_address;
  reg        [2:0]    downsize_d_ctrl_buffer_args_size;
  reg        [31:0]   downsize_d_ctrl_buffer_data_0;
  reg        [31:0]   downsize_d_ctrl_buffer_data_1;
  reg                 downsize_d_ctrl_buffer_corrupt;
  reg                 downsize_d_ctrl_buffer_denied;
  wire       [0:0]    _zz_when_WidthAdapter_l84;
  wire                when_WidthAdapter_l84;
  wire                when_WidthAdapter_l84_1;
  `ifndef SYNTHESIS
  reg [127:0] io_up_a_payload_opcode_string;
  reg [119:0] io_up_d_payload_opcode_string;
  reg [127:0] io_down_a_payload_opcode_string;
  reg [119:0] io_down_d_payload_opcode_string;
  reg [127:0] downsize_d_ctrl_buffer_args_opcode_string;
  `endif


  always @(*) begin
    case(io_down_a_payload_size)
      3'b000 : _zz_downsize_a_ctrl_burstLast = 4'b0000;
      3'b001 : _zz_downsize_a_ctrl_burstLast = 4'b0000;
      3'b010 : _zz_downsize_a_ctrl_burstLast = 4'b0000;
      3'b011 : _zz_downsize_a_ctrl_burstLast = 4'b0001;
      3'b100 : _zz_downsize_a_ctrl_burstLast = 4'b0011;
      3'b101 : _zz_downsize_a_ctrl_burstLast = 4'b0111;
      default : _zz_downsize_a_ctrl_burstLast = 4'b1111;
    endcase
  end

  always @(*) begin
    case(downsize_a_ctrl_sel)
      1'b0 : begin
        _zz_io_down_a_payload_data = io_up_a_payload_data[31 : 0];
        _zz_io_down_a_payload_mask = io_up_a_payload_mask[3 : 0];
      end
      default : begin
        _zz_io_down_a_payload_data = io_up_a_payload_data[63 : 32];
        _zz_io_down_a_payload_mask = io_up_a_payload_mask[7 : 4];
      end
    endcase
  end

  always @(*) begin
    case(io_down_d_payload_size)
      3'b000 : _zz_downsize_d_ctrl_burstLast = 4'b0000;
      3'b001 : _zz_downsize_d_ctrl_burstLast = 4'b0000;
      3'b010 : _zz_downsize_d_ctrl_burstLast = 4'b0000;
      3'b011 : _zz_downsize_d_ctrl_burstLast = 4'b0001;
      3'b100 : _zz_downsize_d_ctrl_burstLast = 4'b0011;
      3'b101 : _zz_downsize_d_ctrl_burstLast = 4'b0111;
      default : _zz_downsize_d_ctrl_burstLast = 4'b1111;
    endcase
  end

  `ifndef SYNTHESIS
  always @(*) begin
    case(io_up_a_payload_opcode)
      A_PUT_FULL_DATA : io_up_a_payload_opcode_string = "PUT_FULL_DATA   ";
      A_PUT_PARTIAL_DATA : io_up_a_payload_opcode_string = "PUT_PARTIAL_DATA";
      A_GET : io_up_a_payload_opcode_string = "GET             ";
      A_ACQUIRE_BLOCK : io_up_a_payload_opcode_string = "ACQUIRE_BLOCK   ";
      A_ACQUIRE_PERM : io_up_a_payload_opcode_string = "ACQUIRE_PERM    ";
      default : io_up_a_payload_opcode_string = "????????????????";
    endcase
  end
  always @(*) begin
    case(io_up_d_payload_opcode)
      D_ACCESS_ACK : io_up_d_payload_opcode_string = "ACCESS_ACK     ";
      D_ACCESS_ACK_DATA : io_up_d_payload_opcode_string = "ACCESS_ACK_DATA";
      D_GRANT : io_up_d_payload_opcode_string = "GRANT          ";
      D_GRANT_DATA : io_up_d_payload_opcode_string = "GRANT_DATA     ";
      D_RELEASE_ACK : io_up_d_payload_opcode_string = "RELEASE_ACK    ";
      default : io_up_d_payload_opcode_string = "???????????????";
    endcase
  end
  always @(*) begin
    case(io_down_a_payload_opcode)
      A_PUT_FULL_DATA : io_down_a_payload_opcode_string = "PUT_FULL_DATA   ";
      A_PUT_PARTIAL_DATA : io_down_a_payload_opcode_string = "PUT_PARTIAL_DATA";
      A_GET : io_down_a_payload_opcode_string = "GET             ";
      A_ACQUIRE_BLOCK : io_down_a_payload_opcode_string = "ACQUIRE_BLOCK   ";
      A_ACQUIRE_PERM : io_down_a_payload_opcode_string = "ACQUIRE_PERM    ";
      default : io_down_a_payload_opcode_string = "????????????????";
    endcase
  end
  always @(*) begin
    case(io_down_d_payload_opcode)
      D_ACCESS_ACK : io_down_d_payload_opcode_string = "ACCESS_ACK     ";
      D_ACCESS_ACK_DATA : io_down_d_payload_opcode_string = "ACCESS_ACK_DATA";
      D_GRANT : io_down_d_payload_opcode_string = "GRANT          ";
      D_GRANT_DATA : io_down_d_payload_opcode_string = "GRANT_DATA     ";
      D_RELEASE_ACK : io_down_d_payload_opcode_string = "RELEASE_ACK    ";
      default : io_down_d_payload_opcode_string = "???????????????";
    endcase
  end
  always @(*) begin
    case(downsize_d_ctrl_buffer_args_opcode)
      A_PUT_FULL_DATA : downsize_d_ctrl_buffer_args_opcode_string = "PUT_FULL_DATA   ";
      A_PUT_PARTIAL_DATA : downsize_d_ctrl_buffer_args_opcode_string = "PUT_PARTIAL_DATA";
      A_GET : downsize_d_ctrl_buffer_args_opcode_string = "GET             ";
      A_ACQUIRE_BLOCK : downsize_d_ctrl_buffer_args_opcode_string = "ACQUIRE_BLOCK   ";
      A_ACQUIRE_PERM : downsize_d_ctrl_buffer_args_opcode_string = "ACQUIRE_PERM    ";
      default : downsize_d_ctrl_buffer_args_opcode_string = "????????????????";
    endcase
  end
  `endif

  assign downsize_a_ctrl_sel = (downsize_a_ctrl_counter + io_up_a_payload_address[2 : 2]);
  assign downsize_a_ctrl_burstLast = ((! ((1'b0 || (A_PUT_FULL_DATA == io_down_a_payload_opcode)) || (A_PUT_PARTIAL_DATA == io_down_a_payload_opcode))) || (io_down_a_tracker_beat == _zz_downsize_a_ctrl_burstLast));
  assign io_down_a_fire = (io_down_a_valid && io_down_a_ready);
  assign io_down_a_valid = io_up_a_valid;
  assign io_down_a_payload_opcode = io_up_a_payload_opcode;
  assign io_down_a_payload_param = io_up_a_payload_param;
  assign io_down_a_payload_source = io_up_a_payload_source;
  always @(*) begin
    io_down_a_payload_address = io_up_a_payload_address;
    io_down_a_payload_address[2 : 2] = downsize_a_ctrl_sel;
  end

  assign io_down_a_payload_size = io_up_a_payload_size;
  assign io_down_a_payload_corrupt = io_up_a_payload_corrupt;
  assign io_up_a_ready = (io_down_a_ready && ((&downsize_a_ctrl_counter) || downsize_a_ctrl_burstLast));
  assign io_down_a_payload_data = _zz_io_down_a_payload_data;
  assign io_down_a_payload_mask = _zz_io_down_a_payload_mask;
  assign downsize_d_ctrl_burstLast = ((! ((1'b0 || (D_ACCESS_ACK_DATA == io_down_d_payload_opcode)) || (D_GRANT_DATA == io_down_d_payload_opcode))) || (io_down_d_tracker_beat == _zz_downsize_d_ctrl_burstLast));
  assign io_down_d_fire = (io_down_d_valid && io_down_d_ready);
  assign downsize_d_sel = io_down_d_tracker_beat[0:0];
  assign downsize_d_ctrl_wordLast = ((&downsize_d_sel) || downsize_d_ctrl_burstLast);
  assign io_up_d_valid = downsize_d_ctrl_buffer_valid;
  assign io_up_d_payload_opcode = downsize_d_ctrl_buffer_args_opcode;
  assign io_up_d_payload_param = downsize_d_ctrl_buffer_args_param;
  assign io_up_d_payload_source = downsize_d_ctrl_buffer_args_source;
  assign io_up_d_payload_size = downsize_d_ctrl_buffer_args_size;
  assign io_up_d_payload_data = {downsize_d_ctrl_buffer_data_1,downsize_d_ctrl_buffer_data_0};
  assign io_up_d_payload_corrupt = downsize_d_ctrl_buffer_corrupt;
  assign io_up_d_payload_denied = downsize_d_ctrl_buffer_denied;
  assign io_down_d_ready = ((! downsize_d_ctrl_buffer_valid) || io_up_d_ready);
  assign _zz_when_WidthAdapter_l84 = (3'b011 <= io_down_d_payload_size);
  assign when_WidthAdapter_l84 = (((downsize_d_sel ^ 1'b0) & _zz_when_WidthAdapter_l84) == 1'b0);
  assign when_WidthAdapter_l84_1 = (((downsize_d_sel ^ 1'b1) & _zz_when_WidthAdapter_l84) == 1'b0);
  always @(posedge clk_cpu or posedge reset_cpu) begin
    if(reset_cpu) begin
      downsize_a_ctrl_counter <= 1'b0;
      io_down_a_tracker_beat <= 4'b0000;
      io_down_d_tracker_beat <= 4'b0000;
      downsize_d_ctrl_buffer_valid <= 1'b0;
      downsize_d_ctrl_buffer_first <= 1'b1;
    end else begin
      if(io_down_a_fire) begin
        io_down_a_tracker_beat <= (io_down_a_tracker_beat + 4'b0001);
        if(downsize_a_ctrl_burstLast) begin
          io_down_a_tracker_beat <= 4'b0000;
        end
      end
      if(io_down_a_fire) begin
        downsize_a_ctrl_counter <= (downsize_a_ctrl_counter + 1'b1);
        if(downsize_a_ctrl_burstLast) begin
          downsize_a_ctrl_counter <= 1'b0;
        end
      end
      if(io_down_d_fire) begin
        io_down_d_tracker_beat <= (io_down_d_tracker_beat + 4'b0001);
        if(downsize_d_ctrl_burstLast) begin
          io_down_d_tracker_beat <= 4'b0000;
        end
      end
      if(io_up_d_ready) begin
        downsize_d_ctrl_buffer_valid <= 1'b0;
      end
      if(io_down_d_fire) begin
        downsize_d_ctrl_buffer_valid <= downsize_d_ctrl_wordLast;
        downsize_d_ctrl_buffer_first <= downsize_d_ctrl_wordLast;
      end
    end
  end

  always @(posedge clk_cpu) begin
    if(io_down_d_fire) begin
      if(downsize_d_ctrl_buffer_first) begin
        downsize_d_ctrl_buffer_args_opcode <= io_down_d_payload_opcode;
        downsize_d_ctrl_buffer_args_param <= io_down_d_payload_param;
        downsize_d_ctrl_buffer_args_source <= io_down_d_payload_source;
        downsize_d_ctrl_buffer_args_size <= io_down_d_payload_size;
        downsize_d_ctrl_buffer_corrupt <= 1'b0;
        downsize_d_ctrl_buffer_denied <= 1'b0;
      end
      if(when_WidthAdapter_l84) begin
        downsize_d_ctrl_buffer_data_0 <= io_down_d_payload_data;
      end
      if(when_WidthAdapter_l84_1) begin
        downsize_d_ctrl_buffer_data_1 <= io_down_d_payload_data;
      end
      if(io_down_d_payload_corrupt) begin
        downsize_d_ctrl_buffer_corrupt <= 1'b1;
      end
      if(io_down_d_payload_denied) begin
        downsize_d_ctrl_buffer_denied <= 1'b1;
      end
    end
  end


endmodule

module Ram (
  input  wire          io_up_a_valid,
  output reg           io_up_a_ready,
  input  wire [2:0]    io_up_a_payload_opcode,
  input  wire [2:0]    io_up_a_payload_param,
  input  wire [2:0]    io_up_a_payload_source,
  input  wire [13:0]   io_up_a_payload_address,
  input  wire [2:0]    io_up_a_payload_size,
  input  wire [3:0]    io_up_a_payload_mask,
  input  wire [31:0]   io_up_a_payload_data,
  input  wire          io_up_a_payload_corrupt,
  output wire          io_up_d_valid,
  input  wire          io_up_d_ready,
  output wire [2:0]    io_up_d_payload_opcode,
  output wire [2:0]    io_up_d_payload_param,
  output wire [2:0]    io_up_d_payload_source,
  output wire [2:0]    io_up_d_payload_size,
  output wire          io_up_d_payload_denied,
  output wire [31:0]   io_up_d_payload_data,
  output wire          io_up_d_payload_corrupt,
  input  wire          clk_cpu,
  input  wire          reset_cpu
);
  localparam A_PUT_FULL_DATA = 3'd0;
  localparam A_PUT_PARTIAL_DATA = 3'd1;
  localparam A_GET = 3'd4;
  localparam A_ACQUIRE_BLOCK = 3'd6;
  localparam A_ACQUIRE_PERM = 3'd7;
  localparam D_ACCESS_ACK = 3'd0;
  localparam D_ACCESS_ACK_DATA = 3'd1;
  localparam D_GRANT = 3'd4;
  localparam D_GRANT_DATA = 3'd5;
  localparam D_RELEASE_ACK = 3'd6;

  wire                mem_en;
  wire       [31:0]   mem_rdData;
  reg        [3:0]    _zz_when_Ram_l54;
  wire       [11:0]   _zz_port_address;
  reg        [3:0]    _zz_io_up_a_tracker_last;
  wire       [7:0]    _zz_ordering_payload_bytes;
  reg                 pipeline_rsp_ready;
  reg        [2:0]    pipeline_rsp_cmd_SIZE;
  reg        [2:0]    pipeline_rsp_cmd_SOURCE;
  reg                 pipeline_rsp_cmd_IS_GET;
  reg                 pipeline_rsp_cmd_LAST;
  wire                pipeline_cmd_ready;
  reg                 pipeline_cmd_LAST;
  reg        [2:0]    pipeline_cmd_SOURCE;
  reg        [2:0]    pipeline_cmd_SIZE;
  reg                 pipeline_cmd_IS_GET;
  wire       [11:0]   port_address;
  wire       [31:0]   port_rdata;
  wire       [31:0]   port_wdata;
  wire                port_enable;
  wire                port_write;
  wire       [3:0]    port_mask;
  reg                 pipeline_cmd_valid;
  wire       [11:0]   pipeline_cmd_addressShifted;
  wire                pipeline_cmd_isFireing;
  reg        [3:0]    pipeline_cmd_fsm_counter;
  reg        [11:0]   pipeline_cmd_fsm_address;
  reg        [2:0]    pipeline_cmd_fsm_size;
  reg        [2:0]    pipeline_cmd_fsm_source;
  reg                 pipeline_cmd_fsm_isGet;
  wire                pipeline_cmd_fsm_busy;
  wire                when_Ram_l42;
  wire                io_up_a_fire;
  wire                when_Ram_l47;
  wire                when_Ram_l54;
  reg                 pipeline_rsp_valid;
  wire                pipeline_rsp_takeIt;
  wire                pipeline_rsp_haltRequest_Ram_l73;
  wire       [2:0]    _zz_io_up_d_payload_opcode;
  reg                 pipeline_cmd_ready_output;
  wire                when_Pipeline_l278;
  wire                when_Connection_l74;
  wire                ordering_valid;
  wire       [6:0]    ordering_payload_bytes;
  reg        [3:0]    io_up_a_tracker_beat;
  wire                io_up_a_tracker_last;
  reg                 ordering_regNext_valid;
  reg        [6:0]    ordering_regNext_payload_bytes;
  `ifndef SYNTHESIS
  reg [127:0] io_up_a_payload_opcode_string;
  reg [119:0] io_up_d_payload_opcode_string;
  reg [119:0] _zz_io_up_d_payload_opcode_string;
  `endif


  assign _zz_port_address = {8'd0, pipeline_cmd_fsm_counter};
  assign _zz_ordering_payload_bytes = ({7'd0,1'b1} <<< io_up_a_payload_size);
  Ram_1wrs #(
    .wordCount      (4096      ),
    .wordWidth      (32        ),
    .readUnderWrite ("dontCare"),
    .duringWrite    ("dontCare"),
    .technology     ("auto"    ),
    .maskWidth      (4         ),
    .maskEnable     (1'b1      )
  ) mem (
    .clk    (clk_cpu           ), //i
    .en     (mem_en            ), //i
    .wr     (port_write        ), //i
    .addr   (port_address[11:0]), //i
    .mask   (port_mask[3:0]    ), //i
    .wrData (port_wdata[31:0]  ), //i
    .rdData (mem_rdData[31:0]  )  //o
  );
  always @(*) begin
    case(pipeline_cmd_SIZE)
      3'b000 : _zz_when_Ram_l54 = 4'b0000;
      3'b001 : _zz_when_Ram_l54 = 4'b0000;
      3'b010 : _zz_when_Ram_l54 = 4'b0000;
      3'b011 : _zz_when_Ram_l54 = 4'b0001;
      3'b100 : _zz_when_Ram_l54 = 4'b0011;
      3'b101 : _zz_when_Ram_l54 = 4'b0111;
      default : _zz_when_Ram_l54 = 4'b1111;
    endcase
  end

  always @(*) begin
    case(io_up_a_payload_size)
      3'b000 : _zz_io_up_a_tracker_last = 4'b0000;
      3'b001 : _zz_io_up_a_tracker_last = 4'b0000;
      3'b010 : _zz_io_up_a_tracker_last = 4'b0000;
      3'b011 : _zz_io_up_a_tracker_last = 4'b0001;
      3'b100 : _zz_io_up_a_tracker_last = 4'b0011;
      3'b101 : _zz_io_up_a_tracker_last = 4'b0111;
      default : _zz_io_up_a_tracker_last = 4'b1111;
    endcase
  end

  `ifndef SYNTHESIS
  always @(*) begin
    case(io_up_a_payload_opcode)
      A_PUT_FULL_DATA : io_up_a_payload_opcode_string = "PUT_FULL_DATA   ";
      A_PUT_PARTIAL_DATA : io_up_a_payload_opcode_string = "PUT_PARTIAL_DATA";
      A_GET : io_up_a_payload_opcode_string = "GET             ";
      A_ACQUIRE_BLOCK : io_up_a_payload_opcode_string = "ACQUIRE_BLOCK   ";
      A_ACQUIRE_PERM : io_up_a_payload_opcode_string = "ACQUIRE_PERM    ";
      default : io_up_a_payload_opcode_string = "????????????????";
    endcase
  end
  always @(*) begin
    case(io_up_d_payload_opcode)
      D_ACCESS_ACK : io_up_d_payload_opcode_string = "ACCESS_ACK     ";
      D_ACCESS_ACK_DATA : io_up_d_payload_opcode_string = "ACCESS_ACK_DATA";
      D_GRANT : io_up_d_payload_opcode_string = "GRANT          ";
      D_GRANT_DATA : io_up_d_payload_opcode_string = "GRANT_DATA     ";
      D_RELEASE_ACK : io_up_d_payload_opcode_string = "RELEASE_ACK    ";
      default : io_up_d_payload_opcode_string = "???????????????";
    endcase
  end
  always @(*) begin
    case(_zz_io_up_d_payload_opcode)
      D_ACCESS_ACK : _zz_io_up_d_payload_opcode_string = "ACCESS_ACK     ";
      D_ACCESS_ACK_DATA : _zz_io_up_d_payload_opcode_string = "ACCESS_ACK_DATA";
      D_GRANT : _zz_io_up_d_payload_opcode_string = "GRANT          ";
      D_GRANT_DATA : _zz_io_up_d_payload_opcode_string = "GRANT_DATA     ";
      D_RELEASE_ACK : _zz_io_up_d_payload_opcode_string = "RELEASE_ACK    ";
      default : _zz_io_up_d_payload_opcode_string = "???????????????";
    endcase
  end
  `endif

  assign port_rdata = mem_rdData;
  always @(*) begin
    pipeline_cmd_IS_GET = (|(io_up_a_payload_opcode == A_GET));
    if(pipeline_cmd_fsm_busy) begin
      pipeline_cmd_IS_GET = pipeline_cmd_fsm_isGet;
    end
  end

  always @(*) begin
    pipeline_cmd_SIZE = io_up_a_payload_size;
    if(pipeline_cmd_fsm_busy) begin
      pipeline_cmd_SIZE = pipeline_cmd_fsm_size;
    end
  end

  always @(*) begin
    pipeline_cmd_SOURCE = io_up_a_payload_source;
    if(pipeline_cmd_fsm_busy) begin
      pipeline_cmd_SOURCE = pipeline_cmd_fsm_source;
    end
  end

  always @(*) begin
    pipeline_cmd_LAST = 1'b1;
    if(when_Ram_l54) begin
      pipeline_cmd_LAST = 1'b0;
    end
  end

  always @(*) begin
    pipeline_cmd_valid = io_up_a_valid;
    if(when_Ram_l42) begin
      pipeline_cmd_valid = 1'b1;
    end
  end

  always @(*) begin
    io_up_a_ready = pipeline_cmd_ready;
    if(when_Ram_l42) begin
      io_up_a_ready = 1'b0;
    end
  end

  assign pipeline_cmd_addressShifted = (io_up_a_payload_address >>> 2'd2);
  assign pipeline_cmd_isFireing = (pipeline_cmd_valid && pipeline_cmd_ready);
  assign port_enable = pipeline_cmd_isFireing;
  assign port_write = (! pipeline_cmd_IS_GET);
  assign port_wdata = io_up_a_payload_data;
  assign port_mask = io_up_a_payload_mask;
  assign pipeline_cmd_fsm_busy = (pipeline_cmd_fsm_counter != 4'b0000);
  assign when_Ram_l42 = (pipeline_cmd_fsm_busy && pipeline_cmd_fsm_isGet);
  assign io_up_a_fire = (io_up_a_valid && io_up_a_ready);
  assign when_Ram_l47 = (io_up_a_fire && (! pipeline_cmd_fsm_busy));
  assign when_Ram_l54 = (pipeline_cmd_fsm_counter != _zz_when_Ram_l54);
  assign port_address = ((pipeline_cmd_fsm_busy ? pipeline_cmd_fsm_address : pipeline_cmd_addressShifted) | _zz_port_address);
  assign pipeline_rsp_takeIt = (pipeline_rsp_cmd_LAST || pipeline_rsp_cmd_IS_GET);
  assign pipeline_rsp_haltRequest_Ram_l73 = ((! io_up_d_ready) && pipeline_rsp_takeIt);
  assign io_up_d_valid = (pipeline_rsp_valid && pipeline_rsp_takeIt);
  assign _zz_io_up_d_payload_opcode = (pipeline_rsp_cmd_IS_GET ? D_ACCESS_ACK_DATA : D_ACCESS_ACK);
  assign io_up_d_payload_opcode = _zz_io_up_d_payload_opcode;
  assign io_up_d_payload_param = 3'b000;
  assign io_up_d_payload_source = pipeline_rsp_cmd_SOURCE;
  assign io_up_d_payload_size = pipeline_rsp_cmd_SIZE;
  assign io_up_d_payload_denied = 1'b0;
  assign io_up_d_payload_corrupt = 1'b0;
  assign io_up_d_payload_data = port_rdata;
  assign pipeline_cmd_ready = pipeline_cmd_ready_output;
  always @(*) begin
    pipeline_rsp_ready = 1'b1;
    if(when_Pipeline_l278) begin
      pipeline_rsp_ready = 1'b0;
    end
  end

  assign when_Pipeline_l278 = (|pipeline_rsp_haltRequest_Ram_l73);
  always @(*) begin
    pipeline_cmd_ready_output = pipeline_rsp_ready;
    if(when_Connection_l74) begin
      pipeline_cmd_ready_output = 1'b1;
    end
  end

  assign when_Connection_l74 = (! pipeline_rsp_valid);
  assign io_up_a_tracker_last = ((! ((1'b0 || (A_PUT_FULL_DATA == io_up_a_payload_opcode)) || (A_PUT_PARTIAL_DATA == io_up_a_payload_opcode))) || (io_up_a_tracker_beat == _zz_io_up_a_tracker_last));
  assign ordering_valid = (io_up_a_fire && io_up_a_tracker_last);
  assign ordering_payload_bytes = _zz_ordering_payload_bytes[6:0];
  assign mem_en = (port_enable && 1'b1);
  always @(posedge clk_cpu or posedge reset_cpu) begin
    if(reset_cpu) begin
      pipeline_cmd_fsm_counter <= 4'b0000;
      pipeline_rsp_valid <= 1'b0;
      io_up_a_tracker_beat <= 4'b0000;
      ordering_regNext_valid <= 1'b0;
    end else begin
      if(pipeline_cmd_isFireing) begin
        pipeline_cmd_fsm_counter <= (pipeline_cmd_fsm_counter + 4'b0001);
        if(pipeline_cmd_LAST) begin
          pipeline_cmd_fsm_counter <= 4'b0000;
        end
      end
      if(pipeline_cmd_ready_output) begin
        pipeline_rsp_valid <= pipeline_cmd_valid;
      end
      if(io_up_a_fire) begin
        io_up_a_tracker_beat <= (io_up_a_tracker_beat + 4'b0001);
        if(io_up_a_tracker_last) begin
          io_up_a_tracker_beat <= 4'b0000;
        end
      end
      ordering_regNext_valid <= ordering_valid;
    end
  end

  always @(posedge clk_cpu) begin
    if(when_Ram_l47) begin
      pipeline_cmd_fsm_size <= io_up_a_payload_size;
      pipeline_cmd_fsm_source <= io_up_a_payload_source;
      pipeline_cmd_fsm_isGet <= (|(io_up_a_payload_opcode == A_GET));
      pipeline_cmd_fsm_address <= pipeline_cmd_addressShifted;
    end
    if(pipeline_cmd_ready_output) begin
      pipeline_rsp_cmd_IS_GET <= pipeline_cmd_IS_GET;
      pipeline_rsp_cmd_SIZE <= pipeline_cmd_SIZE;
      pipeline_rsp_cmd_SOURCE <= pipeline_cmd_SOURCE;
      pipeline_rsp_cmd_LAST <= pipeline_cmd_LAST;
    end
    ordering_regNext_payload_bytes <= ordering_payload_bytes;
  end


endmodule

module Apb3Bridge (
  input  wire          io_up_a_valid,
  output wire          io_up_a_ready,
  input  wire [2:0]    io_up_a_payload_opcode,
  input  wire [2:0]    io_up_a_payload_param,
  input  wire [2:0]    io_up_a_payload_source,
  input  wire [26:0]   io_up_a_payload_address,
  input  wire [2:0]    io_up_a_payload_size,
  input  wire [3:0]    io_up_a_payload_mask,
  input  wire [31:0]   io_up_a_payload_data,
  input  wire          io_up_a_payload_corrupt,
  output wire          io_up_d_valid,
  input  wire          io_up_d_ready,
  output wire [2:0]    io_up_d_payload_opcode,
  output wire [2:0]    io_up_d_payload_param,
  output wire [2:0]    io_up_d_payload_source,
  output wire [2:0]    io_up_d_payload_size,
  output wire          io_up_d_payload_denied,
  output wire [31:0]   io_up_d_payload_data,
  output wire          io_up_d_payload_corrupt,
  output wire [26:0]   io_down_PADDR,
  output reg  [0:0]    io_down_PSEL,
  output wire          io_down_PENABLE,
  input  wire          io_down_PREADY,
  output wire          io_down_PWRITE,
  output wire [31:0]   io_down_PWDATA,
  input  wire [31:0]   io_down_PRDATA,
  input  wire          io_down_PSLVERROR,
  input  wire          clk_cpu,
  input  wire          reset_cpu
);
  localparam A_PUT_FULL_DATA = 3'd0;
  localparam A_PUT_PARTIAL_DATA = 3'd1;
  localparam A_GET = 3'd4;
  localparam A_ACQUIRE_BLOCK = 3'd6;
  localparam A_ACQUIRE_PERM = 3'd7;
  localparam D_ACCESS_ACK = 3'd0;
  localparam D_ACCESS_ACK_DATA = 3'd1;
  localparam D_GRANT = 3'd4;
  localparam D_GRANT_DATA = 3'd5;
  localparam D_RELEASE_ACK = 3'd6;

  reg        [3:0]    _zz_buffered_ready;
  wire       [26:0]   _zz_io_down_PADDR;
  wire       [5:0]    _zz_io_down_PADDR_1;
  wire                buffered_valid;
  wire                buffered_ready;
  wire       [2:0]    buffered_payload_opcode;
  wire       [2:0]    buffered_payload_param;
  wire       [2:0]    buffered_payload_source;
  wire       [26:0]   buffered_payload_address;
  wire       [2:0]    buffered_payload_size;
  wire       [3:0]    buffered_payload_mask;
  wire       [31:0]   buffered_payload_data;
  wire                buffered_payload_corrupt;
  reg                 io_up_a_rValid;
  wire                buffered_fire;
  reg        [2:0]    io_up_a_rData_opcode;
  reg        [2:0]    io_up_a_rData_param;
  reg        [2:0]    io_up_a_rData_source;
  reg        [26:0]   io_up_a_rData_address;
  reg        [2:0]    io_up_a_rData_size;
  reg        [3:0]    io_up_a_rData_mask;
  reg        [31:0]   io_up_a_rData_data;
  reg                 io_up_a_rData_corrupt;
  wire                isGet;
  reg        [3:0]    counter;
  wire                forked_valid;
  wire                forked_ready;
  wire       [2:0]    forked_payload_opcode;
  wire       [2:0]    forked_payload_param;
  wire       [2:0]    forked_payload_source;
  wire       [26:0]   forked_payload_address;
  wire       [2:0]    forked_payload_size;
  wire       [3:0]    forked_payload_mask;
  wire       [31:0]   forked_payload_data;
  wire                forked_payload_corrupt;
  wire                forked_fire;
  reg                 enable;
  wire                rsp_valid;
  wire                rsp_ready;
  wire       [2:0]    rsp_payload_opcode;
  wire       [2:0]    rsp_payload_param;
  wire       [2:0]    rsp_payload_source;
  wire       [2:0]    rsp_payload_size;
  wire                rsp_payload_denied;
  wire       [31:0]   rsp_payload_data;
  wire                rsp_payload_corrupt;
  wire       [2:0]    _zz_rsp_payload_opcode;
  wire                rsp_halfPipe_valid;
  wire                rsp_halfPipe_ready;
  wire       [2:0]    rsp_halfPipe_payload_opcode;
  wire       [2:0]    rsp_halfPipe_payload_param;
  wire       [2:0]    rsp_halfPipe_payload_source;
  wire       [2:0]    rsp_halfPipe_payload_size;
  wire                rsp_halfPipe_payload_denied;
  wire       [31:0]   rsp_halfPipe_payload_data;
  wire                rsp_halfPipe_payload_corrupt;
  reg                 rsp_rValid;
  wire                rsp_halfPipe_fire;
  reg        [2:0]    rsp_rData_opcode;
  reg        [2:0]    rsp_rData_param;
  reg        [2:0]    rsp_rData_source;
  reg        [2:0]    rsp_rData_size;
  reg                 rsp_rData_denied;
  reg        [31:0]   rsp_rData_data;
  reg                 rsp_rData_corrupt;
  `ifndef SYNTHESIS
  reg [127:0] io_up_a_payload_opcode_string;
  reg [119:0] io_up_d_payload_opcode_string;
  reg [127:0] buffered_payload_opcode_string;
  reg [127:0] io_up_a_rData_opcode_string;
  reg [127:0] forked_payload_opcode_string;
  reg [119:0] rsp_payload_opcode_string;
  reg [119:0] _zz_rsp_payload_opcode_string;
  reg [119:0] rsp_halfPipe_payload_opcode_string;
  reg [119:0] rsp_rData_opcode_string;
  `endif


  assign _zz_io_down_PADDR_1 = ({2'd0,counter} <<< 2'd2);
  assign _zz_io_down_PADDR = {21'd0, _zz_io_down_PADDR_1};
  always @(*) begin
    case(buffered_payload_size)
      3'b000 : _zz_buffered_ready = 4'b0000;
      3'b001 : _zz_buffered_ready = 4'b0000;
      3'b010 : _zz_buffered_ready = 4'b0000;
      3'b011 : _zz_buffered_ready = 4'b0001;
      3'b100 : _zz_buffered_ready = 4'b0011;
      3'b101 : _zz_buffered_ready = 4'b0111;
      default : _zz_buffered_ready = 4'b1111;
    endcase
  end

  `ifndef SYNTHESIS
  always @(*) begin
    case(io_up_a_payload_opcode)
      A_PUT_FULL_DATA : io_up_a_payload_opcode_string = "PUT_FULL_DATA   ";
      A_PUT_PARTIAL_DATA : io_up_a_payload_opcode_string = "PUT_PARTIAL_DATA";
      A_GET : io_up_a_payload_opcode_string = "GET             ";
      A_ACQUIRE_BLOCK : io_up_a_payload_opcode_string = "ACQUIRE_BLOCK   ";
      A_ACQUIRE_PERM : io_up_a_payload_opcode_string = "ACQUIRE_PERM    ";
      default : io_up_a_payload_opcode_string = "????????????????";
    endcase
  end
  always @(*) begin
    case(io_up_d_payload_opcode)
      D_ACCESS_ACK : io_up_d_payload_opcode_string = "ACCESS_ACK     ";
      D_ACCESS_ACK_DATA : io_up_d_payload_opcode_string = "ACCESS_ACK_DATA";
      D_GRANT : io_up_d_payload_opcode_string = "GRANT          ";
      D_GRANT_DATA : io_up_d_payload_opcode_string = "GRANT_DATA     ";
      D_RELEASE_ACK : io_up_d_payload_opcode_string = "RELEASE_ACK    ";
      default : io_up_d_payload_opcode_string = "???????????????";
    endcase
  end
  always @(*) begin
    case(buffered_payload_opcode)
      A_PUT_FULL_DATA : buffered_payload_opcode_string = "PUT_FULL_DATA   ";
      A_PUT_PARTIAL_DATA : buffered_payload_opcode_string = "PUT_PARTIAL_DATA";
      A_GET : buffered_payload_opcode_string = "GET             ";
      A_ACQUIRE_BLOCK : buffered_payload_opcode_string = "ACQUIRE_BLOCK   ";
      A_ACQUIRE_PERM : buffered_payload_opcode_string = "ACQUIRE_PERM    ";
      default : buffered_payload_opcode_string = "????????????????";
    endcase
  end
  always @(*) begin
    case(io_up_a_rData_opcode)
      A_PUT_FULL_DATA : io_up_a_rData_opcode_string = "PUT_FULL_DATA   ";
      A_PUT_PARTIAL_DATA : io_up_a_rData_opcode_string = "PUT_PARTIAL_DATA";
      A_GET : io_up_a_rData_opcode_string = "GET             ";
      A_ACQUIRE_BLOCK : io_up_a_rData_opcode_string = "ACQUIRE_BLOCK   ";
      A_ACQUIRE_PERM : io_up_a_rData_opcode_string = "ACQUIRE_PERM    ";
      default : io_up_a_rData_opcode_string = "????????????????";
    endcase
  end
  always @(*) begin
    case(forked_payload_opcode)
      A_PUT_FULL_DATA : forked_payload_opcode_string = "PUT_FULL_DATA   ";
      A_PUT_PARTIAL_DATA : forked_payload_opcode_string = "PUT_PARTIAL_DATA";
      A_GET : forked_payload_opcode_string = "GET             ";
      A_ACQUIRE_BLOCK : forked_payload_opcode_string = "ACQUIRE_BLOCK   ";
      A_ACQUIRE_PERM : forked_payload_opcode_string = "ACQUIRE_PERM    ";
      default : forked_payload_opcode_string = "????????????????";
    endcase
  end
  always @(*) begin
    case(rsp_payload_opcode)
      D_ACCESS_ACK : rsp_payload_opcode_string = "ACCESS_ACK     ";
      D_ACCESS_ACK_DATA : rsp_payload_opcode_string = "ACCESS_ACK_DATA";
      D_GRANT : rsp_payload_opcode_string = "GRANT          ";
      D_GRANT_DATA : rsp_payload_opcode_string = "GRANT_DATA     ";
      D_RELEASE_ACK : rsp_payload_opcode_string = "RELEASE_ACK    ";
      default : rsp_payload_opcode_string = "???????????????";
    endcase
  end
  always @(*) begin
    case(_zz_rsp_payload_opcode)
      D_ACCESS_ACK : _zz_rsp_payload_opcode_string = "ACCESS_ACK     ";
      D_ACCESS_ACK_DATA : _zz_rsp_payload_opcode_string = "ACCESS_ACK_DATA";
      D_GRANT : _zz_rsp_payload_opcode_string = "GRANT          ";
      D_GRANT_DATA : _zz_rsp_payload_opcode_string = "GRANT_DATA     ";
      D_RELEASE_ACK : _zz_rsp_payload_opcode_string = "RELEASE_ACK    ";
      default : _zz_rsp_payload_opcode_string = "???????????????";
    endcase
  end
  always @(*) begin
    case(rsp_halfPipe_payload_opcode)
      D_ACCESS_ACK : rsp_halfPipe_payload_opcode_string = "ACCESS_ACK     ";
      D_ACCESS_ACK_DATA : rsp_halfPipe_payload_opcode_string = "ACCESS_ACK_DATA";
      D_GRANT : rsp_halfPipe_payload_opcode_string = "GRANT          ";
      D_GRANT_DATA : rsp_halfPipe_payload_opcode_string = "GRANT_DATA     ";
      D_RELEASE_ACK : rsp_halfPipe_payload_opcode_string = "RELEASE_ACK    ";
      default : rsp_halfPipe_payload_opcode_string = "???????????????";
    endcase
  end
  always @(*) begin
    case(rsp_rData_opcode)
      D_ACCESS_ACK : rsp_rData_opcode_string = "ACCESS_ACK     ";
      D_ACCESS_ACK_DATA : rsp_rData_opcode_string = "ACCESS_ACK_DATA";
      D_GRANT : rsp_rData_opcode_string = "GRANT          ";
      D_GRANT_DATA : rsp_rData_opcode_string = "GRANT_DATA     ";
      D_RELEASE_ACK : rsp_rData_opcode_string = "RELEASE_ACK    ";
      default : rsp_rData_opcode_string = "???????????????";
    endcase
  end
  `endif

  assign buffered_fire = (buffered_valid && buffered_ready);
  assign io_up_a_ready = (! io_up_a_rValid);
  assign buffered_valid = io_up_a_rValid;
  assign buffered_payload_opcode = io_up_a_rData_opcode;
  assign buffered_payload_param = io_up_a_rData_param;
  assign buffered_payload_source = io_up_a_rData_source;
  assign buffered_payload_address = io_up_a_rData_address;
  assign buffered_payload_size = io_up_a_rData_size;
  assign buffered_payload_mask = io_up_a_rData_mask;
  assign buffered_payload_data = io_up_a_rData_data;
  assign buffered_payload_corrupt = io_up_a_rData_corrupt;
  assign isGet = (buffered_payload_opcode == A_GET);
  assign forked_valid = buffered_valid;
  assign forked_payload_opcode = buffered_payload_opcode;
  assign forked_payload_param = buffered_payload_param;
  assign forked_payload_source = buffered_payload_source;
  assign forked_payload_address = buffered_payload_address;
  assign forked_payload_size = buffered_payload_size;
  assign forked_payload_mask = buffered_payload_mask;
  assign forked_payload_data = buffered_payload_data;
  assign forked_payload_corrupt = buffered_payload_corrupt;
  assign buffered_ready = (forked_ready && ((! isGet) || (counter == _zz_buffered_ready)));
  assign forked_fire = (forked_valid && forked_ready);
  assign forked_ready = (enable && io_down_PREADY);
  always @(*) begin
    io_down_PSEL[0] = buffered_valid;
    if(io_up_d_valid) begin
      io_down_PSEL[0] = 1'b0;
    end
  end

  assign io_down_PENABLE = enable;
  assign io_down_PADDR = (buffered_payload_address | _zz_io_down_PADDR);
  assign io_down_PWRITE = (! isGet);
  assign io_down_PWDATA = buffered_payload_data;
  assign rsp_valid = forked_fire;
  assign _zz_rsp_payload_opcode = (isGet ? D_ACCESS_ACK_DATA : D_ACCESS_ACK);
  assign rsp_payload_opcode = _zz_rsp_payload_opcode;
  assign rsp_payload_param = 3'b000;
  assign rsp_payload_source = buffered_payload_source;
  assign rsp_payload_size = buffered_payload_size;
  assign rsp_payload_data = io_down_PRDATA;
  assign rsp_payload_denied = io_down_PSLVERROR;
  assign rsp_payload_corrupt = 1'b0;
  assign rsp_halfPipe_fire = (rsp_halfPipe_valid && rsp_halfPipe_ready);
  assign rsp_ready = (! rsp_rValid);
  assign rsp_halfPipe_valid = rsp_rValid;
  assign rsp_halfPipe_payload_opcode = rsp_rData_opcode;
  assign rsp_halfPipe_payload_param = rsp_rData_param;
  assign rsp_halfPipe_payload_source = rsp_rData_source;
  assign rsp_halfPipe_payload_size = rsp_rData_size;
  assign rsp_halfPipe_payload_denied = rsp_rData_denied;
  assign rsp_halfPipe_payload_data = rsp_rData_data;
  assign rsp_halfPipe_payload_corrupt = rsp_rData_corrupt;
  assign io_up_d_valid = rsp_halfPipe_valid;
  assign rsp_halfPipe_ready = io_up_d_ready;
  assign io_up_d_payload_opcode = rsp_halfPipe_payload_opcode;
  assign io_up_d_payload_param = rsp_halfPipe_payload_param;
  assign io_up_d_payload_source = rsp_halfPipe_payload_source;
  assign io_up_d_payload_size = rsp_halfPipe_payload_size;
  assign io_up_d_payload_denied = rsp_halfPipe_payload_denied;
  assign io_up_d_payload_data = rsp_halfPipe_payload_data;
  assign io_up_d_payload_corrupt = rsp_halfPipe_payload_corrupt;
  always @(posedge clk_cpu or posedge reset_cpu) begin
    if(reset_cpu) begin
      io_up_a_rValid <= 1'b0;
      counter <= 4'b0000;
      enable <= 1'b0;
      rsp_rValid <= 1'b0;
    end else begin
      if(io_up_a_valid) begin
        io_up_a_rValid <= 1'b1;
      end
      if(buffered_fire) begin
        io_up_a_rValid <= 1'b0;
      end
      if(forked_fire) begin
        counter <= (counter + 4'b0001);
        if(buffered_fire) begin
          counter <= 4'b0000;
        end
      end
      enable <= (enable ? (! io_down_PREADY) : io_down_PSEL[0]);
      if(rsp_valid) begin
        rsp_rValid <= 1'b1;
      end
      if(rsp_halfPipe_fire) begin
        rsp_rValid <= 1'b0;
      end
    end
  end

  always @(posedge clk_cpu) begin
    if(io_up_a_ready) begin
      io_up_a_rData_opcode <= io_up_a_payload_opcode;
      io_up_a_rData_param <= io_up_a_payload_param;
      io_up_a_rData_source <= io_up_a_payload_source;
      io_up_a_rData_address <= io_up_a_payload_address;
      io_up_a_rData_size <= io_up_a_payload_size;
      io_up_a_rData_mask <= io_up_a_payload_mask;
      io_up_a_rData_data <= io_up_a_payload_data;
      io_up_a_rData_corrupt <= io_up_a_payload_corrupt;
    end
    if(rsp_ready) begin
      rsp_rData_opcode <= rsp_payload_opcode;
      rsp_rData_param <= rsp_payload_param;
      rsp_rData_source <= rsp_payload_source;
      rsp_rData_size <= rsp_payload_size;
      rsp_rData_denied <= rsp_payload_denied;
      rsp_rData_data <= rsp_payload_data;
      rsp_rData_corrupt <= rsp_payload_corrupt;
    end
  end


endmodule

module Decoder (
  input  wire          io_up_a_valid,
  output wire          io_up_a_ready,
  input  wire [2:0]    io_up_a_payload_opcode,
  input  wire [2:0]    io_up_a_payload_param,
  input  wire [2:0]    io_up_a_payload_source,
  input  wire [31:0]   io_up_a_payload_address,
  input  wire [2:0]    io_up_a_payload_size,
  input  wire [7:0]    io_up_a_payload_mask,
  input  wire [63:0]   io_up_a_payload_data,
  input  wire          io_up_a_payload_corrupt,
  output wire          io_up_d_valid,
  input  wire          io_up_d_ready,
  output wire [2:0]    io_up_d_payload_opcode,
  output wire [2:0]    io_up_d_payload_param,
  output wire [2:0]    io_up_d_payload_source,
  output wire [2:0]    io_up_d_payload_size,
  output wire          io_up_d_payload_denied,
  output wire [63:0]   io_up_d_payload_data,
  output wire          io_up_d_payload_corrupt,
  output wire          io_downs_0_a_valid,
  input  wire          io_downs_0_a_ready,
  output wire [2:0]    io_downs_0_a_payload_opcode,
  output wire [2:0]    io_downs_0_a_payload_param,
  output wire [2:0]    io_downs_0_a_payload_source,
  output wire [30:0]   io_downs_0_a_payload_address,
  output wire [2:0]    io_downs_0_a_payload_size,
  output wire [7:0]    io_downs_0_a_payload_mask,
  output wire [63:0]   io_downs_0_a_payload_data,
  output wire          io_downs_0_a_payload_corrupt,
  input  wire          io_downs_0_d_valid,
  output wire          io_downs_0_d_ready,
  input  wire [2:0]    io_downs_0_d_payload_opcode,
  input  wire [2:0]    io_downs_0_d_payload_param,
  input  wire [2:0]    io_downs_0_d_payload_source,
  input  wire [2:0]    io_downs_0_d_payload_size,
  input  wire          io_downs_0_d_payload_denied,
  input  wire [63:0]   io_downs_0_d_payload_data,
  input  wire          io_downs_0_d_payload_corrupt,
  output wire          io_downs_1_a_valid,
  input  wire          io_downs_1_a_ready,
  output wire [2:0]    io_downs_1_a_payload_opcode,
  output wire [2:0]    io_downs_1_a_payload_param,
  output wire [2:0]    io_downs_1_a_payload_source,
  output wire [26:0]   io_downs_1_a_payload_address,
  output wire [2:0]    io_downs_1_a_payload_size,
  output wire [7:0]    io_downs_1_a_payload_mask,
  output wire [63:0]   io_downs_1_a_payload_data,
  output wire          io_downs_1_a_payload_corrupt,
  input  wire          io_downs_1_d_valid,
  output wire          io_downs_1_d_ready,
  input  wire [2:0]    io_downs_1_d_payload_opcode,
  input  wire [2:0]    io_downs_1_d_payload_param,
  input  wire [2:0]    io_downs_1_d_payload_source,
  input  wire [2:0]    io_downs_1_d_payload_size,
  input  wire          io_downs_1_d_payload_denied,
  input  wire [63:0]   io_downs_1_d_payload_data,
  input  wire          io_downs_1_d_payload_corrupt,
  input  wire          clk_cpu,
  input  wire          reset_cpu
);
  localparam A_PUT_FULL_DATA = 3'd0;
  localparam A_PUT_PARTIAL_DATA = 3'd1;
  localparam A_GET = 3'd4;
  localparam A_ACQUIRE_BLOCK = 3'd6;
  localparam A_ACQUIRE_PERM = 3'd7;
  localparam D_ACCESS_ACK = 3'd0;
  localparam D_ACCESS_ACK_DATA = 3'd1;
  localparam D_GRANT = 3'd4;
  localparam D_GRANT_DATA = 3'd5;
  localparam D_RELEASE_ACK = 3'd6;

  wire                d_arbiter_io_inputs_0_ready;
  wire                d_arbiter_io_inputs_1_ready;
  wire                d_arbiter_io_output_valid;
  wire       [2:0]    d_arbiter_io_output_payload_opcode;
  wire       [2:0]    d_arbiter_io_output_payload_param;
  wire       [2:0]    d_arbiter_io_output_payload_source;
  wire       [2:0]    d_arbiter_io_output_payload_size;
  wire                d_arbiter_io_output_payload_denied;
  wire       [63:0]   d_arbiter_io_output_payload_data;
  wire                d_arbiter_io_output_payload_corrupt;
  wire       [0:0]    d_arbiter_io_chosen;
  wire       [1:0]    d_arbiter_io_chosenOH;
  wire       [0:0]    _zz_a_logic_0_hit;
  wire       [0:0]    _zz_a_logic_1_hit;
  wire       [31:0]   _zz_downs_1_a_payload_address;
  reg        [1:0]    _zz_1;
  wire       [1:0]    _zz_2;
  wire                downs_0_a_valid;
  wire                downs_0_a_ready;
  wire       [2:0]    downs_0_a_payload_opcode;
  wire       [2:0]    downs_0_a_payload_param;
  wire       [2:0]    downs_0_a_payload_source;
  wire       [30:0]   downs_0_a_payload_address;
  wire       [2:0]    downs_0_a_payload_size;
  wire       [7:0]    downs_0_a_payload_mask;
  wire       [63:0]   downs_0_a_payload_data;
  wire                downs_0_a_payload_corrupt;
  wire                downs_0_d_valid;
  wire                downs_0_d_ready;
  wire       [2:0]    downs_0_d_payload_opcode;
  wire       [2:0]    downs_0_d_payload_param;
  wire       [2:0]    downs_0_d_payload_source;
  wire       [2:0]    downs_0_d_payload_size;
  wire                downs_0_d_payload_denied;
  wire       [63:0]   downs_0_d_payload_data;
  wire                downs_0_d_payload_corrupt;
  wire                downs_1_a_valid;
  wire                downs_1_a_ready;
  wire       [2:0]    downs_1_a_payload_opcode;
  wire       [2:0]    downs_1_a_payload_param;
  wire       [2:0]    downs_1_a_payload_source;
  wire       [26:0]   downs_1_a_payload_address;
  wire       [2:0]    downs_1_a_payload_size;
  wire       [7:0]    downs_1_a_payload_mask;
  wire       [63:0]   downs_1_a_payload_data;
  wire                downs_1_a_payload_corrupt;
  wire                downs_1_d_valid;
  wire                downs_1_d_ready;
  wire       [2:0]    downs_1_d_payload_opcode;
  wire       [2:0]    downs_1_d_payload_param;
  wire       [2:0]    downs_1_d_payload_source;
  wire       [2:0]    downs_1_d_payload_size;
  wire                downs_1_d_payload_denied;
  wire       [63:0]   downs_1_d_payload_data;
  wire                downs_1_d_payload_corrupt;
  wire       [34:0]   a_key;
  wire                a_logic_0_hit;
  wire                a_logic_1_hit;
  wire                a_miss;
  `ifndef SYNTHESIS
  reg [127:0] io_up_a_payload_opcode_string;
  reg [119:0] io_up_d_payload_opcode_string;
  reg [127:0] io_downs_0_a_payload_opcode_string;
  reg [119:0] io_downs_0_d_payload_opcode_string;
  reg [127:0] io_downs_1_a_payload_opcode_string;
  reg [119:0] io_downs_1_d_payload_opcode_string;
  reg [127:0] downs_0_a_payload_opcode_string;
  reg [119:0] downs_0_d_payload_opcode_string;
  reg [127:0] downs_1_a_payload_opcode_string;
  reg [119:0] downs_1_d_payload_opcode_string;
  `endif


  assign _zz_a_logic_0_hit = (|((a_key & 35'h080000000) == 35'h0));
  assign _zz_a_logic_1_hit = (|((a_key & 35'h080000000) == 35'h080000000));
  assign _zz_downs_1_a_payload_address = (io_up_a_payload_address - 32'h80000000);
  assign _zz_2 = {io_downs_1_a_valid,io_downs_0_a_valid};
  StreamArbiter_7 d_arbiter (
    .io_inputs_0_valid           (downs_0_d_valid                        ), //i
    .io_inputs_0_ready           (d_arbiter_io_inputs_0_ready            ), //o
    .io_inputs_0_payload_opcode  (downs_0_d_payload_opcode[2:0]          ), //i
    .io_inputs_0_payload_param   (downs_0_d_payload_param[2:0]           ), //i
    .io_inputs_0_payload_source  (downs_0_d_payload_source[2:0]          ), //i
    .io_inputs_0_payload_size    (downs_0_d_payload_size[2:0]            ), //i
    .io_inputs_0_payload_denied  (downs_0_d_payload_denied               ), //i
    .io_inputs_0_payload_data    (downs_0_d_payload_data[63:0]           ), //i
    .io_inputs_0_payload_corrupt (downs_0_d_payload_corrupt              ), //i
    .io_inputs_1_valid           (downs_1_d_valid                        ), //i
    .io_inputs_1_ready           (d_arbiter_io_inputs_1_ready            ), //o
    .io_inputs_1_payload_opcode  (downs_1_d_payload_opcode[2:0]          ), //i
    .io_inputs_1_payload_param   (downs_1_d_payload_param[2:0]           ), //i
    .io_inputs_1_payload_source  (downs_1_d_payload_source[2:0]          ), //i
    .io_inputs_1_payload_size    (downs_1_d_payload_size[2:0]            ), //i
    .io_inputs_1_payload_denied  (downs_1_d_payload_denied               ), //i
    .io_inputs_1_payload_data    (downs_1_d_payload_data[63:0]           ), //i
    .io_inputs_1_payload_corrupt (downs_1_d_payload_corrupt              ), //i
    .io_output_valid             (d_arbiter_io_output_valid              ), //o
    .io_output_ready             (io_up_d_ready                          ), //i
    .io_output_payload_opcode    (d_arbiter_io_output_payload_opcode[2:0]), //o
    .io_output_payload_param     (d_arbiter_io_output_payload_param[2:0] ), //o
    .io_output_payload_source    (d_arbiter_io_output_payload_source[2:0]), //o
    .io_output_payload_size      (d_arbiter_io_output_payload_size[2:0]  ), //o
    .io_output_payload_denied    (d_arbiter_io_output_payload_denied     ), //o
    .io_output_payload_data      (d_arbiter_io_output_payload_data[63:0] ), //o
    .io_output_payload_corrupt   (d_arbiter_io_output_payload_corrupt    ), //o
    .io_chosen                   (d_arbiter_io_chosen                    ), //o
    .io_chosenOH                 (d_arbiter_io_chosenOH[1:0]             ), //o
    .clk_cpu                     (clk_cpu                                ), //i
    .reset_cpu                   (reset_cpu                              )  //i
  );
  always @(*) begin
    case(_zz_2)
      2'b00 : _zz_1 = 2'b00;
      2'b01 : _zz_1 = 2'b01;
      2'b10 : _zz_1 = 2'b01;
      default : _zz_1 = 2'b10;
    endcase
  end

  `ifndef SYNTHESIS
  always @(*) begin
    case(io_up_a_payload_opcode)
      A_PUT_FULL_DATA : io_up_a_payload_opcode_string = "PUT_FULL_DATA   ";
      A_PUT_PARTIAL_DATA : io_up_a_payload_opcode_string = "PUT_PARTIAL_DATA";
      A_GET : io_up_a_payload_opcode_string = "GET             ";
      A_ACQUIRE_BLOCK : io_up_a_payload_opcode_string = "ACQUIRE_BLOCK   ";
      A_ACQUIRE_PERM : io_up_a_payload_opcode_string = "ACQUIRE_PERM    ";
      default : io_up_a_payload_opcode_string = "????????????????";
    endcase
  end
  always @(*) begin
    case(io_up_d_payload_opcode)
      D_ACCESS_ACK : io_up_d_payload_opcode_string = "ACCESS_ACK     ";
      D_ACCESS_ACK_DATA : io_up_d_payload_opcode_string = "ACCESS_ACK_DATA";
      D_GRANT : io_up_d_payload_opcode_string = "GRANT          ";
      D_GRANT_DATA : io_up_d_payload_opcode_string = "GRANT_DATA     ";
      D_RELEASE_ACK : io_up_d_payload_opcode_string = "RELEASE_ACK    ";
      default : io_up_d_payload_opcode_string = "???????????????";
    endcase
  end
  always @(*) begin
    case(io_downs_0_a_payload_opcode)
      A_PUT_FULL_DATA : io_downs_0_a_payload_opcode_string = "PUT_FULL_DATA   ";
      A_PUT_PARTIAL_DATA : io_downs_0_a_payload_opcode_string = "PUT_PARTIAL_DATA";
      A_GET : io_downs_0_a_payload_opcode_string = "GET             ";
      A_ACQUIRE_BLOCK : io_downs_0_a_payload_opcode_string = "ACQUIRE_BLOCK   ";
      A_ACQUIRE_PERM : io_downs_0_a_payload_opcode_string = "ACQUIRE_PERM    ";
      default : io_downs_0_a_payload_opcode_string = "????????????????";
    endcase
  end
  always @(*) begin
    case(io_downs_0_d_payload_opcode)
      D_ACCESS_ACK : io_downs_0_d_payload_opcode_string = "ACCESS_ACK     ";
      D_ACCESS_ACK_DATA : io_downs_0_d_payload_opcode_string = "ACCESS_ACK_DATA";
      D_GRANT : io_downs_0_d_payload_opcode_string = "GRANT          ";
      D_GRANT_DATA : io_downs_0_d_payload_opcode_string = "GRANT_DATA     ";
      D_RELEASE_ACK : io_downs_0_d_payload_opcode_string = "RELEASE_ACK    ";
      default : io_downs_0_d_payload_opcode_string = "???????????????";
    endcase
  end
  always @(*) begin
    case(io_downs_1_a_payload_opcode)
      A_PUT_FULL_DATA : io_downs_1_a_payload_opcode_string = "PUT_FULL_DATA   ";
      A_PUT_PARTIAL_DATA : io_downs_1_a_payload_opcode_string = "PUT_PARTIAL_DATA";
      A_GET : io_downs_1_a_payload_opcode_string = "GET             ";
      A_ACQUIRE_BLOCK : io_downs_1_a_payload_opcode_string = "ACQUIRE_BLOCK   ";
      A_ACQUIRE_PERM : io_downs_1_a_payload_opcode_string = "ACQUIRE_PERM    ";
      default : io_downs_1_a_payload_opcode_string = "????????????????";
    endcase
  end
  always @(*) begin
    case(io_downs_1_d_payload_opcode)
      D_ACCESS_ACK : io_downs_1_d_payload_opcode_string = "ACCESS_ACK     ";
      D_ACCESS_ACK_DATA : io_downs_1_d_payload_opcode_string = "ACCESS_ACK_DATA";
      D_GRANT : io_downs_1_d_payload_opcode_string = "GRANT          ";
      D_GRANT_DATA : io_downs_1_d_payload_opcode_string = "GRANT_DATA     ";
      D_RELEASE_ACK : io_downs_1_d_payload_opcode_string = "RELEASE_ACK    ";
      default : io_downs_1_d_payload_opcode_string = "???????????????";
    endcase
  end
  always @(*) begin
    case(downs_0_a_payload_opcode)
      A_PUT_FULL_DATA : downs_0_a_payload_opcode_string = "PUT_FULL_DATA   ";
      A_PUT_PARTIAL_DATA : downs_0_a_payload_opcode_string = "PUT_PARTIAL_DATA";
      A_GET : downs_0_a_payload_opcode_string = "GET             ";
      A_ACQUIRE_BLOCK : downs_0_a_payload_opcode_string = "ACQUIRE_BLOCK   ";
      A_ACQUIRE_PERM : downs_0_a_payload_opcode_string = "ACQUIRE_PERM    ";
      default : downs_0_a_payload_opcode_string = "????????????????";
    endcase
  end
  always @(*) begin
    case(downs_0_d_payload_opcode)
      D_ACCESS_ACK : downs_0_d_payload_opcode_string = "ACCESS_ACK     ";
      D_ACCESS_ACK_DATA : downs_0_d_payload_opcode_string = "ACCESS_ACK_DATA";
      D_GRANT : downs_0_d_payload_opcode_string = "GRANT          ";
      D_GRANT_DATA : downs_0_d_payload_opcode_string = "GRANT_DATA     ";
      D_RELEASE_ACK : downs_0_d_payload_opcode_string = "RELEASE_ACK    ";
      default : downs_0_d_payload_opcode_string = "???????????????";
    endcase
  end
  always @(*) begin
    case(downs_1_a_payload_opcode)
      A_PUT_FULL_DATA : downs_1_a_payload_opcode_string = "PUT_FULL_DATA   ";
      A_PUT_PARTIAL_DATA : downs_1_a_payload_opcode_string = "PUT_PARTIAL_DATA";
      A_GET : downs_1_a_payload_opcode_string = "GET             ";
      A_ACQUIRE_BLOCK : downs_1_a_payload_opcode_string = "ACQUIRE_BLOCK   ";
      A_ACQUIRE_PERM : downs_1_a_payload_opcode_string = "ACQUIRE_PERM    ";
      default : downs_1_a_payload_opcode_string = "????????????????";
    endcase
  end
  always @(*) begin
    case(downs_1_d_payload_opcode)
      D_ACCESS_ACK : downs_1_d_payload_opcode_string = "ACCESS_ACK     ";
      D_ACCESS_ACK_DATA : downs_1_d_payload_opcode_string = "ACCESS_ACK_DATA";
      D_GRANT : downs_1_d_payload_opcode_string = "GRANT          ";
      D_GRANT_DATA : downs_1_d_payload_opcode_string = "GRANT_DATA     ";
      D_RELEASE_ACK : downs_1_d_payload_opcode_string = "RELEASE_ACK    ";
      default : downs_1_d_payload_opcode_string = "???????????????";
    endcase
  end
  `endif

  assign io_downs_0_a_valid = downs_0_a_valid;
  assign downs_0_a_ready = io_downs_0_a_ready;
  assign io_downs_0_a_payload_opcode = downs_0_a_payload_opcode;
  assign io_downs_0_a_payload_param = downs_0_a_payload_param;
  assign io_downs_0_a_payload_source = downs_0_a_payload_source;
  assign io_downs_0_a_payload_address = downs_0_a_payload_address;
  assign io_downs_0_a_payload_size = downs_0_a_payload_size;
  assign io_downs_0_a_payload_mask = downs_0_a_payload_mask;
  assign io_downs_0_a_payload_data = downs_0_a_payload_data;
  assign io_downs_0_a_payload_corrupt = downs_0_a_payload_corrupt;
  assign downs_0_d_valid = io_downs_0_d_valid;
  assign io_downs_0_d_ready = downs_0_d_ready;
  assign downs_0_d_payload_opcode = io_downs_0_d_payload_opcode;
  assign downs_0_d_payload_param = io_downs_0_d_payload_param;
  assign downs_0_d_payload_source = io_downs_0_d_payload_source;
  assign downs_0_d_payload_size = io_downs_0_d_payload_size;
  assign downs_0_d_payload_denied = io_downs_0_d_payload_denied;
  assign downs_0_d_payload_data = io_downs_0_d_payload_data;
  assign downs_0_d_payload_corrupt = io_downs_0_d_payload_corrupt;
  assign io_downs_1_a_valid = downs_1_a_valid;
  assign downs_1_a_ready = io_downs_1_a_ready;
  assign io_downs_1_a_payload_opcode = downs_1_a_payload_opcode;
  assign io_downs_1_a_payload_param = downs_1_a_payload_param;
  assign io_downs_1_a_payload_source = downs_1_a_payload_source;
  assign io_downs_1_a_payload_address = downs_1_a_payload_address;
  assign io_downs_1_a_payload_size = downs_1_a_payload_size;
  assign io_downs_1_a_payload_mask = downs_1_a_payload_mask;
  assign io_downs_1_a_payload_data = downs_1_a_payload_data;
  assign io_downs_1_a_payload_corrupt = downs_1_a_payload_corrupt;
  assign downs_1_d_valid = io_downs_1_d_valid;
  assign io_downs_1_d_ready = downs_1_d_ready;
  assign downs_1_d_payload_opcode = io_downs_1_d_payload_opcode;
  assign downs_1_d_payload_param = io_downs_1_d_payload_param;
  assign downs_1_d_payload_source = io_downs_1_d_payload_source;
  assign downs_1_d_payload_size = io_downs_1_d_payload_size;
  assign downs_1_d_payload_denied = io_downs_1_d_payload_denied;
  assign downs_1_d_payload_data = io_downs_1_d_payload_data;
  assign downs_1_d_payload_corrupt = io_downs_1_d_payload_corrupt;
  assign a_key = {io_up_a_payload_opcode,io_up_a_payload_address};
  assign a_logic_0_hit = _zz_a_logic_0_hit[0];
  assign downs_0_a_valid = (io_up_a_valid && a_logic_0_hit);
  assign downs_0_a_payload_opcode = io_up_a_payload_opcode;
  assign downs_0_a_payload_param = io_up_a_payload_param;
  assign downs_0_a_payload_source = io_up_a_payload_source;
  assign downs_0_a_payload_mask = io_up_a_payload_mask;
  assign downs_0_a_payload_data = io_up_a_payload_data;
  assign downs_0_a_payload_corrupt = io_up_a_payload_corrupt;
  assign downs_0_a_payload_address = io_up_a_payload_address[30:0];
  assign downs_0_a_payload_size = io_up_a_payload_size;
  assign a_logic_1_hit = _zz_a_logic_1_hit[0];
  assign downs_1_a_valid = (io_up_a_valid && a_logic_1_hit);
  assign downs_1_a_payload_opcode = io_up_a_payload_opcode;
  assign downs_1_a_payload_param = io_up_a_payload_param;
  assign downs_1_a_payload_source = io_up_a_payload_source;
  assign downs_1_a_payload_mask = io_up_a_payload_mask;
  assign downs_1_a_payload_data = io_up_a_payload_data;
  assign downs_1_a_payload_corrupt = io_up_a_payload_corrupt;
  assign downs_1_a_payload_address = _zz_downs_1_a_payload_address[26:0];
  assign downs_1_a_payload_size = io_up_a_payload_size;
  assign io_up_a_ready = (|{(downs_1_a_ready && a_logic_1_hit),(downs_0_a_ready && a_logic_0_hit)});
  assign a_miss = (! (|{a_logic_1_hit,a_logic_0_hit}));
  assign downs_0_d_ready = d_arbiter_io_inputs_0_ready;
  assign downs_1_d_ready = d_arbiter_io_inputs_1_ready;
  assign io_up_d_valid = d_arbiter_io_output_valid;
  assign io_up_d_payload_opcode = d_arbiter_io_output_payload_opcode;
  assign io_up_d_payload_param = d_arbiter_io_output_payload_param;
  assign io_up_d_payload_source = d_arbiter_io_output_payload_source;
  assign io_up_d_payload_size = d_arbiter_io_output_payload_size;
  assign io_up_d_payload_denied = d_arbiter_io_output_payload_denied;
  assign io_up_d_payload_data = d_arbiter_io_output_payload_data;
  assign io_up_d_payload_corrupt = d_arbiter_io_output_payload_corrupt;
  always @(posedge clk_cpu or posedge reset_cpu) begin
    if(reset_cpu) begin
    end else begin
      `ifndef SYNTHESIS
        `ifdef FORMAL
          assert((! (io_up_a_valid && a_miss))); // Decoder.scala:L106
        `else
          if(!(! (io_up_a_valid && a_miss))) begin
            $display("FAILURE Tilelink decoder miss ???"); // Decoder.scala:L106
            $finish;
          end
        `endif
      `endif
      `ifndef SYNTHESIS
        `ifdef FORMAL
          assert((! (io_up_a_valid && (_zz_1 != 2'b01)))); // Decoder.scala:L107
        `else
          if(!(! (io_up_a_valid && (_zz_1 != 2'b01)))) begin
            $display("FAILURE Tilelink decoder miss ???"); // Decoder.scala:L107
            $finish;
          end
        `endif
      `endif
    end
  end


endmodule

module Axi4SharedCC (
  input  wire          io_input_arw_valid,
  output wire          io_input_arw_ready,
  input  wire [26:0]   io_input_arw_payload_addr,
  input  wire [2:0]    io_input_arw_payload_id,
  input  wire [7:0]    io_input_arw_payload_len,
  input  wire [2:0]    io_input_arw_payload_size,
  input  wire [1:0]    io_input_arw_payload_burst,
  input  wire          io_input_arw_payload_allStrb,
  input  wire          io_input_arw_payload_write,
  input  wire          io_input_w_valid,
  output wire          io_input_w_ready,
  input  wire [63:0]   io_input_w_payload_data,
  input  wire [7:0]    io_input_w_payload_strb,
  input  wire          io_input_w_payload_last,
  output wire          io_input_b_valid,
  input  wire          io_input_b_ready,
  output wire [2:0]    io_input_b_payload_id,
  output wire [1:0]    io_input_b_payload_resp,
  output wire          io_input_r_valid,
  input  wire          io_input_r_ready,
  output wire [63:0]   io_input_r_payload_data,
  output wire [2:0]    io_input_r_payload_id,
  output wire [1:0]    io_input_r_payload_resp,
  output wire          io_input_r_payload_last,
  output wire          io_output_arw_valid,
  input  wire          io_output_arw_ready,
  output wire [26:0]   io_output_arw_payload_addr,
  output wire [2:0]    io_output_arw_payload_id,
  output wire [7:0]    io_output_arw_payload_len,
  output wire [2:0]    io_output_arw_payload_size,
  output wire [1:0]    io_output_arw_payload_burst,
  output wire          io_output_arw_payload_allStrb,
  output wire          io_output_arw_payload_write,
  output wire          io_output_w_valid,
  input  wire          io_output_w_ready,
  output wire [63:0]   io_output_w_payload_data,
  output wire [7:0]    io_output_w_payload_strb,
  output wire          io_output_w_payload_last,
  input  wire          io_output_b_valid,
  output wire          io_output_b_ready,
  input  wire [2:0]    io_output_b_payload_id,
  input  wire [1:0]    io_output_b_payload_resp,
  input  wire          io_output_r_valid,
  output wire          io_output_r_ready,
  input  wire [63:0]   io_output_r_payload_data,
  input  wire [2:0]    io_output_r_payload_id,
  input  wire [1:0]    io_output_r_payload_resp,
  input  wire          io_output_r_payload_last,
  input  wire          clk_cpu,
  input  wire          reset_cpu,
  input  wire          clk_ram_bus,
  input  wire          reset_ram
);

  wire                io_input_arw_queue_io_push_ready;
  wire                io_input_arw_queue_io_pop_valid;
  wire       [26:0]   io_input_arw_queue_io_pop_payload_addr;
  wire       [2:0]    io_input_arw_queue_io_pop_payload_id;
  wire       [7:0]    io_input_arw_queue_io_pop_payload_len;
  wire       [2:0]    io_input_arw_queue_io_pop_payload_size;
  wire       [1:0]    io_input_arw_queue_io_pop_payload_burst;
  wire                io_input_arw_queue_io_pop_payload_allStrb;
  wire                io_input_arw_queue_io_pop_payload_write;
  wire       [1:0]    io_input_arw_queue_io_pushOccupancy;
  wire       [1:0]    io_input_arw_queue_io_popOccupancy;
  wire                io_input_arw_queue_ram_axi_cc_toplevel_board_ctrl_reset_cpu_synchronized_1;
  wire                io_output_r_queue_io_push_ready;
  wire                io_output_r_queue_io_pop_valid;
  wire       [63:0]   io_output_r_queue_io_pop_payload_data;
  wire       [2:0]    io_output_r_queue_io_pop_payload_id;
  wire       [1:0]    io_output_r_queue_io_pop_payload_resp;
  wire                io_output_r_queue_io_pop_payload_last;
  wire       [7:0]    io_output_r_queue_io_pushOccupancy;
  wire       [7:0]    io_output_r_queue_io_popOccupancy;
  wire                io_output_r_queue_ram_axi_cc_toplevel_board_ctrl_reset_ram_synchronized_1;
  wire                io_input_w_queue_io_push_ready;
  wire                io_input_w_queue_io_pop_valid;
  wire       [63:0]   io_input_w_queue_io_pop_payload_data;
  wire       [7:0]    io_input_w_queue_io_pop_payload_strb;
  wire                io_input_w_queue_io_pop_payload_last;
  wire       [4:0]    io_input_w_queue_io_pushOccupancy;
  wire       [4:0]    io_input_w_queue_io_popOccupancy;
  wire                io_output_b_queue_io_push_ready;
  wire                io_output_b_queue_io_pop_valid;
  wire       [2:0]    io_output_b_queue_io_pop_payload_id;
  wire       [1:0]    io_output_b_queue_io_pop_payload_resp;
  wire       [1:0]    io_output_b_queue_io_pushOccupancy;
  wire       [1:0]    io_output_b_queue_io_popOccupancy;

  StreamFifoCC io_input_arw_queue (
    .io_push_valid                                           (io_input_arw_valid                                                        ), //i
    .io_push_ready                                           (io_input_arw_queue_io_push_ready                                          ), //o
    .io_push_payload_addr                                    (io_input_arw_payload_addr[26:0]                                           ), //i
    .io_push_payload_id                                      (io_input_arw_payload_id[2:0]                                              ), //i
    .io_push_payload_len                                     (io_input_arw_payload_len[7:0]                                             ), //i
    .io_push_payload_size                                    (io_input_arw_payload_size[2:0]                                            ), //i
    .io_push_payload_burst                                   (io_input_arw_payload_burst[1:0]                                           ), //i
    .io_push_payload_allStrb                                 (io_input_arw_payload_allStrb                                              ), //i
    .io_push_payload_write                                   (io_input_arw_payload_write                                                ), //i
    .io_pop_valid                                            (io_input_arw_queue_io_pop_valid                                           ), //o
    .io_pop_ready                                            (io_output_arw_ready                                                       ), //i
    .io_pop_payload_addr                                     (io_input_arw_queue_io_pop_payload_addr[26:0]                              ), //o
    .io_pop_payload_id                                       (io_input_arw_queue_io_pop_payload_id[2:0]                                 ), //o
    .io_pop_payload_len                                      (io_input_arw_queue_io_pop_payload_len[7:0]                                ), //o
    .io_pop_payload_size                                     (io_input_arw_queue_io_pop_payload_size[2:0]                               ), //o
    .io_pop_payload_burst                                    (io_input_arw_queue_io_pop_payload_burst[1:0]                              ), //o
    .io_pop_payload_allStrb                                  (io_input_arw_queue_io_pop_payload_allStrb                                 ), //o
    .io_pop_payload_write                                    (io_input_arw_queue_io_pop_payload_write                                   ), //o
    .io_pushOccupancy                                        (io_input_arw_queue_io_pushOccupancy[1:0]                                  ), //o
    .io_popOccupancy                                         (io_input_arw_queue_io_popOccupancy[1:0]                                   ), //o
    .clk_cpu                                                 (clk_cpu                                                                   ), //i
    .reset_cpu                                               (reset_cpu                                                                 ), //i
    .clk_ram_bus                                             (clk_ram_bus                                                               ), //i
    .ram_axi_cc_toplevel_board_ctrl_reset_cpu_synchronized_1 (io_input_arw_queue_ram_axi_cc_toplevel_board_ctrl_reset_cpu_synchronized_1)  //o
  );
  StreamFifoCC_1 io_output_r_queue (
    .io_push_valid                                           (io_output_r_valid                                                        ), //i
    .io_push_ready                                           (io_output_r_queue_io_push_ready                                          ), //o
    .io_push_payload_data                                    (io_output_r_payload_data[63:0]                                           ), //i
    .io_push_payload_id                                      (io_output_r_payload_id[2:0]                                              ), //i
    .io_push_payload_resp                                    (io_output_r_payload_resp[1:0]                                            ), //i
    .io_push_payload_last                                    (io_output_r_payload_last                                                 ), //i
    .io_pop_valid                                            (io_output_r_queue_io_pop_valid                                           ), //o
    .io_pop_ready                                            (io_input_r_ready                                                         ), //i
    .io_pop_payload_data                                     (io_output_r_queue_io_pop_payload_data[63:0]                              ), //o
    .io_pop_payload_id                                       (io_output_r_queue_io_pop_payload_id[2:0]                                 ), //o
    .io_pop_payload_resp                                     (io_output_r_queue_io_pop_payload_resp[1:0]                               ), //o
    .io_pop_payload_last                                     (io_output_r_queue_io_pop_payload_last                                    ), //o
    .io_pushOccupancy                                        (io_output_r_queue_io_pushOccupancy[7:0]                                  ), //o
    .io_popOccupancy                                         (io_output_r_queue_io_popOccupancy[7:0]                                   ), //o
    .clk_ram_bus                                             (clk_ram_bus                                                              ), //i
    .reset_ram                                               (reset_ram                                                                ), //i
    .clk_cpu                                                 (clk_cpu                                                                  ), //i
    .ram_axi_cc_toplevel_board_ctrl_reset_ram_synchronized_1 (io_output_r_queue_ram_axi_cc_toplevel_board_ctrl_reset_ram_synchronized_1)  //o
  );
  StreamFifoCC_2 io_input_w_queue (
    .io_push_valid                                           (io_input_w_valid                                                          ), //i
    .io_push_ready                                           (io_input_w_queue_io_push_ready                                            ), //o
    .io_push_payload_data                                    (io_input_w_payload_data[63:0]                                             ), //i
    .io_push_payload_strb                                    (io_input_w_payload_strb[7:0]                                              ), //i
    .io_push_payload_last                                    (io_input_w_payload_last                                                   ), //i
    .io_pop_valid                                            (io_input_w_queue_io_pop_valid                                             ), //o
    .io_pop_ready                                            (io_output_w_ready                                                         ), //i
    .io_pop_payload_data                                     (io_input_w_queue_io_pop_payload_data[63:0]                                ), //o
    .io_pop_payload_strb                                     (io_input_w_queue_io_pop_payload_strb[7:0]                                 ), //o
    .io_pop_payload_last                                     (io_input_w_queue_io_pop_payload_last                                      ), //o
    .io_pushOccupancy                                        (io_input_w_queue_io_pushOccupancy[4:0]                                    ), //o
    .io_popOccupancy                                         (io_input_w_queue_io_popOccupancy[4:0]                                     ), //o
    .clk_cpu                                                 (clk_cpu                                                                   ), //i
    .reset_cpu                                               (reset_cpu                                                                 ), //i
    .clk_ram_bus                                             (clk_ram_bus                                                               ), //i
    .ram_axi_cc_toplevel_board_ctrl_reset_cpu_synchronized_1 (io_input_arw_queue_ram_axi_cc_toplevel_board_ctrl_reset_cpu_synchronized_1)  //i
  );
  StreamFifoCC_3 io_output_b_queue (
    .io_push_valid                                           (io_output_b_valid                                                        ), //i
    .io_push_ready                                           (io_output_b_queue_io_push_ready                                          ), //o
    .io_push_payload_id                                      (io_output_b_payload_id[2:0]                                              ), //i
    .io_push_payload_resp                                    (io_output_b_payload_resp[1:0]                                            ), //i
    .io_pop_valid                                            (io_output_b_queue_io_pop_valid                                           ), //o
    .io_pop_ready                                            (io_input_b_ready                                                         ), //i
    .io_pop_payload_id                                       (io_output_b_queue_io_pop_payload_id[2:0]                                 ), //o
    .io_pop_payload_resp                                     (io_output_b_queue_io_pop_payload_resp[1:0]                               ), //o
    .io_pushOccupancy                                        (io_output_b_queue_io_pushOccupancy[1:0]                                  ), //o
    .io_popOccupancy                                         (io_output_b_queue_io_popOccupancy[1:0]                                   ), //o
    .clk_ram_bus                                             (clk_ram_bus                                                              ), //i
    .reset_ram                                               (reset_ram                                                                ), //i
    .clk_cpu                                                 (clk_cpu                                                                  ), //i
    .ram_axi_cc_toplevel_board_ctrl_reset_ram_synchronized_1 (io_output_r_queue_ram_axi_cc_toplevel_board_ctrl_reset_ram_synchronized_1)  //i
  );
  assign io_input_arw_ready = io_input_arw_queue_io_push_ready;
  assign io_output_arw_valid = io_input_arw_queue_io_pop_valid;
  assign io_output_arw_payload_addr = io_input_arw_queue_io_pop_payload_addr;
  assign io_output_arw_payload_id = io_input_arw_queue_io_pop_payload_id;
  assign io_output_arw_payload_len = io_input_arw_queue_io_pop_payload_len;
  assign io_output_arw_payload_size = io_input_arw_queue_io_pop_payload_size;
  assign io_output_arw_payload_burst = io_input_arw_queue_io_pop_payload_burst;
  assign io_output_arw_payload_allStrb = io_input_arw_queue_io_pop_payload_allStrb;
  assign io_output_arw_payload_write = io_input_arw_queue_io_pop_payload_write;
  assign io_output_r_ready = io_output_r_queue_io_push_ready;
  assign io_input_r_valid = io_output_r_queue_io_pop_valid;
  assign io_input_r_payload_data = io_output_r_queue_io_pop_payload_data;
  assign io_input_r_payload_id = io_output_r_queue_io_pop_payload_id;
  assign io_input_r_payload_resp = io_output_r_queue_io_pop_payload_resp;
  assign io_input_r_payload_last = io_output_r_queue_io_pop_payload_last;
  assign io_input_w_ready = io_input_w_queue_io_push_ready;
  assign io_output_w_valid = io_input_w_queue_io_pop_valid;
  assign io_output_w_payload_data = io_input_w_queue_io_pop_payload_data;
  assign io_output_w_payload_strb = io_input_w_queue_io_pop_payload_strb;
  assign io_output_w_payload_last = io_input_w_queue_io_pop_payload_last;
  assign io_output_b_ready = io_output_b_queue_io_push_ready;
  assign io_input_b_valid = io_output_b_queue_io_pop_valid;
  assign io_input_b_payload_id = io_output_b_queue_io_pop_payload_id;
  assign io_input_b_payload_resp = io_output_b_queue_io_pop_payload_resp;

endmodule

module StreamArbiter_9 (
  input  wire          io_inputs_0_valid,
  output wire          io_inputs_0_ready,
  input  wire [26:0]   io_inputs_0_payload_addr,
  input  wire [2:0]    io_inputs_0_payload_id,
  input  wire [7:0]    io_inputs_0_payload_len,
  input  wire [2:0]    io_inputs_0_payload_size,
  input  wire [1:0]    io_inputs_0_payload_burst,
  input  wire          io_inputs_0_payload_allStrb,
  input  wire          io_inputs_1_valid,
  output wire          io_inputs_1_ready,
  input  wire [26:0]   io_inputs_1_payload_addr,
  input  wire [2:0]    io_inputs_1_payload_id,
  input  wire [7:0]    io_inputs_1_payload_len,
  input  wire [2:0]    io_inputs_1_payload_size,
  input  wire [1:0]    io_inputs_1_payload_burst,
  input  wire          io_inputs_1_payload_allStrb,
  output wire          io_output_valid,
  input  wire          io_output_ready,
  output wire [26:0]   io_output_payload_addr,
  output wire [2:0]    io_output_payload_id,
  output wire [7:0]    io_output_payload_len,
  output wire [2:0]    io_output_payload_size,
  output wire [1:0]    io_output_payload_burst,
  output wire          io_output_payload_allStrb,
  output wire [0:0]    io_chosen,
  output wire [1:0]    io_chosenOH,
  input  wire          clk_cpu,
  input  wire          reset_cpu
);

  wire       [3:0]    _zz__zz_maskProposal_0_2;
  wire       [3:0]    _zz__zz_maskProposal_0_2_1;
  wire       [1:0]    _zz__zz_maskProposal_0_2_2;
  reg                 locked;
  wire                maskProposal_0;
  wire                maskProposal_1;
  reg                 maskLocked_0;
  reg                 maskLocked_1;
  wire                maskRouted_0;
  wire                maskRouted_1;
  wire       [1:0]    _zz_maskProposal_0;
  wire       [3:0]    _zz_maskProposal_0_1;
  wire       [3:0]    _zz_maskProposal_0_2;
  wire       [1:0]    _zz_maskProposal_0_3;
  wire                io_output_fire;
  wire                _zz_io_chosen;

  assign _zz__zz_maskProposal_0_2 = (_zz_maskProposal_0_1 - _zz__zz_maskProposal_0_2_1);
  assign _zz__zz_maskProposal_0_2_2 = {maskLocked_0,maskLocked_1};
  assign _zz__zz_maskProposal_0_2_1 = {2'd0, _zz__zz_maskProposal_0_2_2};
  assign maskRouted_0 = (locked ? maskLocked_0 : maskProposal_0);
  assign maskRouted_1 = (locked ? maskLocked_1 : maskProposal_1);
  assign _zz_maskProposal_0 = {io_inputs_1_valid,io_inputs_0_valid};
  assign _zz_maskProposal_0_1 = {_zz_maskProposal_0,_zz_maskProposal_0};
  assign _zz_maskProposal_0_2 = (_zz_maskProposal_0_1 & (~ _zz__zz_maskProposal_0_2));
  assign _zz_maskProposal_0_3 = (_zz_maskProposal_0_2[3 : 2] | _zz_maskProposal_0_2[1 : 0]);
  assign maskProposal_0 = _zz_maskProposal_0_3[0];
  assign maskProposal_1 = _zz_maskProposal_0_3[1];
  assign io_output_fire = (io_output_valid && io_output_ready);
  assign io_output_valid = ((io_inputs_0_valid && maskRouted_0) || (io_inputs_1_valid && maskRouted_1));
  assign io_output_payload_addr = (maskRouted_0 ? io_inputs_0_payload_addr : io_inputs_1_payload_addr);
  assign io_output_payload_id = (maskRouted_0 ? io_inputs_0_payload_id : io_inputs_1_payload_id);
  assign io_output_payload_len = (maskRouted_0 ? io_inputs_0_payload_len : io_inputs_1_payload_len);
  assign io_output_payload_size = (maskRouted_0 ? io_inputs_0_payload_size : io_inputs_1_payload_size);
  assign io_output_payload_burst = (maskRouted_0 ? io_inputs_0_payload_burst : io_inputs_1_payload_burst);
  assign io_output_payload_allStrb = (maskRouted_0 ? io_inputs_0_payload_allStrb : io_inputs_1_payload_allStrb);
  assign io_inputs_0_ready = (maskRouted_0 && io_output_ready);
  assign io_inputs_1_ready = (maskRouted_1 && io_output_ready);
  assign io_chosenOH = {maskRouted_1,maskRouted_0};
  assign _zz_io_chosen = io_chosenOH[1];
  assign io_chosen = _zz_io_chosen;
  always @(posedge clk_cpu or posedge reset_cpu) begin
    if(reset_cpu) begin
      locked <= 1'b0;
      maskLocked_0 <= 1'b0;
      maskLocked_1 <= 1'b1;
    end else begin
      if(io_output_valid) begin
        maskLocked_0 <= maskRouted_0;
        maskLocked_1 <= maskRouted_1;
      end
      if(io_output_valid) begin
        locked <= 1'b1;
      end
      if(io_output_fire) begin
        locked <= 1'b0;
      end
    end
  end


endmodule

module WidthAdapter (
  input  wire          io_up_a_valid,
  output wire          io_up_a_ready,
  input  wire [2:0]    io_up_a_payload_opcode,
  input  wire [2:0]    io_up_a_payload_param,
  input  wire [31:0]   io_up_a_payload_address,
  input  wire [1:0]    io_up_a_payload_size,
  input  wire [3:0]    io_up_a_payload_mask,
  input  wire [31:0]   io_up_a_payload_data,
  input  wire          io_up_a_payload_corrupt,
  output wire          io_up_d_valid,
  input  wire          io_up_d_ready,
  output wire [2:0]    io_up_d_payload_opcode,
  output wire [2:0]    io_up_d_payload_param,
  output wire [1:0]    io_up_d_payload_size,
  output wire          io_up_d_payload_denied,
  output wire [31:0]   io_up_d_payload_data,
  output wire          io_up_d_payload_corrupt,
  output wire          io_down_a_valid,
  input  wire          io_down_a_ready,
  output wire [2:0]    io_down_a_payload_opcode,
  output wire [2:0]    io_down_a_payload_param,
  output wire [31:0]   io_down_a_payload_address,
  output wire [1:0]    io_down_a_payload_size,
  output wire [7:0]    io_down_a_payload_mask,
  output wire [63:0]   io_down_a_payload_data,
  output wire          io_down_a_payload_corrupt,
  input  wire          io_down_d_valid,
  output wire          io_down_d_ready,
  input  wire [2:0]    io_down_d_payload_opcode,
  input  wire [2:0]    io_down_d_payload_param,
  input  wire [1:0]    io_down_d_payload_size,
  input  wire          io_down_d_payload_denied,
  input  wire [63:0]   io_down_d_payload_data,
  input  wire          io_down_d_payload_corrupt,
  input  wire          clk_cpu,
  input  wire          reset_cpu
);
  localparam A_PUT_FULL_DATA = 3'd0;
  localparam A_PUT_PARTIAL_DATA = 3'd1;
  localparam A_GET = 3'd4;
  localparam A_ACQUIRE_BLOCK = 3'd6;
  localparam A_ACQUIRE_PERM = 3'd7;
  localparam D_ACCESS_ACK = 3'd0;
  localparam D_ACCESS_ACK_DATA = 3'd1;
  localparam D_GRANT = 3'd4;
  localparam D_GRANT_DATA = 3'd5;
  localparam D_RELEASE_ACK = 3'd6;

  wire                upsize_d_ctx_io_add_valid;
  wire       [0:0]    upsize_d_ctx_io_add_payload_context;
  wire                upsize_d_ctx_io_remove_valid;
  wire                upsize_d_ctx_io_add_ready;
  wire       [0:0]    upsize_d_ctx_io_query_context;
  reg        [31:0]   _zz_io_up_d_payload_data;
  reg                 upsize_iaHalt;
  wire                _zz_io_up_a_ready;
  wire                upsize_ia_valid;
  wire                upsize_ia_ready;
  wire       [2:0]    upsize_ia_payload_opcode;
  wire       [2:0]    upsize_ia_payload_param;
  wire       [31:0]   upsize_ia_payload_address;
  wire       [1:0]    upsize_ia_payload_size;
  wire       [3:0]    upsize_ia_payload_mask;
  wire       [31:0]   upsize_ia_payload_data;
  wire                upsize_ia_payload_corrupt;
  wire       [0:0]    _zz_upsize_a_ctrl_wordLast;
  wire                upsize_a_ctrl_burstLast;
  wire                upsize_ia_fire;
  wire                upsize_a_ctrl_wordLast;
  reg                 upsize_a_ctrl_buffer_valid;
  reg                 upsize_a_ctrl_buffer_first;
  reg        [2:0]    upsize_a_ctrl_buffer_args_opcode;
  reg        [2:0]    upsize_a_ctrl_buffer_args_param;
  reg        [31:0]   upsize_a_ctrl_buffer_args_address;
  reg        [1:0]    upsize_a_ctrl_buffer_args_size;
  reg        [31:0]   upsize_a_ctrl_buffer_data_0;
  reg        [31:0]   upsize_a_ctrl_buffer_data_1;
  reg        [3:0]    upsize_a_ctrl_buffer_mask_0;
  reg        [3:0]    upsize_a_ctrl_buffer_mask_1;
  reg                 upsize_a_ctrl_buffer_corrupt;
  wire       [1:0]    _zz_1;
  wire       [1:0]    _zz_2;
  wire                io_up_a_fire;
  wire                io_up_a_tracker_last;
  wire                when_ContextBuffer_l19;
  wire                io_up_d_fire;
  wire                upsize_d_ctrl_burstLast;
  reg        [0:0]    upsize_d_ctrl_counter;
  wire       [0:0]    upsize_d_ctrl_sel;
  `ifndef SYNTHESIS
  reg [127:0] io_up_a_payload_opcode_string;
  reg [119:0] io_up_d_payload_opcode_string;
  reg [127:0] io_down_a_payload_opcode_string;
  reg [119:0] io_down_d_payload_opcode_string;
  reg [127:0] upsize_ia_payload_opcode_string;
  reg [127:0] upsize_a_ctrl_buffer_args_opcode_string;
  `endif


  ContextAsyncBufferFull_1 upsize_d_ctx (
    .io_add_valid           (upsize_d_ctx_io_add_valid          ), //i
    .io_add_ready           (upsize_d_ctx_io_add_ready          ), //o
    .io_add_payload_context (upsize_d_ctx_io_add_payload_context), //i
    .io_remove_valid        (upsize_d_ctx_io_remove_valid       ), //i
    .io_query_context       (upsize_d_ctx_io_query_context      ), //o
    .clk_cpu                (clk_cpu                            ), //i
    .reset_cpu              (reset_cpu                          )  //i
  );
  always @(*) begin
    case(upsize_d_ctrl_sel)
      1'b0 : _zz_io_up_d_payload_data = io_down_d_payload_data[31 : 0];
      default : _zz_io_up_d_payload_data = io_down_d_payload_data[63 : 32];
    endcase
  end

  `ifndef SYNTHESIS
  always @(*) begin
    case(io_up_a_payload_opcode)
      A_PUT_FULL_DATA : io_up_a_payload_opcode_string = "PUT_FULL_DATA   ";
      A_PUT_PARTIAL_DATA : io_up_a_payload_opcode_string = "PUT_PARTIAL_DATA";
      A_GET : io_up_a_payload_opcode_string = "GET             ";
      A_ACQUIRE_BLOCK : io_up_a_payload_opcode_string = "ACQUIRE_BLOCK   ";
      A_ACQUIRE_PERM : io_up_a_payload_opcode_string = "ACQUIRE_PERM    ";
      default : io_up_a_payload_opcode_string = "????????????????";
    endcase
  end
  always @(*) begin
    case(io_up_d_payload_opcode)
      D_ACCESS_ACK : io_up_d_payload_opcode_string = "ACCESS_ACK     ";
      D_ACCESS_ACK_DATA : io_up_d_payload_opcode_string = "ACCESS_ACK_DATA";
      D_GRANT : io_up_d_payload_opcode_string = "GRANT          ";
      D_GRANT_DATA : io_up_d_payload_opcode_string = "GRANT_DATA     ";
      D_RELEASE_ACK : io_up_d_payload_opcode_string = "RELEASE_ACK    ";
      default : io_up_d_payload_opcode_string = "???????????????";
    endcase
  end
  always @(*) begin
    case(io_down_a_payload_opcode)
      A_PUT_FULL_DATA : io_down_a_payload_opcode_string = "PUT_FULL_DATA   ";
      A_PUT_PARTIAL_DATA : io_down_a_payload_opcode_string = "PUT_PARTIAL_DATA";
      A_GET : io_down_a_payload_opcode_string = "GET             ";
      A_ACQUIRE_BLOCK : io_down_a_payload_opcode_string = "ACQUIRE_BLOCK   ";
      A_ACQUIRE_PERM : io_down_a_payload_opcode_string = "ACQUIRE_PERM    ";
      default : io_down_a_payload_opcode_string = "????????????????";
    endcase
  end
  always @(*) begin
    case(io_down_d_payload_opcode)
      D_ACCESS_ACK : io_down_d_payload_opcode_string = "ACCESS_ACK     ";
      D_ACCESS_ACK_DATA : io_down_d_payload_opcode_string = "ACCESS_ACK_DATA";
      D_GRANT : io_down_d_payload_opcode_string = "GRANT          ";
      D_GRANT_DATA : io_down_d_payload_opcode_string = "GRANT_DATA     ";
      D_RELEASE_ACK : io_down_d_payload_opcode_string = "RELEASE_ACK    ";
      default : io_down_d_payload_opcode_string = "???????????????";
    endcase
  end
  always @(*) begin
    case(upsize_ia_payload_opcode)
      A_PUT_FULL_DATA : upsize_ia_payload_opcode_string = "PUT_FULL_DATA   ";
      A_PUT_PARTIAL_DATA : upsize_ia_payload_opcode_string = "PUT_PARTIAL_DATA";
      A_GET : upsize_ia_payload_opcode_string = "GET             ";
      A_ACQUIRE_BLOCK : upsize_ia_payload_opcode_string = "ACQUIRE_BLOCK   ";
      A_ACQUIRE_PERM : upsize_ia_payload_opcode_string = "ACQUIRE_PERM    ";
      default : upsize_ia_payload_opcode_string = "????????????????";
    endcase
  end
  always @(*) begin
    case(upsize_a_ctrl_buffer_args_opcode)
      A_PUT_FULL_DATA : upsize_a_ctrl_buffer_args_opcode_string = "PUT_FULL_DATA   ";
      A_PUT_PARTIAL_DATA : upsize_a_ctrl_buffer_args_opcode_string = "PUT_PARTIAL_DATA";
      A_GET : upsize_a_ctrl_buffer_args_opcode_string = "GET             ";
      A_ACQUIRE_BLOCK : upsize_a_ctrl_buffer_args_opcode_string = "ACQUIRE_BLOCK   ";
      A_ACQUIRE_PERM : upsize_a_ctrl_buffer_args_opcode_string = "ACQUIRE_PERM    ";
      default : upsize_a_ctrl_buffer_args_opcode_string = "????????????????";
    endcase
  end
  `endif

  always @(*) begin
    upsize_iaHalt = 1'b0;
    if(when_ContextBuffer_l19) begin
      upsize_iaHalt = 1'b1;
    end
  end

  assign _zz_io_up_a_ready = (! upsize_iaHalt);
  assign upsize_ia_valid = (io_up_a_valid && _zz_io_up_a_ready);
  assign io_up_a_ready = (upsize_ia_ready && _zz_io_up_a_ready);
  assign upsize_ia_payload_opcode = io_up_a_payload_opcode;
  assign upsize_ia_payload_param = io_up_a_payload_param;
  assign upsize_ia_payload_address = io_up_a_payload_address;
  assign upsize_ia_payload_size = io_up_a_payload_size;
  assign upsize_ia_payload_mask = io_up_a_payload_mask;
  assign upsize_ia_payload_data = io_up_a_payload_data;
  assign upsize_ia_payload_corrupt = io_up_a_payload_corrupt;
  assign _zz_upsize_a_ctrl_wordLast = upsize_ia_payload_address[2 : 2];
  assign upsize_a_ctrl_burstLast = ((! ((1'b0 || (A_PUT_FULL_DATA == upsize_ia_payload_opcode)) || (A_PUT_PARTIAL_DATA == upsize_ia_payload_opcode))) || 1'b1);
  assign upsize_ia_fire = (upsize_ia_valid && upsize_ia_ready);
  assign upsize_a_ctrl_wordLast = ((&_zz_upsize_a_ctrl_wordLast) || upsize_a_ctrl_burstLast);
  assign io_down_a_valid = upsize_a_ctrl_buffer_valid;
  assign io_down_a_payload_opcode = upsize_a_ctrl_buffer_args_opcode;
  assign io_down_a_payload_param = upsize_a_ctrl_buffer_args_param;
  assign io_down_a_payload_address = upsize_a_ctrl_buffer_args_address;
  assign io_down_a_payload_size = upsize_a_ctrl_buffer_args_size;
  assign io_down_a_payload_mask = {upsize_a_ctrl_buffer_mask_1,upsize_a_ctrl_buffer_mask_0};
  assign io_down_a_payload_data = {upsize_a_ctrl_buffer_data_1,upsize_a_ctrl_buffer_data_0};
  assign io_down_a_payload_corrupt = upsize_a_ctrl_buffer_corrupt;
  assign upsize_ia_ready = ((! upsize_a_ctrl_buffer_valid) || io_down_a_ready);
  assign _zz_1 = ({1'd0,1'b1} <<< _zz_upsize_a_ctrl_wordLast);
  assign _zz_2 = ({1'd0,1'b1} <<< _zz_upsize_a_ctrl_wordLast);
  assign io_up_a_fire = (io_up_a_valid && io_up_a_ready);
  assign io_up_a_tracker_last = ((! ((1'b0 || (A_PUT_FULL_DATA == io_up_a_payload_opcode)) || (A_PUT_PARTIAL_DATA == io_up_a_payload_opcode))) || 1'b1);
  assign upsize_d_ctx_io_add_valid = (io_up_a_fire && io_up_a_tracker_last);
  assign when_ContextBuffer_l19 = (! upsize_d_ctx_io_add_ready);
  assign io_up_d_fire = (io_up_d_valid && io_up_d_ready);
  assign upsize_d_ctrl_burstLast = ((! ((1'b0 || (D_ACCESS_ACK_DATA == io_up_d_payload_opcode)) || (D_GRANT_DATA == io_up_d_payload_opcode))) || 1'b1);
  assign upsize_d_ctx_io_remove_valid = ((io_up_d_fire && upsize_d_ctrl_burstLast) && (|{(io_up_d_payload_opcode == D_GRANT_DATA),{(io_up_d_payload_opcode == D_GRANT),{(io_up_d_payload_opcode == D_ACCESS_ACK_DATA),(io_up_d_payload_opcode == D_ACCESS_ACK)}}}));
  assign upsize_d_ctx_io_add_payload_context = io_up_a_payload_address[2 : 2];
  assign upsize_d_ctrl_sel = (upsize_d_ctrl_counter + upsize_d_ctx_io_query_context);
  assign io_up_d_valid = io_down_d_valid;
  assign io_up_d_payload_opcode = io_down_d_payload_opcode;
  assign io_up_d_payload_param = io_down_d_payload_param;
  assign io_up_d_payload_size = io_down_d_payload_size;
  assign io_up_d_payload_denied = io_down_d_payload_denied;
  assign io_up_d_payload_corrupt = io_down_d_payload_corrupt;
  assign io_down_d_ready = (io_up_d_ready && ((&upsize_d_ctrl_counter) || upsize_d_ctrl_burstLast));
  assign io_up_d_payload_data = _zz_io_up_d_payload_data;
  always @(posedge clk_cpu or posedge reset_cpu) begin
    if(reset_cpu) begin
      upsize_a_ctrl_buffer_valid <= 1'b0;
      upsize_a_ctrl_buffer_first <= 1'b1;
      upsize_d_ctrl_counter <= 1'b0;
    end else begin
      if(io_down_a_ready) begin
        upsize_a_ctrl_buffer_valid <= 1'b0;
      end
      if(upsize_ia_fire) begin
        upsize_a_ctrl_buffer_valid <= upsize_a_ctrl_wordLast;
        upsize_a_ctrl_buffer_first <= upsize_a_ctrl_wordLast;
      end
      if(io_up_d_fire) begin
        upsize_d_ctrl_counter <= (upsize_d_ctrl_counter + 1'b1);
        if(upsize_d_ctrl_burstLast) begin
          upsize_d_ctrl_counter <= 1'b0;
        end
      end
    end
  end

  always @(posedge clk_cpu) begin
    if(upsize_ia_fire) begin
      if(upsize_a_ctrl_buffer_first) begin
        upsize_a_ctrl_buffer_args_opcode <= upsize_ia_payload_opcode;
        upsize_a_ctrl_buffer_args_param <= upsize_ia_payload_param;
        upsize_a_ctrl_buffer_args_address <= upsize_ia_payload_address;
        upsize_a_ctrl_buffer_args_size <= upsize_ia_payload_size;
        upsize_a_ctrl_buffer_corrupt <= 1'b0;
        upsize_a_ctrl_buffer_mask_0 <= 4'b0000;
        upsize_a_ctrl_buffer_mask_1 <= 4'b0000;
      end
      if(_zz_1[0]) begin
        upsize_a_ctrl_buffer_data_0 <= upsize_ia_payload_data;
      end
      if(_zz_1[1]) begin
        upsize_a_ctrl_buffer_data_1 <= upsize_ia_payload_data;
      end
      if(_zz_2[0]) begin
        upsize_a_ctrl_buffer_mask_0 <= upsize_ia_payload_mask;
      end
      if(_zz_2[1]) begin
        upsize_a_ctrl_buffer_mask_1 <= upsize_ia_payload_mask;
      end
      if(upsize_ia_payload_corrupt) begin
        upsize_a_ctrl_buffer_corrupt <= 1'b1;
      end
    end
  end


endmodule

module Axi4Bridge (
  input  wire          io_up_a_valid,
  output wire          io_up_a_ready,
  input  wire [2:0]    io_up_a_payload_opcode,
  input  wire [2:0]    io_up_a_payload_param,
  input  wire [2:0]    io_up_a_payload_source,
  input  wire [26:0]   io_up_a_payload_address,
  input  wire [2:0]    io_up_a_payload_size,
  input  wire [7:0]    io_up_a_payload_mask,
  input  wire [63:0]   io_up_a_payload_data,
  input  wire          io_up_a_payload_corrupt,
  output wire          io_up_d_valid,
  input  wire          io_up_d_ready,
  output wire [2:0]    io_up_d_payload_opcode,
  output wire [2:0]    io_up_d_payload_param,
  output wire [2:0]    io_up_d_payload_source,
  output wire [2:0]    io_up_d_payload_size,
  output wire          io_up_d_payload_denied,
  output wire [63:0]   io_up_d_payload_data,
  output wire          io_up_d_payload_corrupt,
  output wire          io_down_aw_valid,
  input  wire          io_down_aw_ready,
  output wire [26:0]   io_down_aw_payload_addr,
  output wire [2:0]    io_down_aw_payload_id,
  output wire [7:0]    io_down_aw_payload_len,
  output wire [2:0]    io_down_aw_payload_size,
  output wire [1:0]    io_down_aw_payload_burst,
  output wire          io_down_aw_payload_allStrb,
  output wire          io_down_w_valid,
  input  wire          io_down_w_ready,
  output wire [63:0]   io_down_w_payload_data,
  output wire [7:0]    io_down_w_payload_strb,
  output wire          io_down_w_payload_last,
  input  wire          io_down_b_valid,
  output wire          io_down_b_ready,
  input  wire [2:0]    io_down_b_payload_id,
  input  wire [1:0]    io_down_b_payload_resp,
  output wire          io_down_ar_valid,
  input  wire          io_down_ar_ready,
  output wire [26:0]   io_down_ar_payload_addr,
  output wire [2:0]    io_down_ar_payload_id,
  output wire [7:0]    io_down_ar_payload_len,
  output wire [2:0]    io_down_ar_payload_size,
  output wire [1:0]    io_down_ar_payload_burst,
  input  wire          io_down_r_valid,
  output wire          io_down_r_ready,
  input  wire [63:0]   io_down_r_payload_data,
  input  wire [2:0]    io_down_r_payload_id,
  input  wire [1:0]    io_down_r_payload_resp,
  input  wire          io_down_r_payload_last,
  input  wire          clk_cpu,
  input  wire          reset_cpu
);
  localparam A_PUT_FULL_DATA = 3'd0;
  localparam A_PUT_PARTIAL_DATA = 3'd1;
  localparam A_GET = 3'd4;
  localparam A_ACQUIRE_BLOCK = 3'd6;
  localparam A_ACQUIRE_PERM = 3'd7;
  localparam D_ACCESS_ACK = 3'd0;
  localparam D_ACCESS_ACK_DATA = 3'd1;
  localparam D_GRANT = 3'd4;
  localparam D_GRANT_DATA = 3'd5;
  localparam D_RELEASE_ACK = 3'd6;

  wire                a_ctx_io_add_valid;
  wire                a_ctx_io_remove_valid;
  wire                d_arbiter_io_inputs_0_payload_denied;
  wire                d_arbiter_io_inputs_1_payload_denied;
  wire                a_ctx_io_add_ready;
  wire       [2:0]    a_ctx_io_query_context;
  wire                d_arbiter_io_inputs_0_ready;
  wire                d_arbiter_io_inputs_1_ready;
  wire                d_arbiter_io_output_valid;
  wire       [2:0]    d_arbiter_io_output_payload_source;
  wire                d_arbiter_io_output_payload_denied;
  wire                d_arbiter_io_output_payload_last;
  wire       [0:0]    d_arbiter_io_chosen;
  wire       [1:0]    d_arbiter_io_chosenOH;
  reg        [2:0]    _zz_io_up_a_tracker_last;
  reg        [2:0]    _zz_io_up_d_tracker_last;
  reg        [2:0]    _zz_a_cmdFork_tracker_last;
  reg        [2:0]    _zz_a_cmd_len;
  reg        [2:0]    _zz_a_cmd_sizePerBeat;
  reg        [2:0]    _zz_a_data_buffer_tracker_last;
  reg                 a_ctxFull;
  wire                _zz_io_up_a_ready;
  wire                a_halted_valid;
  reg                 a_halted_ready;
  wire       [2:0]    a_halted_payload_opcode;
  wire       [2:0]    a_halted_payload_param;
  wire       [2:0]    a_halted_payload_source;
  wire       [26:0]   a_halted_payload_address;
  wire       [2:0]    a_halted_payload_size;
  wire       [7:0]    a_halted_payload_mask;
  wire       [63:0]   a_halted_payload_data;
  wire                a_halted_payload_corrupt;
  wire                io_up_a_fire;
  reg        [2:0]    io_up_a_tracker_beat;
  wire                io_up_a_tracker_last;
  wire                when_ContextBuffer_l19;
  wire                io_up_d_fire;
  reg        [2:0]    io_up_d_tracker_beat;
  wire                io_up_d_tracker_last;
  wire                a_cmdFork_valid;
  reg                 a_cmdFork_ready;
  wire       [2:0]    a_cmdFork_payload_opcode;
  wire       [2:0]    a_cmdFork_payload_param;
  wire       [2:0]    a_cmdFork_payload_source;
  wire       [26:0]   a_cmdFork_payload_address;
  wire       [2:0]    a_cmdFork_payload_size;
  wire       [7:0]    a_cmdFork_payload_mask;
  wire       [63:0]   a_cmdFork_payload_data;
  wire                a_cmdFork_payload_corrupt;
  wire                a_dataFork_valid;
  reg                 a_dataFork_ready;
  wire       [2:0]    a_dataFork_payload_opcode;
  wire       [2:0]    a_dataFork_payload_param;
  wire       [2:0]    a_dataFork_payload_source;
  wire       [26:0]   a_dataFork_payload_address;
  wire       [2:0]    a_dataFork_payload_size;
  wire       [7:0]    a_dataFork_payload_mask;
  wire       [63:0]   a_dataFork_payload_data;
  wire                a_dataFork_payload_corrupt;
  reg                 a_halted_fork2_logic_linkEnable_0;
  reg                 a_halted_fork2_logic_linkEnable_1;
  wire                when_Stream_l1084;
  wire                when_Stream_l1084_1;
  wire                a_cmdFork_fire;
  wire                a_dataFork_fire;
  reg        [2:0]    a_cmdFork_tracker_beat;
  wire                a_cmdFork_tracker_last;
  wire                when_Stream_l466;
  reg                 a_cmd_filtred_valid;
  wire                a_cmd_filtred_ready;
  wire       [2:0]    a_cmd_filtred_payload_opcode;
  wire       [2:0]    a_cmd_filtred_payload_param;
  wire       [2:0]    a_cmd_filtred_payload_source;
  wire       [26:0]   a_cmd_filtred_payload_address;
  wire       [2:0]    a_cmd_filtred_payload_size;
  wire       [7:0]    a_cmd_filtred_payload_mask;
  wire       [63:0]   a_cmd_filtred_payload_data;
  wire                a_cmd_filtred_payload_corrupt;
  wire                a_cmd_buffered_valid;
  wire                a_cmd_buffered_ready;
  wire       [2:0]    a_cmd_buffered_payload_opcode;
  wire       [2:0]    a_cmd_buffered_payload_param;
  wire       [2:0]    a_cmd_buffered_payload_source;
  wire       [26:0]   a_cmd_buffered_payload_address;
  wire       [2:0]    a_cmd_buffered_payload_size;
  wire       [7:0]    a_cmd_buffered_payload_mask;
  wire       [63:0]   a_cmd_buffered_payload_data;
  wire                a_cmd_buffered_payload_corrupt;
  reg                 a_cmd_filtred_rValid;
  wire                a_cmd_buffered_fire;
  reg        [2:0]    a_cmd_filtred_rData_opcode;
  reg        [2:0]    a_cmd_filtred_rData_param;
  reg        [2:0]    a_cmd_filtred_rData_source;
  reg        [26:0]   a_cmd_filtred_rData_address;
  reg        [2:0]    a_cmd_filtred_rData_size;
  reg        [7:0]    a_cmd_filtred_rData_mask;
  reg        [63:0]   a_cmd_filtred_rData_data;
  reg                 a_cmd_filtred_rData_corrupt;
  wire                a_cmd_isGet;
  wire       [7:0]    a_cmd_len;
  wire       [2:0]    a_cmd_sizePerBeat;
  wire                when_Stream_l466_1;
  reg                 a_data_filtred_valid;
  reg                 a_data_filtred_ready;
  wire       [2:0]    a_data_filtred_payload_opcode;
  wire       [2:0]    a_data_filtred_payload_param;
  wire       [2:0]    a_data_filtred_payload_source;
  wire       [26:0]   a_data_filtred_payload_address;
  wire       [2:0]    a_data_filtred_payload_size;
  wire       [7:0]    a_data_filtred_payload_mask;
  wire       [63:0]   a_data_filtred_payload_data;
  wire                a_data_filtred_payload_corrupt;
  wire                a_data_buffer_valid;
  wire                a_data_buffer_ready;
  wire       [2:0]    a_data_buffer_payload_opcode;
  wire       [2:0]    a_data_buffer_payload_param;
  wire       [2:0]    a_data_buffer_payload_source;
  wire       [26:0]   a_data_buffer_payload_address;
  wire       [2:0]    a_data_buffer_payload_size;
  wire       [7:0]    a_data_buffer_payload_mask;
  wire       [63:0]   a_data_buffer_payload_data;
  wire                a_data_buffer_payload_corrupt;
  reg                 a_data_filtred_rValid;
  reg        [2:0]    a_data_filtred_rData_opcode;
  reg        [2:0]    a_data_filtred_rData_param;
  reg        [2:0]    a_data_filtred_rData_source;
  reg        [26:0]   a_data_filtred_rData_address;
  reg        [2:0]    a_data_filtred_rData_size;
  reg        [7:0]    a_data_filtred_rData_mask;
  reg        [63:0]   a_data_filtred_rData_data;
  reg                 a_data_filtred_rData_corrupt;
  wire                when_Stream_l393;
  reg        [2:0]    a_data_buffer_tracker_beat;
  wire                a_data_buffer_tracker_last;
  wire                a_data_buffer_fire;
  wire       [2:0]    _zz_io_up_d_payload_opcode;
  `ifndef SYNTHESIS
  reg [127:0] io_up_a_payload_opcode_string;
  reg [119:0] io_up_d_payload_opcode_string;
  reg [127:0] a_halted_payload_opcode_string;
  reg [127:0] a_cmdFork_payload_opcode_string;
  reg [127:0] a_dataFork_payload_opcode_string;
  reg [127:0] a_cmd_filtred_payload_opcode_string;
  reg [127:0] a_cmd_buffered_payload_opcode_string;
  reg [127:0] a_cmd_filtred_rData_opcode_string;
  reg [127:0] a_data_filtred_payload_opcode_string;
  reg [127:0] a_data_buffer_payload_opcode_string;
  reg [127:0] a_data_filtred_rData_opcode_string;
  reg [119:0] _zz_io_up_d_payload_opcode_string;
  `endif


  ContextAsyncBufferFull a_ctx (
    .io_add_valid           (a_ctx_io_add_valid         ), //i
    .io_add_ready           (a_ctx_io_add_ready         ), //o
    .io_add_payload_id      (io_up_a_payload_source[2:0]), //i
    .io_add_payload_context (io_up_a_payload_size[2:0]  ), //i
    .io_remove_valid        (a_ctx_io_remove_valid      ), //i
    .io_remove_payload_id   (io_up_d_payload_source[2:0]), //i
    .io_query_id            (io_up_d_payload_source[2:0]), //i
    .io_query_context       (a_ctx_io_query_context[2:0]), //o
    .clk_cpu                (clk_cpu                    ), //i
    .reset_cpu              (reset_cpu                  )  //i
  );
  StreamArbiter_6 d_arbiter (
    .io_inputs_0_valid          (io_down_b_valid                        ), //i
    .io_inputs_0_ready          (d_arbiter_io_inputs_0_ready            ), //o
    .io_inputs_0_payload_source (io_down_b_payload_id[2:0]              ), //i
    .io_inputs_0_payload_denied (d_arbiter_io_inputs_0_payload_denied   ), //i
    .io_inputs_0_payload_last   (1'b1                                   ), //i
    .io_inputs_1_valid          (io_down_r_valid                        ), //i
    .io_inputs_1_ready          (d_arbiter_io_inputs_1_ready            ), //o
    .io_inputs_1_payload_source (io_down_r_payload_id[2:0]              ), //i
    .io_inputs_1_payload_denied (d_arbiter_io_inputs_1_payload_denied   ), //i
    .io_inputs_1_payload_last   (io_down_r_payload_last                 ), //i
    .io_output_valid            (d_arbiter_io_output_valid              ), //o
    .io_output_ready            (io_up_d_ready                          ), //i
    .io_output_payload_source   (d_arbiter_io_output_payload_source[2:0]), //o
    .io_output_payload_denied   (d_arbiter_io_output_payload_denied     ), //o
    .io_output_payload_last     (d_arbiter_io_output_payload_last       ), //o
    .io_chosen                  (d_arbiter_io_chosen                    ), //o
    .io_chosenOH                (d_arbiter_io_chosenOH[1:0]             ), //o
    .clk_cpu                    (clk_cpu                                ), //i
    .reset_cpu                  (reset_cpu                              )  //i
  );
  always @(*) begin
    case(io_up_a_payload_size)
      3'b000 : _zz_io_up_a_tracker_last = 3'b000;
      3'b001 : _zz_io_up_a_tracker_last = 3'b000;
      3'b010 : _zz_io_up_a_tracker_last = 3'b000;
      3'b011 : _zz_io_up_a_tracker_last = 3'b000;
      3'b100 : _zz_io_up_a_tracker_last = 3'b001;
      3'b101 : _zz_io_up_a_tracker_last = 3'b011;
      default : _zz_io_up_a_tracker_last = 3'b111;
    endcase
  end

  always @(*) begin
    case(io_up_d_payload_size)
      3'b000 : _zz_io_up_d_tracker_last = 3'b000;
      3'b001 : _zz_io_up_d_tracker_last = 3'b000;
      3'b010 : _zz_io_up_d_tracker_last = 3'b000;
      3'b011 : _zz_io_up_d_tracker_last = 3'b000;
      3'b100 : _zz_io_up_d_tracker_last = 3'b001;
      3'b101 : _zz_io_up_d_tracker_last = 3'b011;
      default : _zz_io_up_d_tracker_last = 3'b111;
    endcase
  end

  always @(*) begin
    case(a_cmdFork_payload_size)
      3'b000 : _zz_a_cmdFork_tracker_last = 3'b000;
      3'b001 : _zz_a_cmdFork_tracker_last = 3'b000;
      3'b010 : _zz_a_cmdFork_tracker_last = 3'b000;
      3'b011 : _zz_a_cmdFork_tracker_last = 3'b000;
      3'b100 : _zz_a_cmdFork_tracker_last = 3'b001;
      3'b101 : _zz_a_cmdFork_tracker_last = 3'b011;
      default : _zz_a_cmdFork_tracker_last = 3'b111;
    endcase
  end

  always @(*) begin
    case(a_cmd_buffered_payload_size)
      3'b000 : begin
        _zz_a_cmd_len = 3'b000;
        _zz_a_cmd_sizePerBeat = 3'b000;
      end
      3'b001 : begin
        _zz_a_cmd_len = 3'b000;
        _zz_a_cmd_sizePerBeat = 3'b001;
      end
      3'b010 : begin
        _zz_a_cmd_len = 3'b000;
        _zz_a_cmd_sizePerBeat = 3'b010;
      end
      3'b011 : begin
        _zz_a_cmd_len = 3'b000;
        _zz_a_cmd_sizePerBeat = 3'b011;
      end
      3'b100 : begin
        _zz_a_cmd_len = 3'b001;
        _zz_a_cmd_sizePerBeat = 3'b011;
      end
      3'b101 : begin
        _zz_a_cmd_len = 3'b011;
        _zz_a_cmd_sizePerBeat = 3'b011;
      end
      default : begin
        _zz_a_cmd_len = 3'b111;
        _zz_a_cmd_sizePerBeat = 3'b011;
      end
    endcase
  end

  always @(*) begin
    case(a_data_buffer_payload_size)
      3'b000 : _zz_a_data_buffer_tracker_last = 3'b000;
      3'b001 : _zz_a_data_buffer_tracker_last = 3'b000;
      3'b010 : _zz_a_data_buffer_tracker_last = 3'b000;
      3'b011 : _zz_a_data_buffer_tracker_last = 3'b000;
      3'b100 : _zz_a_data_buffer_tracker_last = 3'b001;
      3'b101 : _zz_a_data_buffer_tracker_last = 3'b011;
      default : _zz_a_data_buffer_tracker_last = 3'b111;
    endcase
  end

  `ifndef SYNTHESIS
  always @(*) begin
    case(io_up_a_payload_opcode)
      A_PUT_FULL_DATA : io_up_a_payload_opcode_string = "PUT_FULL_DATA   ";
      A_PUT_PARTIAL_DATA : io_up_a_payload_opcode_string = "PUT_PARTIAL_DATA";
      A_GET : io_up_a_payload_opcode_string = "GET             ";
      A_ACQUIRE_BLOCK : io_up_a_payload_opcode_string = "ACQUIRE_BLOCK   ";
      A_ACQUIRE_PERM : io_up_a_payload_opcode_string = "ACQUIRE_PERM    ";
      default : io_up_a_payload_opcode_string = "????????????????";
    endcase
  end
  always @(*) begin
    case(io_up_d_payload_opcode)
      D_ACCESS_ACK : io_up_d_payload_opcode_string = "ACCESS_ACK     ";
      D_ACCESS_ACK_DATA : io_up_d_payload_opcode_string = "ACCESS_ACK_DATA";
      D_GRANT : io_up_d_payload_opcode_string = "GRANT          ";
      D_GRANT_DATA : io_up_d_payload_opcode_string = "GRANT_DATA     ";
      D_RELEASE_ACK : io_up_d_payload_opcode_string = "RELEASE_ACK    ";
      default : io_up_d_payload_opcode_string = "???????????????";
    endcase
  end
  always @(*) begin
    case(a_halted_payload_opcode)
      A_PUT_FULL_DATA : a_halted_payload_opcode_string = "PUT_FULL_DATA   ";
      A_PUT_PARTIAL_DATA : a_halted_payload_opcode_string = "PUT_PARTIAL_DATA";
      A_GET : a_halted_payload_opcode_string = "GET             ";
      A_ACQUIRE_BLOCK : a_halted_payload_opcode_string = "ACQUIRE_BLOCK   ";
      A_ACQUIRE_PERM : a_halted_payload_opcode_string = "ACQUIRE_PERM    ";
      default : a_halted_payload_opcode_string = "????????????????";
    endcase
  end
  always @(*) begin
    case(a_cmdFork_payload_opcode)
      A_PUT_FULL_DATA : a_cmdFork_payload_opcode_string = "PUT_FULL_DATA   ";
      A_PUT_PARTIAL_DATA : a_cmdFork_payload_opcode_string = "PUT_PARTIAL_DATA";
      A_GET : a_cmdFork_payload_opcode_string = "GET             ";
      A_ACQUIRE_BLOCK : a_cmdFork_payload_opcode_string = "ACQUIRE_BLOCK   ";
      A_ACQUIRE_PERM : a_cmdFork_payload_opcode_string = "ACQUIRE_PERM    ";
      default : a_cmdFork_payload_opcode_string = "????????????????";
    endcase
  end
  always @(*) begin
    case(a_dataFork_payload_opcode)
      A_PUT_FULL_DATA : a_dataFork_payload_opcode_string = "PUT_FULL_DATA   ";
      A_PUT_PARTIAL_DATA : a_dataFork_payload_opcode_string = "PUT_PARTIAL_DATA";
      A_GET : a_dataFork_payload_opcode_string = "GET             ";
      A_ACQUIRE_BLOCK : a_dataFork_payload_opcode_string = "ACQUIRE_BLOCK   ";
      A_ACQUIRE_PERM : a_dataFork_payload_opcode_string = "ACQUIRE_PERM    ";
      default : a_dataFork_payload_opcode_string = "????????????????";
    endcase
  end
  always @(*) begin
    case(a_cmd_filtred_payload_opcode)
      A_PUT_FULL_DATA : a_cmd_filtred_payload_opcode_string = "PUT_FULL_DATA   ";
      A_PUT_PARTIAL_DATA : a_cmd_filtred_payload_opcode_string = "PUT_PARTIAL_DATA";
      A_GET : a_cmd_filtred_payload_opcode_string = "GET             ";
      A_ACQUIRE_BLOCK : a_cmd_filtred_payload_opcode_string = "ACQUIRE_BLOCK   ";
      A_ACQUIRE_PERM : a_cmd_filtred_payload_opcode_string = "ACQUIRE_PERM    ";
      default : a_cmd_filtred_payload_opcode_string = "????????????????";
    endcase
  end
  always @(*) begin
    case(a_cmd_buffered_payload_opcode)
      A_PUT_FULL_DATA : a_cmd_buffered_payload_opcode_string = "PUT_FULL_DATA   ";
      A_PUT_PARTIAL_DATA : a_cmd_buffered_payload_opcode_string = "PUT_PARTIAL_DATA";
      A_GET : a_cmd_buffered_payload_opcode_string = "GET             ";
      A_ACQUIRE_BLOCK : a_cmd_buffered_payload_opcode_string = "ACQUIRE_BLOCK   ";
      A_ACQUIRE_PERM : a_cmd_buffered_payload_opcode_string = "ACQUIRE_PERM    ";
      default : a_cmd_buffered_payload_opcode_string = "????????????????";
    endcase
  end
  always @(*) begin
    case(a_cmd_filtred_rData_opcode)
      A_PUT_FULL_DATA : a_cmd_filtred_rData_opcode_string = "PUT_FULL_DATA   ";
      A_PUT_PARTIAL_DATA : a_cmd_filtred_rData_opcode_string = "PUT_PARTIAL_DATA";
      A_GET : a_cmd_filtred_rData_opcode_string = "GET             ";
      A_ACQUIRE_BLOCK : a_cmd_filtred_rData_opcode_string = "ACQUIRE_BLOCK   ";
      A_ACQUIRE_PERM : a_cmd_filtred_rData_opcode_string = "ACQUIRE_PERM    ";
      default : a_cmd_filtred_rData_opcode_string = "????????????????";
    endcase
  end
  always @(*) begin
    case(a_data_filtred_payload_opcode)
      A_PUT_FULL_DATA : a_data_filtred_payload_opcode_string = "PUT_FULL_DATA   ";
      A_PUT_PARTIAL_DATA : a_data_filtred_payload_opcode_string = "PUT_PARTIAL_DATA";
      A_GET : a_data_filtred_payload_opcode_string = "GET             ";
      A_ACQUIRE_BLOCK : a_data_filtred_payload_opcode_string = "ACQUIRE_BLOCK   ";
      A_ACQUIRE_PERM : a_data_filtred_payload_opcode_string = "ACQUIRE_PERM    ";
      default : a_data_filtred_payload_opcode_string = "????????????????";
    endcase
  end
  always @(*) begin
    case(a_data_buffer_payload_opcode)
      A_PUT_FULL_DATA : a_data_buffer_payload_opcode_string = "PUT_FULL_DATA   ";
      A_PUT_PARTIAL_DATA : a_data_buffer_payload_opcode_string = "PUT_PARTIAL_DATA";
      A_GET : a_data_buffer_payload_opcode_string = "GET             ";
      A_ACQUIRE_BLOCK : a_data_buffer_payload_opcode_string = "ACQUIRE_BLOCK   ";
      A_ACQUIRE_PERM : a_data_buffer_payload_opcode_string = "ACQUIRE_PERM    ";
      default : a_data_buffer_payload_opcode_string = "????????????????";
    endcase
  end
  always @(*) begin
    case(a_data_filtred_rData_opcode)
      A_PUT_FULL_DATA : a_data_filtred_rData_opcode_string = "PUT_FULL_DATA   ";
      A_PUT_PARTIAL_DATA : a_data_filtred_rData_opcode_string = "PUT_PARTIAL_DATA";
      A_GET : a_data_filtred_rData_opcode_string = "GET             ";
      A_ACQUIRE_BLOCK : a_data_filtred_rData_opcode_string = "ACQUIRE_BLOCK   ";
      A_ACQUIRE_PERM : a_data_filtred_rData_opcode_string = "ACQUIRE_PERM    ";
      default : a_data_filtred_rData_opcode_string = "????????????????";
    endcase
  end
  always @(*) begin
    case(_zz_io_up_d_payload_opcode)
      D_ACCESS_ACK : _zz_io_up_d_payload_opcode_string = "ACCESS_ACK     ";
      D_ACCESS_ACK_DATA : _zz_io_up_d_payload_opcode_string = "ACCESS_ACK_DATA";
      D_GRANT : _zz_io_up_d_payload_opcode_string = "GRANT          ";
      D_GRANT_DATA : _zz_io_up_d_payload_opcode_string = "GRANT_DATA     ";
      D_RELEASE_ACK : _zz_io_up_d_payload_opcode_string = "RELEASE_ACK    ";
      default : _zz_io_up_d_payload_opcode_string = "???????????????";
    endcase
  end
  `endif

  always @(*) begin
    a_ctxFull = 1'b0;
    if(when_ContextBuffer_l19) begin
      a_ctxFull = 1'b1;
    end
  end

  assign _zz_io_up_a_ready = (! a_ctxFull);
  assign a_halted_valid = (io_up_a_valid && _zz_io_up_a_ready);
  assign io_up_a_ready = (a_halted_ready && _zz_io_up_a_ready);
  assign a_halted_payload_opcode = io_up_a_payload_opcode;
  assign a_halted_payload_param = io_up_a_payload_param;
  assign a_halted_payload_source = io_up_a_payload_source;
  assign a_halted_payload_address = io_up_a_payload_address;
  assign a_halted_payload_size = io_up_a_payload_size;
  assign a_halted_payload_mask = io_up_a_payload_mask;
  assign a_halted_payload_data = io_up_a_payload_data;
  assign a_halted_payload_corrupt = io_up_a_payload_corrupt;
  assign io_up_a_fire = (io_up_a_valid && io_up_a_ready);
  assign io_up_a_tracker_last = ((! ((1'b0 || (A_PUT_FULL_DATA == io_up_a_payload_opcode)) || (A_PUT_PARTIAL_DATA == io_up_a_payload_opcode))) || (io_up_a_tracker_beat == _zz_io_up_a_tracker_last));
  assign a_ctx_io_add_valid = (io_up_a_fire && io_up_a_tracker_last);
  assign when_ContextBuffer_l19 = (! a_ctx_io_add_ready);
  assign io_up_d_fire = (io_up_d_valid && io_up_d_ready);
  assign io_up_d_tracker_last = ((! ((1'b0 || (D_ACCESS_ACK_DATA == io_up_d_payload_opcode)) || (D_GRANT_DATA == io_up_d_payload_opcode))) || (io_up_d_tracker_beat == _zz_io_up_d_tracker_last));
  assign a_ctx_io_remove_valid = ((io_up_d_fire && io_up_d_tracker_last) && (|{(io_up_d_payload_opcode == D_GRANT_DATA),{(io_up_d_payload_opcode == D_GRANT),{(io_up_d_payload_opcode == D_ACCESS_ACK_DATA),(io_up_d_payload_opcode == D_ACCESS_ACK)}}}));
  always @(*) begin
    a_halted_ready = 1'b1;
    if(when_Stream_l1084) begin
      a_halted_ready = 1'b0;
    end
    if(when_Stream_l1084_1) begin
      a_halted_ready = 1'b0;
    end
  end

  assign when_Stream_l1084 = ((! a_cmdFork_ready) && a_halted_fork2_logic_linkEnable_0);
  assign when_Stream_l1084_1 = ((! a_dataFork_ready) && a_halted_fork2_logic_linkEnable_1);
  assign a_cmdFork_valid = (a_halted_valid && a_halted_fork2_logic_linkEnable_0);
  assign a_cmdFork_payload_opcode = a_halted_payload_opcode;
  assign a_cmdFork_payload_param = a_halted_payload_param;
  assign a_cmdFork_payload_source = a_halted_payload_source;
  assign a_cmdFork_payload_address = a_halted_payload_address;
  assign a_cmdFork_payload_size = a_halted_payload_size;
  assign a_cmdFork_payload_mask = a_halted_payload_mask;
  assign a_cmdFork_payload_data = a_halted_payload_data;
  assign a_cmdFork_payload_corrupt = a_halted_payload_corrupt;
  assign a_cmdFork_fire = (a_cmdFork_valid && a_cmdFork_ready);
  assign a_dataFork_valid = (a_halted_valid && a_halted_fork2_logic_linkEnable_1);
  assign a_dataFork_payload_opcode = a_halted_payload_opcode;
  assign a_dataFork_payload_param = a_halted_payload_param;
  assign a_dataFork_payload_source = a_halted_payload_source;
  assign a_dataFork_payload_address = a_halted_payload_address;
  assign a_dataFork_payload_size = a_halted_payload_size;
  assign a_dataFork_payload_mask = a_halted_payload_mask;
  assign a_dataFork_payload_data = a_halted_payload_data;
  assign a_dataFork_payload_corrupt = a_halted_payload_corrupt;
  assign a_dataFork_fire = (a_dataFork_valid && a_dataFork_ready);
  assign a_cmdFork_tracker_last = ((! ((1'b0 || (A_PUT_FULL_DATA == a_cmdFork_payload_opcode)) || (A_PUT_PARTIAL_DATA == a_cmdFork_payload_opcode))) || (a_cmdFork_tracker_beat == _zz_a_cmdFork_tracker_last));
  assign when_Stream_l466 = (! (a_cmdFork_tracker_beat == 3'b000));
  always @(*) begin
    a_cmd_filtred_valid = a_cmdFork_valid;
    if(when_Stream_l466) begin
      a_cmd_filtred_valid = 1'b0;
    end
  end

  always @(*) begin
    a_cmdFork_ready = a_cmd_filtred_ready;
    if(when_Stream_l466) begin
      a_cmdFork_ready = 1'b1;
    end
  end

  assign a_cmd_filtred_payload_opcode = a_cmdFork_payload_opcode;
  assign a_cmd_filtred_payload_param = a_cmdFork_payload_param;
  assign a_cmd_filtred_payload_source = a_cmdFork_payload_source;
  assign a_cmd_filtred_payload_address = a_cmdFork_payload_address;
  assign a_cmd_filtred_payload_size = a_cmdFork_payload_size;
  assign a_cmd_filtred_payload_mask = a_cmdFork_payload_mask;
  assign a_cmd_filtred_payload_data = a_cmdFork_payload_data;
  assign a_cmd_filtred_payload_corrupt = a_cmdFork_payload_corrupt;
  assign a_cmd_buffered_fire = (a_cmd_buffered_valid && a_cmd_buffered_ready);
  assign a_cmd_filtred_ready = (! a_cmd_filtred_rValid);
  assign a_cmd_buffered_valid = a_cmd_filtred_rValid;
  assign a_cmd_buffered_payload_opcode = a_cmd_filtred_rData_opcode;
  assign a_cmd_buffered_payload_param = a_cmd_filtred_rData_param;
  assign a_cmd_buffered_payload_source = a_cmd_filtred_rData_source;
  assign a_cmd_buffered_payload_address = a_cmd_filtred_rData_address;
  assign a_cmd_buffered_payload_size = a_cmd_filtred_rData_size;
  assign a_cmd_buffered_payload_mask = a_cmd_filtred_rData_mask;
  assign a_cmd_buffered_payload_data = a_cmd_filtred_rData_data;
  assign a_cmd_buffered_payload_corrupt = a_cmd_filtred_rData_corrupt;
  assign a_cmd_isGet = (a_cmd_buffered_payload_opcode == A_GET);
  assign io_down_aw_valid = (a_cmd_buffered_valid && (! a_cmd_isGet));
  assign io_down_ar_valid = (a_cmd_buffered_valid && a_cmd_isGet);
  assign a_cmd_buffered_ready = (a_cmd_isGet ? io_down_ar_ready : io_down_aw_ready);
  assign a_cmd_len = {5'd0, _zz_a_cmd_len};
  assign a_cmd_sizePerBeat = _zz_a_cmd_sizePerBeat;
  assign io_down_aw_payload_addr = a_cmd_buffered_payload_address;
  assign io_down_aw_payload_id = a_cmd_buffered_payload_source;
  assign io_down_aw_payload_len = a_cmd_len;
  assign io_down_aw_payload_size = a_cmd_sizePerBeat;
  assign io_down_aw_payload_burst = 2'b01;
  assign io_down_ar_payload_addr = a_cmd_buffered_payload_address;
  assign io_down_ar_payload_id = a_cmd_buffered_payload_source;
  assign io_down_ar_payload_len = a_cmd_len;
  assign io_down_ar_payload_size = a_cmd_sizePerBeat;
  assign io_down_ar_payload_burst = 2'b01;
  assign io_down_aw_payload_allStrb = (a_cmd_buffered_payload_opcode == A_PUT_FULL_DATA);
  assign when_Stream_l466_1 = (! ((a_dataFork_payload_opcode == A_PUT_FULL_DATA) || (a_dataFork_payload_opcode == A_PUT_PARTIAL_DATA)));
  always @(*) begin
    a_data_filtred_valid = a_dataFork_valid;
    if(when_Stream_l466_1) begin
      a_data_filtred_valid = 1'b0;
    end
  end

  always @(*) begin
    a_dataFork_ready = a_data_filtred_ready;
    if(when_Stream_l466_1) begin
      a_dataFork_ready = 1'b1;
    end
  end

  assign a_data_filtred_payload_opcode = a_dataFork_payload_opcode;
  assign a_data_filtred_payload_param = a_dataFork_payload_param;
  assign a_data_filtred_payload_source = a_dataFork_payload_source;
  assign a_data_filtred_payload_address = a_dataFork_payload_address;
  assign a_data_filtred_payload_size = a_dataFork_payload_size;
  assign a_data_filtred_payload_mask = a_dataFork_payload_mask;
  assign a_data_filtred_payload_data = a_dataFork_payload_data;
  assign a_data_filtred_payload_corrupt = a_dataFork_payload_corrupt;
  always @(*) begin
    a_data_filtred_ready = a_data_buffer_ready;
    if(when_Stream_l393) begin
      a_data_filtred_ready = 1'b1;
    end
  end

  assign when_Stream_l393 = (! a_data_buffer_valid);
  assign a_data_buffer_valid = a_data_filtred_rValid;
  assign a_data_buffer_payload_opcode = a_data_filtred_rData_opcode;
  assign a_data_buffer_payload_param = a_data_filtred_rData_param;
  assign a_data_buffer_payload_source = a_data_filtred_rData_source;
  assign a_data_buffer_payload_address = a_data_filtred_rData_address;
  assign a_data_buffer_payload_size = a_data_filtred_rData_size;
  assign a_data_buffer_payload_mask = a_data_filtred_rData_mask;
  assign a_data_buffer_payload_data = a_data_filtred_rData_data;
  assign a_data_buffer_payload_corrupt = a_data_filtred_rData_corrupt;
  assign io_down_w_valid = a_data_buffer_valid;
  assign a_data_buffer_ready = io_down_w_ready;
  assign io_down_w_payload_data = a_data_buffer_payload_data;
  assign io_down_w_payload_strb = a_data_buffer_payload_mask;
  assign a_data_buffer_tracker_last = ((! ((1'b0 || (A_PUT_FULL_DATA == a_data_buffer_payload_opcode)) || (A_PUT_PARTIAL_DATA == a_data_buffer_payload_opcode))) || (a_data_buffer_tracker_beat == _zz_a_data_buffer_tracker_last));
  assign a_data_buffer_fire = (a_data_buffer_valid && a_data_buffer_ready);
  assign io_down_w_payload_last = a_data_buffer_tracker_last;
  assign io_down_b_ready = d_arbiter_io_inputs_0_ready;
  assign d_arbiter_io_inputs_0_payload_denied = (! (io_down_b_payload_resp == 2'b00));
  assign io_down_r_ready = d_arbiter_io_inputs_1_ready;
  assign d_arbiter_io_inputs_1_payload_denied = (! (io_down_r_payload_resp == 2'b00));
  assign io_up_d_valid = d_arbiter_io_output_valid;
  assign _zz_io_up_d_payload_opcode = (d_arbiter_io_chosen[0] ? D_ACCESS_ACK_DATA : D_ACCESS_ACK);
  assign io_up_d_payload_opcode = _zz_io_up_d_payload_opcode;
  assign io_up_d_payload_param = 3'b000;
  assign io_up_d_payload_source = d_arbiter_io_output_payload_source;
  assign io_up_d_payload_denied = d_arbiter_io_output_payload_denied;
  assign io_up_d_payload_data = io_down_r_payload_data;
  assign io_up_d_payload_corrupt = 1'b0;
  assign io_up_d_payload_size = a_ctx_io_query_context;
  always @(posedge clk_cpu or posedge reset_cpu) begin
    if(reset_cpu) begin
      io_up_a_tracker_beat <= 3'b000;
      io_up_d_tracker_beat <= 3'b000;
      a_halted_fork2_logic_linkEnable_0 <= 1'b1;
      a_halted_fork2_logic_linkEnable_1 <= 1'b1;
      a_cmdFork_tracker_beat <= 3'b000;
      a_cmd_filtred_rValid <= 1'b0;
      a_data_filtred_rValid <= 1'b0;
      a_data_buffer_tracker_beat <= 3'b000;
    end else begin
      if(io_up_a_fire) begin
        io_up_a_tracker_beat <= (io_up_a_tracker_beat + 3'b001);
        if(io_up_a_tracker_last) begin
          io_up_a_tracker_beat <= 3'b000;
        end
      end
      if(io_up_d_fire) begin
        io_up_d_tracker_beat <= (io_up_d_tracker_beat + 3'b001);
        if(io_up_d_tracker_last) begin
          io_up_d_tracker_beat <= 3'b000;
        end
      end
      if(a_cmdFork_fire) begin
        a_halted_fork2_logic_linkEnable_0 <= 1'b0;
      end
      if(a_dataFork_fire) begin
        a_halted_fork2_logic_linkEnable_1 <= 1'b0;
      end
      if(a_halted_ready) begin
        a_halted_fork2_logic_linkEnable_0 <= 1'b1;
        a_halted_fork2_logic_linkEnable_1 <= 1'b1;
      end
      if(a_cmdFork_fire) begin
        a_cmdFork_tracker_beat <= (a_cmdFork_tracker_beat + 3'b001);
        if(a_cmdFork_tracker_last) begin
          a_cmdFork_tracker_beat <= 3'b000;
        end
      end
      if(a_cmd_filtred_valid) begin
        a_cmd_filtred_rValid <= 1'b1;
      end
      if(a_cmd_buffered_fire) begin
        a_cmd_filtred_rValid <= 1'b0;
      end
      if(a_data_filtred_ready) begin
        a_data_filtred_rValid <= a_data_filtred_valid;
      end
      if(a_data_buffer_fire) begin
        a_data_buffer_tracker_beat <= (a_data_buffer_tracker_beat + 3'b001);
        if(a_data_buffer_tracker_last) begin
          a_data_buffer_tracker_beat <= 3'b000;
        end
      end
    end
  end

  always @(posedge clk_cpu) begin
    if(a_cmd_filtred_ready) begin
      a_cmd_filtred_rData_opcode <= a_cmd_filtred_payload_opcode;
      a_cmd_filtred_rData_param <= a_cmd_filtred_payload_param;
      a_cmd_filtred_rData_source <= a_cmd_filtred_payload_source;
      a_cmd_filtred_rData_address <= a_cmd_filtred_payload_address;
      a_cmd_filtred_rData_size <= a_cmd_filtred_payload_size;
      a_cmd_filtred_rData_mask <= a_cmd_filtred_payload_mask;
      a_cmd_filtred_rData_data <= a_cmd_filtred_payload_data;
      a_cmd_filtred_rData_corrupt <= a_cmd_filtred_payload_corrupt;
    end
    if(a_data_filtred_ready) begin
      a_data_filtred_rData_opcode <= a_data_filtred_payload_opcode;
      a_data_filtred_rData_param <= a_data_filtred_payload_param;
      a_data_filtred_rData_source <= a_data_filtred_payload_source;
      a_data_filtred_rData_address <= a_data_filtred_payload_address;
      a_data_filtred_rData_size <= a_data_filtred_payload_size;
      a_data_filtred_rData_mask <= a_data_filtred_payload_mask;
      a_data_filtred_rData_data <= a_data_filtred_payload_data;
      a_data_filtred_rData_corrupt <= a_data_filtred_payload_corrupt;
    end
  end


endmodule

module Arbiter (
  input  wire          io_ups_0_a_valid,
  output wire          io_ups_0_a_ready,
  input  wire [2:0]    io_ups_0_a_payload_opcode,
  input  wire [2:0]    io_ups_0_a_payload_param,
  input  wire [31:0]   io_ups_0_a_payload_address,
  input  wire [2:0]    io_ups_0_a_payload_size,
  output wire          io_ups_0_d_valid,
  input  wire          io_ups_0_d_ready,
  output wire [2:0]    io_ups_0_d_payload_opcode,
  output wire [2:0]    io_ups_0_d_payload_param,
  output wire [2:0]    io_ups_0_d_payload_size,
  output wire          io_ups_0_d_payload_denied,
  output wire [63:0]   io_ups_0_d_payload_data,
  output wire          io_ups_0_d_payload_corrupt,
  input  wire          io_ups_1_a_valid,
  output wire          io_ups_1_a_ready,
  input  wire [2:0]    io_ups_1_a_payload_opcode,
  input  wire [2:0]    io_ups_1_a_payload_param,
  input  wire [31:0]   io_ups_1_a_payload_address,
  input  wire [1:0]    io_ups_1_a_payload_size,
  input  wire [7:0]    io_ups_1_a_payload_mask,
  input  wire [63:0]   io_ups_1_a_payload_data,
  input  wire          io_ups_1_a_payload_corrupt,
  output wire          io_ups_1_d_valid,
  input  wire          io_ups_1_d_ready,
  output wire [2:0]    io_ups_1_d_payload_opcode,
  output wire [2:0]    io_ups_1_d_payload_param,
  output wire [1:0]    io_ups_1_d_payload_size,
  output wire          io_ups_1_d_payload_denied,
  output wire [63:0]   io_ups_1_d_payload_data,
  output wire          io_ups_1_d_payload_corrupt,
  input  wire          io_ups_2_a_valid,
  output wire          io_ups_2_a_ready,
  input  wire [2:0]    io_ups_2_a_payload_opcode,
  input  wire [2:0]    io_ups_2_a_payload_param,
  input  wire [0:0]    io_ups_2_a_payload_source,
  input  wire [31:0]   io_ups_2_a_payload_address,
  input  wire [2:0]    io_ups_2_a_payload_size,
  input  wire [7:0]    io_ups_2_a_payload_mask,
  input  wire [63:0]   io_ups_2_a_payload_data,
  input  wire          io_ups_2_a_payload_corrupt,
  output wire          io_ups_2_d_valid,
  input  wire          io_ups_2_d_ready,
  output wire [2:0]    io_ups_2_d_payload_opcode,
  output wire [2:0]    io_ups_2_d_payload_param,
  output wire [0:0]    io_ups_2_d_payload_source,
  output wire [2:0]    io_ups_2_d_payload_size,
  output wire          io_ups_2_d_payload_denied,
  output wire [63:0]   io_ups_2_d_payload_data,
  output wire          io_ups_2_d_payload_corrupt,
  output wire          io_down_a_valid,
  input  wire          io_down_a_ready,
  output wire [2:0]    io_down_a_payload_opcode,
  output wire [2:0]    io_down_a_payload_param,
  output wire [2:0]    io_down_a_payload_source,
  output wire [31:0]   io_down_a_payload_address,
  output wire [2:0]    io_down_a_payload_size,
  output wire [7:0]    io_down_a_payload_mask,
  output wire [63:0]   io_down_a_payload_data,
  output wire          io_down_a_payload_corrupt,
  input  wire          io_down_d_valid,
  output wire          io_down_d_ready,
  input  wire [2:0]    io_down_d_payload_opcode,
  input  wire [2:0]    io_down_d_payload_param,
  input  wire [2:0]    io_down_d_payload_source,
  input  wire [2:0]    io_down_d_payload_size,
  input  wire          io_down_d_payload_denied,
  input  wire [63:0]   io_down_d_payload_data,
  input  wire          io_down_d_payload_corrupt,
  input  wire          clk_cpu,
  input  wire          reset_cpu
);
  localparam A_PUT_FULL_DATA = 3'd0;
  localparam A_PUT_PARTIAL_DATA = 3'd1;
  localparam A_GET = 3'd4;
  localparam A_ACQUIRE_BLOCK = 3'd6;
  localparam A_ACQUIRE_PERM = 3'd7;
  localparam D_ACCESS_ACK = 3'd0;
  localparam D_ACCESS_ACK_DATA = 3'd1;
  localparam D_GRANT = 3'd4;
  localparam D_GRANT_DATA = 3'd5;
  localparam D_RELEASE_ACK = 3'd6;

  wire       [2:0]    a_arbiter_io_inputs_1_payload_size;
  wire                a_arbiter_io_inputs_0_ready;
  wire                a_arbiter_io_inputs_1_ready;
  wire                a_arbiter_io_inputs_2_ready;
  wire                a_arbiter_io_output_valid;
  wire       [2:0]    a_arbiter_io_output_payload_opcode;
  wire       [2:0]    a_arbiter_io_output_payload_param;
  wire       [2:0]    a_arbiter_io_output_payload_source;
  wire       [31:0]   a_arbiter_io_output_payload_address;
  wire       [2:0]    a_arbiter_io_output_payload_size;
  wire       [7:0]    a_arbiter_io_output_payload_mask;
  wire       [63:0]   a_arbiter_io_output_payload_data;
  wire                a_arbiter_io_output_payload_corrupt;
  wire       [1:0]    a_arbiter_io_chosen;
  wire       [2:0]    a_arbiter_io_chosenOH;
  wire       [2:0]    _zz_ups_2_a_payload_source;
  reg                 _zz_io_down_d_ready;
  wire                ups_0_a_valid;
  wire                ups_0_a_ready;
  wire       [2:0]    ups_0_a_payload_opcode;
  wire       [2:0]    ups_0_a_payload_param;
  wire       [2:0]    ups_0_a_payload_source;
  wire       [31:0]   ups_0_a_payload_address;
  wire       [2:0]    ups_0_a_payload_size;
  wire                ups_0_d_valid;
  wire                ups_0_d_ready;
  wire       [2:0]    ups_0_d_payload_opcode;
  wire       [2:0]    ups_0_d_payload_param;
  wire       [2:0]    ups_0_d_payload_source;
  wire       [2:0]    ups_0_d_payload_size;
  wire                ups_0_d_payload_denied;
  wire       [63:0]   ups_0_d_payload_data;
  wire                ups_0_d_payload_corrupt;
  wire                ups_1_a_valid;
  wire                ups_1_a_ready;
  wire       [2:0]    ups_1_a_payload_opcode;
  wire       [2:0]    ups_1_a_payload_param;
  wire       [2:0]    ups_1_a_payload_source;
  wire       [31:0]   ups_1_a_payload_address;
  wire       [1:0]    ups_1_a_payload_size;
  wire       [7:0]    ups_1_a_payload_mask;
  wire       [63:0]   ups_1_a_payload_data;
  wire                ups_1_a_payload_corrupt;
  wire                ups_1_d_valid;
  wire                ups_1_d_ready;
  wire       [2:0]    ups_1_d_payload_opcode;
  wire       [2:0]    ups_1_d_payload_param;
  wire       [2:0]    ups_1_d_payload_source;
  wire       [1:0]    ups_1_d_payload_size;
  wire                ups_1_d_payload_denied;
  wire       [63:0]   ups_1_d_payload_data;
  wire                ups_1_d_payload_corrupt;
  wire                ups_2_a_valid;
  wire                ups_2_a_ready;
  wire       [2:0]    ups_2_a_payload_opcode;
  wire       [2:0]    ups_2_a_payload_param;
  wire       [2:0]    ups_2_a_payload_source;
  wire       [31:0]   ups_2_a_payload_address;
  wire       [2:0]    ups_2_a_payload_size;
  wire       [7:0]    ups_2_a_payload_mask;
  wire       [63:0]   ups_2_a_payload_data;
  wire                ups_2_a_payload_corrupt;
  wire                ups_2_d_valid;
  wire                ups_2_d_ready;
  wire       [2:0]    ups_2_d_payload_opcode;
  wire       [2:0]    ups_2_d_payload_param;
  wire       [2:0]    ups_2_d_payload_source;
  wire       [2:0]    ups_2_d_payload_size;
  wire                ups_2_d_payload_denied;
  wire       [63:0]   ups_2_d_payload_data;
  wire                ups_2_d_payload_corrupt;
  wire       [1:0]    d_sel;
  `ifndef SYNTHESIS
  reg [127:0] io_ups_0_a_payload_opcode_string;
  reg [119:0] io_ups_0_d_payload_opcode_string;
  reg [127:0] io_ups_1_a_payload_opcode_string;
  reg [119:0] io_ups_1_d_payload_opcode_string;
  reg [127:0] io_ups_2_a_payload_opcode_string;
  reg [119:0] io_ups_2_d_payload_opcode_string;
  reg [127:0] io_down_a_payload_opcode_string;
  reg [119:0] io_down_d_payload_opcode_string;
  reg [127:0] ups_0_a_payload_opcode_string;
  reg [119:0] ups_0_d_payload_opcode_string;
  reg [127:0] ups_1_a_payload_opcode_string;
  reg [119:0] ups_1_d_payload_opcode_string;
  reg [127:0] ups_2_a_payload_opcode_string;
  reg [119:0] ups_2_d_payload_opcode_string;
  `endif


  assign _zz_ups_2_a_payload_source = {2'd0, io_ups_2_a_payload_source};
  StreamArbiter_5 a_arbiter (
    .io_inputs_0_valid           (ups_0_a_valid                                                       ), //i
    .io_inputs_0_ready           (a_arbiter_io_inputs_0_ready                                         ), //o
    .io_inputs_0_payload_opcode  (ups_0_a_payload_opcode[2:0]                                         ), //i
    .io_inputs_0_payload_param   (ups_0_a_payload_param[2:0]                                          ), //i
    .io_inputs_0_payload_source  (ups_0_a_payload_source[2:0]                                         ), //i
    .io_inputs_0_payload_address (ups_0_a_payload_address[31:0]                                       ), //i
    .io_inputs_0_payload_size    (ups_0_a_payload_size[2:0]                                           ), //i
    .io_inputs_0_payload_mask    (8'bxxxxxxxx                                                         ), //i
    .io_inputs_0_payload_data    (64'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx), //i
    .io_inputs_0_payload_corrupt (1'b0                                                                ), //i
    .io_inputs_1_valid           (ups_1_a_valid                                                       ), //i
    .io_inputs_1_ready           (a_arbiter_io_inputs_1_ready                                         ), //o
    .io_inputs_1_payload_opcode  (ups_1_a_payload_opcode[2:0]                                         ), //i
    .io_inputs_1_payload_param   (ups_1_a_payload_param[2:0]                                          ), //i
    .io_inputs_1_payload_source  (ups_1_a_payload_source[2:0]                                         ), //i
    .io_inputs_1_payload_address (ups_1_a_payload_address[31:0]                                       ), //i
    .io_inputs_1_payload_size    (a_arbiter_io_inputs_1_payload_size[2:0]                             ), //i
    .io_inputs_1_payload_mask    (ups_1_a_payload_mask[7:0]                                           ), //i
    .io_inputs_1_payload_data    (ups_1_a_payload_data[63:0]                                          ), //i
    .io_inputs_1_payload_corrupt (ups_1_a_payload_corrupt                                             ), //i
    .io_inputs_2_valid           (ups_2_a_valid                                                       ), //i
    .io_inputs_2_ready           (a_arbiter_io_inputs_2_ready                                         ), //o
    .io_inputs_2_payload_opcode  (ups_2_a_payload_opcode[2:0]                                         ), //i
    .io_inputs_2_payload_param   (ups_2_a_payload_param[2:0]                                          ), //i
    .io_inputs_2_payload_source  (ups_2_a_payload_source[2:0]                                         ), //i
    .io_inputs_2_payload_address (ups_2_a_payload_address[31:0]                                       ), //i
    .io_inputs_2_payload_size    (ups_2_a_payload_size[2:0]                                           ), //i
    .io_inputs_2_payload_mask    (ups_2_a_payload_mask[7:0]                                           ), //i
    .io_inputs_2_payload_data    (ups_2_a_payload_data[63:0]                                          ), //i
    .io_inputs_2_payload_corrupt (ups_2_a_payload_corrupt                                             ), //i
    .io_output_valid             (a_arbiter_io_output_valid                                           ), //o
    .io_output_ready             (io_down_a_ready                                                     ), //i
    .io_output_payload_opcode    (a_arbiter_io_output_payload_opcode[2:0]                             ), //o
    .io_output_payload_param     (a_arbiter_io_output_payload_param[2:0]                              ), //o
    .io_output_payload_source    (a_arbiter_io_output_payload_source[2:0]                             ), //o
    .io_output_payload_address   (a_arbiter_io_output_payload_address[31:0]                           ), //o
    .io_output_payload_size      (a_arbiter_io_output_payload_size[2:0]                               ), //o
    .io_output_payload_mask      (a_arbiter_io_output_payload_mask[7:0]                               ), //o
    .io_output_payload_data      (a_arbiter_io_output_payload_data[63:0]                              ), //o
    .io_output_payload_corrupt   (a_arbiter_io_output_payload_corrupt                                 ), //o
    .io_chosen                   (a_arbiter_io_chosen[1:0]                                            ), //o
    .io_chosenOH                 (a_arbiter_io_chosenOH[2:0]                                          ), //o
    .clk_cpu                     (clk_cpu                                                             ), //i
    .reset_cpu                   (reset_cpu                                                           )  //i
  );
  always @(*) begin
    case(d_sel)
      2'b00 : _zz_io_down_d_ready = ups_0_d_ready;
      2'b01 : _zz_io_down_d_ready = ups_1_d_ready;
      default : _zz_io_down_d_ready = ups_2_d_ready;
    endcase
  end

  `ifndef SYNTHESIS
  always @(*) begin
    case(io_ups_0_a_payload_opcode)
      A_PUT_FULL_DATA : io_ups_0_a_payload_opcode_string = "PUT_FULL_DATA   ";
      A_PUT_PARTIAL_DATA : io_ups_0_a_payload_opcode_string = "PUT_PARTIAL_DATA";
      A_GET : io_ups_0_a_payload_opcode_string = "GET             ";
      A_ACQUIRE_BLOCK : io_ups_0_a_payload_opcode_string = "ACQUIRE_BLOCK   ";
      A_ACQUIRE_PERM : io_ups_0_a_payload_opcode_string = "ACQUIRE_PERM    ";
      default : io_ups_0_a_payload_opcode_string = "????????????????";
    endcase
  end
  always @(*) begin
    case(io_ups_0_d_payload_opcode)
      D_ACCESS_ACK : io_ups_0_d_payload_opcode_string = "ACCESS_ACK     ";
      D_ACCESS_ACK_DATA : io_ups_0_d_payload_opcode_string = "ACCESS_ACK_DATA";
      D_GRANT : io_ups_0_d_payload_opcode_string = "GRANT          ";
      D_GRANT_DATA : io_ups_0_d_payload_opcode_string = "GRANT_DATA     ";
      D_RELEASE_ACK : io_ups_0_d_payload_opcode_string = "RELEASE_ACK    ";
      default : io_ups_0_d_payload_opcode_string = "???????????????";
    endcase
  end
  always @(*) begin
    case(io_ups_1_a_payload_opcode)
      A_PUT_FULL_DATA : io_ups_1_a_payload_opcode_string = "PUT_FULL_DATA   ";
      A_PUT_PARTIAL_DATA : io_ups_1_a_payload_opcode_string = "PUT_PARTIAL_DATA";
      A_GET : io_ups_1_a_payload_opcode_string = "GET             ";
      A_ACQUIRE_BLOCK : io_ups_1_a_payload_opcode_string = "ACQUIRE_BLOCK   ";
      A_ACQUIRE_PERM : io_ups_1_a_payload_opcode_string = "ACQUIRE_PERM    ";
      default : io_ups_1_a_payload_opcode_string = "????????????????";
    endcase
  end
  always @(*) begin
    case(io_ups_1_d_payload_opcode)
      D_ACCESS_ACK : io_ups_1_d_payload_opcode_string = "ACCESS_ACK     ";
      D_ACCESS_ACK_DATA : io_ups_1_d_payload_opcode_string = "ACCESS_ACK_DATA";
      D_GRANT : io_ups_1_d_payload_opcode_string = "GRANT          ";
      D_GRANT_DATA : io_ups_1_d_payload_opcode_string = "GRANT_DATA     ";
      D_RELEASE_ACK : io_ups_1_d_payload_opcode_string = "RELEASE_ACK    ";
      default : io_ups_1_d_payload_opcode_string = "???????????????";
    endcase
  end
  always @(*) begin
    case(io_ups_2_a_payload_opcode)
      A_PUT_FULL_DATA : io_ups_2_a_payload_opcode_string = "PUT_FULL_DATA   ";
      A_PUT_PARTIAL_DATA : io_ups_2_a_payload_opcode_string = "PUT_PARTIAL_DATA";
      A_GET : io_ups_2_a_payload_opcode_string = "GET             ";
      A_ACQUIRE_BLOCK : io_ups_2_a_payload_opcode_string = "ACQUIRE_BLOCK   ";
      A_ACQUIRE_PERM : io_ups_2_a_payload_opcode_string = "ACQUIRE_PERM    ";
      default : io_ups_2_a_payload_opcode_string = "????????????????";
    endcase
  end
  always @(*) begin
    case(io_ups_2_d_payload_opcode)
      D_ACCESS_ACK : io_ups_2_d_payload_opcode_string = "ACCESS_ACK     ";
      D_ACCESS_ACK_DATA : io_ups_2_d_payload_opcode_string = "ACCESS_ACK_DATA";
      D_GRANT : io_ups_2_d_payload_opcode_string = "GRANT          ";
      D_GRANT_DATA : io_ups_2_d_payload_opcode_string = "GRANT_DATA     ";
      D_RELEASE_ACK : io_ups_2_d_payload_opcode_string = "RELEASE_ACK    ";
      default : io_ups_2_d_payload_opcode_string = "???????????????";
    endcase
  end
  always @(*) begin
    case(io_down_a_payload_opcode)
      A_PUT_FULL_DATA : io_down_a_payload_opcode_string = "PUT_FULL_DATA   ";
      A_PUT_PARTIAL_DATA : io_down_a_payload_opcode_string = "PUT_PARTIAL_DATA";
      A_GET : io_down_a_payload_opcode_string = "GET             ";
      A_ACQUIRE_BLOCK : io_down_a_payload_opcode_string = "ACQUIRE_BLOCK   ";
      A_ACQUIRE_PERM : io_down_a_payload_opcode_string = "ACQUIRE_PERM    ";
      default : io_down_a_payload_opcode_string = "????????????????";
    endcase
  end
  always @(*) begin
    case(io_down_d_payload_opcode)
      D_ACCESS_ACK : io_down_d_payload_opcode_string = "ACCESS_ACK     ";
      D_ACCESS_ACK_DATA : io_down_d_payload_opcode_string = "ACCESS_ACK_DATA";
      D_GRANT : io_down_d_payload_opcode_string = "GRANT          ";
      D_GRANT_DATA : io_down_d_payload_opcode_string = "GRANT_DATA     ";
      D_RELEASE_ACK : io_down_d_payload_opcode_string = "RELEASE_ACK    ";
      default : io_down_d_payload_opcode_string = "???????????????";
    endcase
  end
  always @(*) begin
    case(ups_0_a_payload_opcode)
      A_PUT_FULL_DATA : ups_0_a_payload_opcode_string = "PUT_FULL_DATA   ";
      A_PUT_PARTIAL_DATA : ups_0_a_payload_opcode_string = "PUT_PARTIAL_DATA";
      A_GET : ups_0_a_payload_opcode_string = "GET             ";
      A_ACQUIRE_BLOCK : ups_0_a_payload_opcode_string = "ACQUIRE_BLOCK   ";
      A_ACQUIRE_PERM : ups_0_a_payload_opcode_string = "ACQUIRE_PERM    ";
      default : ups_0_a_payload_opcode_string = "????????????????";
    endcase
  end
  always @(*) begin
    case(ups_0_d_payload_opcode)
      D_ACCESS_ACK : ups_0_d_payload_opcode_string = "ACCESS_ACK     ";
      D_ACCESS_ACK_DATA : ups_0_d_payload_opcode_string = "ACCESS_ACK_DATA";
      D_GRANT : ups_0_d_payload_opcode_string = "GRANT          ";
      D_GRANT_DATA : ups_0_d_payload_opcode_string = "GRANT_DATA     ";
      D_RELEASE_ACK : ups_0_d_payload_opcode_string = "RELEASE_ACK    ";
      default : ups_0_d_payload_opcode_string = "???????????????";
    endcase
  end
  always @(*) begin
    case(ups_1_a_payload_opcode)
      A_PUT_FULL_DATA : ups_1_a_payload_opcode_string = "PUT_FULL_DATA   ";
      A_PUT_PARTIAL_DATA : ups_1_a_payload_opcode_string = "PUT_PARTIAL_DATA";
      A_GET : ups_1_a_payload_opcode_string = "GET             ";
      A_ACQUIRE_BLOCK : ups_1_a_payload_opcode_string = "ACQUIRE_BLOCK   ";
      A_ACQUIRE_PERM : ups_1_a_payload_opcode_string = "ACQUIRE_PERM    ";
      default : ups_1_a_payload_opcode_string = "????????????????";
    endcase
  end
  always @(*) begin
    case(ups_1_d_payload_opcode)
      D_ACCESS_ACK : ups_1_d_payload_opcode_string = "ACCESS_ACK     ";
      D_ACCESS_ACK_DATA : ups_1_d_payload_opcode_string = "ACCESS_ACK_DATA";
      D_GRANT : ups_1_d_payload_opcode_string = "GRANT          ";
      D_GRANT_DATA : ups_1_d_payload_opcode_string = "GRANT_DATA     ";
      D_RELEASE_ACK : ups_1_d_payload_opcode_string = "RELEASE_ACK    ";
      default : ups_1_d_payload_opcode_string = "???????????????";
    endcase
  end
  always @(*) begin
    case(ups_2_a_payload_opcode)
      A_PUT_FULL_DATA : ups_2_a_payload_opcode_string = "PUT_FULL_DATA   ";
      A_PUT_PARTIAL_DATA : ups_2_a_payload_opcode_string = "PUT_PARTIAL_DATA";
      A_GET : ups_2_a_payload_opcode_string = "GET             ";
      A_ACQUIRE_BLOCK : ups_2_a_payload_opcode_string = "ACQUIRE_BLOCK   ";
      A_ACQUIRE_PERM : ups_2_a_payload_opcode_string = "ACQUIRE_PERM    ";
      default : ups_2_a_payload_opcode_string = "????????????????";
    endcase
  end
  always @(*) begin
    case(ups_2_d_payload_opcode)
      D_ACCESS_ACK : ups_2_d_payload_opcode_string = "ACCESS_ACK     ";
      D_ACCESS_ACK_DATA : ups_2_d_payload_opcode_string = "ACCESS_ACK_DATA";
      D_GRANT : ups_2_d_payload_opcode_string = "GRANT          ";
      D_GRANT_DATA : ups_2_d_payload_opcode_string = "GRANT_DATA     ";
      D_RELEASE_ACK : ups_2_d_payload_opcode_string = "RELEASE_ACK    ";
      default : ups_2_d_payload_opcode_string = "???????????????";
    endcase
  end
  `endif

  assign ups_0_a_valid = io_ups_0_a_valid;
  assign io_ups_0_a_ready = ups_0_a_ready;
  assign ups_0_a_payload_opcode = io_ups_0_a_payload_opcode;
  assign ups_0_a_payload_param = io_ups_0_a_payload_param;
  assign ups_0_a_payload_address = io_ups_0_a_payload_address;
  assign ups_0_a_payload_size = io_ups_0_a_payload_size;
  assign io_ups_0_d_valid = ups_0_d_valid;
  assign ups_0_d_ready = io_ups_0_d_ready;
  assign io_ups_0_d_payload_opcode = ups_0_d_payload_opcode;
  assign io_ups_0_d_payload_param = ups_0_d_payload_param;
  assign io_ups_0_d_payload_size = ups_0_d_payload_size;
  assign io_ups_0_d_payload_denied = ups_0_d_payload_denied;
  assign io_ups_0_d_payload_data = ups_0_d_payload_data;
  assign io_ups_0_d_payload_corrupt = ups_0_d_payload_corrupt;
  assign ups_0_a_payload_source = (3'b000 | 3'b000);
  assign ups_1_a_valid = io_ups_1_a_valid;
  assign io_ups_1_a_ready = ups_1_a_ready;
  assign ups_1_a_payload_opcode = io_ups_1_a_payload_opcode;
  assign ups_1_a_payload_param = io_ups_1_a_payload_param;
  assign ups_1_a_payload_address = io_ups_1_a_payload_address;
  assign ups_1_a_payload_size = io_ups_1_a_payload_size;
  assign ups_1_a_payload_mask = io_ups_1_a_payload_mask;
  assign ups_1_a_payload_data = io_ups_1_a_payload_data;
  assign ups_1_a_payload_corrupt = io_ups_1_a_payload_corrupt;
  assign io_ups_1_d_valid = ups_1_d_valid;
  assign ups_1_d_ready = io_ups_1_d_ready;
  assign io_ups_1_d_payload_opcode = ups_1_d_payload_opcode;
  assign io_ups_1_d_payload_param = ups_1_d_payload_param;
  assign io_ups_1_d_payload_size = ups_1_d_payload_size;
  assign io_ups_1_d_payload_denied = ups_1_d_payload_denied;
  assign io_ups_1_d_payload_data = ups_1_d_payload_data;
  assign io_ups_1_d_payload_corrupt = ups_1_d_payload_corrupt;
  assign ups_1_a_payload_source = (3'b000 | 3'b010);
  assign ups_2_a_valid = io_ups_2_a_valid;
  assign io_ups_2_a_ready = ups_2_a_ready;
  assign ups_2_a_payload_opcode = io_ups_2_a_payload_opcode;
  assign ups_2_a_payload_param = io_ups_2_a_payload_param;
  assign ups_2_a_payload_address = io_ups_2_a_payload_address;
  assign ups_2_a_payload_size = io_ups_2_a_payload_size;
  assign ups_2_a_payload_mask = io_ups_2_a_payload_mask;
  assign ups_2_a_payload_data = io_ups_2_a_payload_data;
  assign ups_2_a_payload_corrupt = io_ups_2_a_payload_corrupt;
  assign io_ups_2_d_valid = ups_2_d_valid;
  assign ups_2_d_ready = io_ups_2_d_ready;
  assign io_ups_2_d_payload_opcode = ups_2_d_payload_opcode;
  assign io_ups_2_d_payload_param = ups_2_d_payload_param;
  assign io_ups_2_d_payload_size = ups_2_d_payload_size;
  assign io_ups_2_d_payload_denied = ups_2_d_payload_denied;
  assign io_ups_2_d_payload_data = ups_2_d_payload_data;
  assign io_ups_2_d_payload_corrupt = ups_2_d_payload_corrupt;
  assign ups_2_a_payload_source = (_zz_ups_2_a_payload_source | 3'b100);
  assign io_ups_2_d_payload_source = ups_2_d_payload_source[0:0];
  assign ups_0_a_ready = a_arbiter_io_inputs_0_ready;
  assign ups_1_a_ready = a_arbiter_io_inputs_1_ready;
  assign a_arbiter_io_inputs_1_payload_size = {1'd0, ups_1_a_payload_size};
  assign ups_2_a_ready = a_arbiter_io_inputs_2_ready;
  assign io_down_a_valid = a_arbiter_io_output_valid;
  assign io_down_a_payload_opcode = a_arbiter_io_output_payload_opcode;
  assign io_down_a_payload_param = a_arbiter_io_output_payload_param;
  assign io_down_a_payload_source = a_arbiter_io_output_payload_source;
  assign io_down_a_payload_address = a_arbiter_io_output_payload_address;
  assign io_down_a_payload_size = a_arbiter_io_output_payload_size;
  assign io_down_a_payload_mask = a_arbiter_io_output_payload_mask;
  assign io_down_a_payload_data = a_arbiter_io_output_payload_data;
  assign io_down_a_payload_corrupt = a_arbiter_io_output_payload_corrupt;
  assign d_sel = io_down_d_payload_source[2 : 1];
  assign io_down_d_ready = _zz_io_down_d_ready;
  assign ups_0_d_valid = (io_down_d_valid && (d_sel == 2'b00));
  assign ups_0_d_payload_opcode = io_down_d_payload_opcode;
  assign ups_0_d_payload_param = io_down_d_payload_param;
  assign ups_0_d_payload_source = io_down_d_payload_source;
  assign ups_0_d_payload_denied = io_down_d_payload_denied;
  assign ups_0_d_payload_size = io_down_d_payload_size;
  assign ups_0_d_payload_data = io_down_d_payload_data;
  assign ups_0_d_payload_corrupt = io_down_d_payload_corrupt;
  assign ups_1_d_valid = (io_down_d_valid && (d_sel == 2'b01));
  assign ups_1_d_payload_opcode = io_down_d_payload_opcode;
  assign ups_1_d_payload_param = io_down_d_payload_param;
  assign ups_1_d_payload_source = io_down_d_payload_source;
  assign ups_1_d_payload_denied = io_down_d_payload_denied;
  assign ups_1_d_payload_size = io_down_d_payload_size[1:0];
  assign ups_1_d_payload_data = io_down_d_payload_data;
  assign ups_1_d_payload_corrupt = io_down_d_payload_corrupt;
  assign ups_2_d_valid = (io_down_d_valid && (d_sel == 2'b10));
  assign ups_2_d_payload_opcode = io_down_d_payload_opcode;
  assign ups_2_d_payload_param = io_down_d_payload_param;
  assign ups_2_d_payload_source = io_down_d_payload_source;
  assign ups_2_d_payload_denied = io_down_d_payload_denied;
  assign ups_2_d_payload_size = io_down_d_payload_size;
  assign ups_2_d_payload_data = io_down_d_payload_data;
  assign ups_2_d_payload_corrupt = io_down_d_payload_corrupt;

endmodule

module VexiiRiscv (
  input  wire [63:0]   PrivilegedPlugin_logic_rdtime,
  input  wire          PrivilegedPlugin_logic_harts_0_int_m_timer /* verilator public */ ,
  input  wire          PrivilegedPlugin_logic_harts_0_int_m_software /* verilator public */ ,
  input  wire          PrivilegedPlugin_logic_harts_0_int_m_external /* verilator public */ ,
  input  wire          PrivilegedPlugin_logic_harts_0_int_s_external /* verilator public */ ,
  output wire          FetchL1TileLinkPlugin_logic_down_a_valid,
  input  wire          FetchL1TileLinkPlugin_logic_down_a_ready,
  output wire [2:0]    FetchL1TileLinkPlugin_logic_down_a_payload_opcode,
  output wire [2:0]    FetchL1TileLinkPlugin_logic_down_a_payload_param,
  output wire [31:0]   FetchL1TileLinkPlugin_logic_down_a_payload_address,
  output wire [2:0]    FetchL1TileLinkPlugin_logic_down_a_payload_size,
  input  wire          FetchL1TileLinkPlugin_logic_down_d_valid,
  output wire          FetchL1TileLinkPlugin_logic_down_d_ready,
  input  wire [2:0]    FetchL1TileLinkPlugin_logic_down_d_payload_opcode,
  input  wire [2:0]    FetchL1TileLinkPlugin_logic_down_d_payload_param,
  input  wire [2:0]    FetchL1TileLinkPlugin_logic_down_d_payload_size,
  input  wire          FetchL1TileLinkPlugin_logic_down_d_payload_denied,
  input  wire [63:0]   FetchL1TileLinkPlugin_logic_down_d_payload_data,
  input  wire          FetchL1TileLinkPlugin_logic_down_d_payload_corrupt,
  output reg           LsuL1TileLinkPlugin_logic_down_a_valid,
  input  wire          LsuL1TileLinkPlugin_logic_down_a_ready,
  output reg  [2:0]    LsuL1TileLinkPlugin_logic_down_a_payload_opcode,
  output wire [2:0]    LsuL1TileLinkPlugin_logic_down_a_payload_param,
  output reg  [0:0]    LsuL1TileLinkPlugin_logic_down_a_payload_source,
  output reg  [31:0]   LsuL1TileLinkPlugin_logic_down_a_payload_address,
  output wire [2:0]    LsuL1TileLinkPlugin_logic_down_a_payload_size,
  output wire [7:0]    LsuL1TileLinkPlugin_logic_down_a_payload_mask,
  output wire [63:0]   LsuL1TileLinkPlugin_logic_down_a_payload_data,
  output wire          LsuL1TileLinkPlugin_logic_down_a_payload_corrupt,
  input  wire          LsuL1TileLinkPlugin_logic_down_d_valid,
  output wire          LsuL1TileLinkPlugin_logic_down_d_ready,
  input  wire [2:0]    LsuL1TileLinkPlugin_logic_down_d_payload_opcode,
  input  wire [2:0]    LsuL1TileLinkPlugin_logic_down_d_payload_param,
  input  wire [0:0]    LsuL1TileLinkPlugin_logic_down_d_payload_source,
  input  wire [2:0]    LsuL1TileLinkPlugin_logic_down_d_payload_size,
  input  wire          LsuL1TileLinkPlugin_logic_down_d_payload_denied,
  input  wire [63:0]   LsuL1TileLinkPlugin_logic_down_d_payload_data,
  input  wire          LsuL1TileLinkPlugin_logic_down_d_payload_corrupt,
  output wire          LsuTileLinkPlugin_logic_bridge_down_a_valid,
  input  wire          LsuTileLinkPlugin_logic_bridge_down_a_ready,
  output wire [2:0]    LsuTileLinkPlugin_logic_bridge_down_a_payload_opcode,
  output wire [2:0]    LsuTileLinkPlugin_logic_bridge_down_a_payload_param,
  output wire [31:0]   LsuTileLinkPlugin_logic_bridge_down_a_payload_address,
  output wire [1:0]    LsuTileLinkPlugin_logic_bridge_down_a_payload_size,
  output wire [3:0]    LsuTileLinkPlugin_logic_bridge_down_a_payload_mask,
  output wire [31:0]   LsuTileLinkPlugin_logic_bridge_down_a_payload_data,
  output wire          LsuTileLinkPlugin_logic_bridge_down_a_payload_corrupt,
  input  wire          LsuTileLinkPlugin_logic_bridge_down_d_valid,
  output wire          LsuTileLinkPlugin_logic_bridge_down_d_ready,
  input  wire [2:0]    LsuTileLinkPlugin_logic_bridge_down_d_payload_opcode,
  input  wire [2:0]    LsuTileLinkPlugin_logic_bridge_down_d_payload_param,
  input  wire [1:0]    LsuTileLinkPlugin_logic_bridge_down_d_payload_size,
  input  wire          LsuTileLinkPlugin_logic_bridge_down_d_payload_denied,
  input  wire [31:0]   LsuTileLinkPlugin_logic_bridge_down_d_payload_data,
  input  wire          LsuTileLinkPlugin_logic_bridge_down_d_payload_corrupt,
  input  wire          clk_cpu,
  input  wire          reset_cpu
);
  localparam IntAluPlugin_AluBitwiseCtrlEnum_XOR_1 = 2'd0;
  localparam IntAluPlugin_AluBitwiseCtrlEnum_OR_1 = 2'd1;
  localparam IntAluPlugin_AluBitwiseCtrlEnum_AND_1 = 2'd2;
  localparam IntAluPlugin_AluBitwiseCtrlEnum_ZERO = 2'd3;
  localparam BranchPlugin_BranchCtrlEnum_B = 2'd0;
  localparam BranchPlugin_BranchCtrlEnum_JAL = 2'd1;
  localparam BranchPlugin_BranchCtrlEnum_JALR = 2'd2;
  localparam EnvPluginOp_ECALL = 3'd0;
  localparam EnvPluginOp_EBREAK = 3'd1;
  localparam EnvPluginOp_PRIV_RET = 3'd2;
  localparam EnvPluginOp_FENCE_I = 3'd3;
  localparam EnvPluginOp_SFENCE_VMA = 3'd4;
  localparam EnvPluginOp_WFI = 3'd5;
  localparam A_PUT_FULL_DATA = 3'd0;
  localparam A_PUT_PARTIAL_DATA = 3'd1;
  localparam A_GET = 3'd4;
  localparam A_ACQUIRE_BLOCK = 3'd6;
  localparam A_ACQUIRE_PERM = 3'd7;
  localparam D_ACCESS_ACK = 3'd0;
  localparam D_ACCESS_ACK_DATA = 3'd1;
  localparam D_GRANT = 3'd4;
  localparam D_GRANT_DATA = 3'd5;
  localparam D_RELEASE_ACK = 3'd6;
  localparam LsuL1CmdOpcode_LSU = 3'd0;
  localparam LsuL1CmdOpcode_ACCESS_1 = 3'd1;
  localparam LsuL1CmdOpcode_STORE_BUFFER = 3'd2;
  localparam LsuL1CmdOpcode_FLUSH = 3'd3;
  localparam LsuL1CmdOpcode_PREFETCH = 3'd4;
  localparam LsuPlugin_logic_flusher_enumDef_IDLE = 2'd0;
  localparam LsuPlugin_logic_flusher_enumDef_CMD = 2'd1;
  localparam LsuPlugin_logic_flusher_enumDef_COMPLETION = 2'd2;
  localparam TrapPlugin_logic_harts_0_trap_fsm_enumDef_RESET = 4'd0;
  localparam TrapPlugin_logic_harts_0_trap_fsm_enumDef_RUNNING = 4'd1;
  localparam TrapPlugin_logic_harts_0_trap_fsm_enumDef_PROCESS_1 = 4'd2;
  localparam TrapPlugin_logic_harts_0_trap_fsm_enumDef_TRAP_EPC = 4'd3;
  localparam TrapPlugin_logic_harts_0_trap_fsm_enumDef_TRAP_TVAL = 4'd4;
  localparam TrapPlugin_logic_harts_0_trap_fsm_enumDef_TRAP_TVEC = 4'd5;
  localparam TrapPlugin_logic_harts_0_trap_fsm_enumDef_TRAP_APPLY = 4'd6;
  localparam TrapPlugin_logic_harts_0_trap_fsm_enumDef_XRET_EPC = 4'd7;
  localparam TrapPlugin_logic_harts_0_trap_fsm_enumDef_XRET_APPLY = 4'd8;
  localparam TrapPlugin_logic_harts_0_trap_fsm_enumDef_ATS_RSP = 4'd9;
  localparam TrapPlugin_logic_harts_0_trap_fsm_enumDef_JUMP = 4'd10;
  localparam TrapPlugin_logic_harts_0_trap_fsm_enumDef_LSU_FLUSH = 4'd11;
  localparam TrapPlugin_logic_harts_0_trap_fsm_enumDef_FETCH_FLUSH = 4'd12;
  localparam MmuPlugin_logic_refill_enumDef_BOOT = 3'd0;
  localparam MmuPlugin_logic_refill_enumDef_IDLE = 3'd1;
  localparam MmuPlugin_logic_refill_enumDef_CMD_0 = 3'd2;
  localparam MmuPlugin_logic_refill_enumDef_CMD_1 = 3'd3;
  localparam MmuPlugin_logic_refill_enumDef_RSP_0 = 3'd4;
  localparam MmuPlugin_logic_refill_enumDef_RSP_1 = 3'd5;
  localparam CsrAccessPlugin_logic_fsm_enumDef_IDLE = 2'd0;
  localparam CsrAccessPlugin_logic_fsm_enumDef_READ = 2'd1;
  localparam CsrAccessPlugin_logic_fsm_enumDef_WRITE = 2'd2;
  localparam CsrAccessPlugin_logic_fsm_enumDef_COMPLETION = 2'd3;

  reg                 early0_DivPlugin_logic_processing_div_io_cmd_valid;
  reg                 LsuPlugin_logic_flusher_arbiter_io_output_ready;
  wire                LsuPlugin_logic_onAddress0_arbiter_io_output_ready;
  reg                 MmuPlugin_logic_refill_arbiter_io_output_ready;
  reg                 MmuPlugin_logic_invalidate_arbiter_io_output_ready;
  reg                 integer_RegFilePlugin_logic_regfile_fpga_io_writes_0_valid;
  reg        [4:0]    integer_RegFilePlugin_logic_regfile_fpga_io_writes_0_address;
  reg        [31:0]   integer_RegFilePlugin_logic_regfile_fpga_io_writes_0_data;
  wire       [30:0]   BtbPlugin_logic_ras_mem_stack_spinal_port0;
  reg        [63:0]   FetchL1Plugin_logic_banks_0_mem_spinal_port1;
  reg        [63:0]   FetchL1Plugin_logic_banks_1_mem_spinal_port1;
  reg        [21:0]   FetchL1Plugin_logic_ways_0_mem_spinal_port1;
  reg        [21:0]   FetchL1Plugin_logic_ways_1_mem_spinal_port1;
  reg        [0:0]    FetchL1Plugin_logic_plru_mem_spinal_port1;
  reg        [7:0]    GSharePlugin_logic_mem_counter_spinal_port1;
  reg        [101:0]  BtbPlugin_logic_mem_spinal_port1;
  reg        [63:0]   LsuL1Plugin_logic_banks_0_mem_spinal_port1;
  reg        [63:0]   LsuL1Plugin_logic_banks_1_mem_spinal_port1;
  reg        [21:0]   LsuL1Plugin_logic_ways_0_mem_spinal_port1;
  reg        [21:0]   LsuL1Plugin_logic_ways_1_mem_spinal_port1;
  reg        [2:0]    LsuL1Plugin_logic_shared_mem_spinal_port1;
  reg        [63:0]   LsuL1Plugin_logic_writeback_victimBuffer_spinal_port1;
  wire       [38:0]   FetchL1Plugin_logic_translationStorage_logic_sl_0_ways_0_spinal_port1;
  wire       [38:0]   FetchL1Plugin_logic_translationStorage_logic_sl_0_ways_1_spinal_port1;
  wire       [18:0]   FetchL1Plugin_logic_translationStorage_logic_sl_1_ways_0_spinal_port1;
  wire       [38:0]   LsuPlugin_logic_translationStorage_logic_sl_0_ways_0_spinal_port1;
  wire       [38:0]   LsuPlugin_logic_translationStorage_logic_sl_0_ways_1_spinal_port1;
  wire       [18:0]   LsuPlugin_logic_translationStorage_logic_sl_1_ways_0_spinal_port1;
  reg        [31:0]   CsrRamPlugin_logic_mem_spinal_port1;
  wire                early0_DivPlugin_logic_processing_div_io_cmd_ready;
  wire                early0_DivPlugin_logic_processing_div_io_rsp_valid;
  wire       [31:0]   early0_DivPlugin_logic_processing_div_io_rsp_payload_result;
  wire       [31:0]   early0_DivPlugin_logic_processing_div_io_rsp_payload_remain;
  wire                LsuPlugin_logic_flusher_arbiter_io_inputs_0_ready;
  wire                LsuPlugin_logic_flusher_arbiter_io_output_valid;
  wire       [0:0]    LsuPlugin_logic_flusher_arbiter_io_chosenOH;
  wire                streamArbiter_10_io_inputs_0_ready;
  wire                streamArbiter_10_io_inputs_1_ready;
  wire                streamArbiter_10_io_output_valid;
  wire       [31:0]   streamArbiter_10_io_output_payload_pcOnLastSlice;
  wire       [31:0]   streamArbiter_10_io_output_payload_pcTarget;
  wire                streamArbiter_10_io_output_payload_taken;
  wire                streamArbiter_10_io_output_payload_isBranch;
  wire                streamArbiter_10_io_output_payload_isPush;
  wire                streamArbiter_10_io_output_payload_isPop;
  wire                streamArbiter_10_io_output_payload_wasWrong;
  wire                streamArbiter_10_io_output_payload_badPredictedTarget;
  wire       [11:0]   streamArbiter_10_io_output_payload_history;
  wire       [15:0]   streamArbiter_10_io_output_payload_uopId;
  wire       [1:0]    streamArbiter_10_io_output_payload_ctx_GSharePlugin_GSHARE_COUNTER_0;
  wire       [1:0]    streamArbiter_10_io_output_payload_ctx_GSharePlugin_GSHARE_COUNTER_1;
  wire       [1:0]    streamArbiter_10_io_output_payload_ctx_GSharePlugin_GSHARE_COUNTER_2;
  wire       [1:0]    streamArbiter_10_io_output_payload_ctx_GSharePlugin_GSHARE_COUNTER_3;
  wire       [0:0]    streamArbiter_10_io_chosen;
  wire       [1:0]    streamArbiter_10_io_chosenOH;
  wire                LsuPlugin_logic_onAddress0_arbiter_io_inputs_0_ready;
  wire                LsuPlugin_logic_onAddress0_arbiter_io_inputs_1_ready;
  wire                LsuPlugin_logic_onAddress0_arbiter_io_inputs_2_ready;
  wire                LsuPlugin_logic_onAddress0_arbiter_io_output_valid;
  wire       [2:0]    LsuPlugin_logic_onAddress0_arbiter_io_output_payload_op;
  wire       [31:0]   LsuPlugin_logic_onAddress0_arbiter_io_output_payload_address;
  wire       [1:0]    LsuPlugin_logic_onAddress0_arbiter_io_output_payload_size;
  wire                LsuPlugin_logic_onAddress0_arbiter_io_output_payload_load;
  wire                LsuPlugin_logic_onAddress0_arbiter_io_output_payload_store;
  wire                LsuPlugin_logic_onAddress0_arbiter_io_output_payload_atomic;
  wire       [11:0]   LsuPlugin_logic_onAddress0_arbiter_io_output_payload_storeId;
  wire       [1:0]    LsuPlugin_logic_onAddress0_arbiter_io_chosen;
  wire       [2:0]    LsuPlugin_logic_onAddress0_arbiter_io_chosenOH;
  wire                MmuPlugin_logic_refill_arbiter_io_inputs_0_ready;
  wire                MmuPlugin_logic_refill_arbiter_io_output_valid;
  wire       [31:0]   MmuPlugin_logic_refill_arbiter_io_output_payload_address;
  wire       [0:0]    MmuPlugin_logic_refill_arbiter_io_output_payload_storageId;
  wire       [0:0]    MmuPlugin_logic_refill_arbiter_io_chosenOH;
  wire                MmuPlugin_logic_invalidate_arbiter_io_inputs_0_ready;
  wire                MmuPlugin_logic_invalidate_arbiter_io_output_valid;
  wire       [0:0]    MmuPlugin_logic_invalidate_arbiter_io_chosenOH;
  wire       [31:0]   integer_RegFilePlugin_logic_regfile_fpga_io_reads_0_data;
  wire       [31:0]   integer_RegFilePlugin_logic_regfile_fpga_io_reads_1_data;
  wire       [31:0]   integer_RegFilePlugin_logic_regfile_fpga_io_reads_2_data;
  wire       [31:0]   integer_RegFilePlugin_logic_regfile_fpga_io_reads_3_data;
  wire       [31:0]   _zz_early0_IntAluPlugin_logic_alu_result;
  wire       [31:0]   _zz_early0_IntAluPlugin_logic_alu_result_1;
  wire       [31:0]   _zz_early0_IntAluPlugin_logic_alu_result_2;
  wire       [31:0]   _zz_early0_IntAluPlugin_logic_alu_result_3;
  wire       [31:0]   _zz_early0_IntAluPlugin_logic_alu_result_4;
  wire       [0:0]    _zz_early0_IntAluPlugin_logic_alu_result_5;
  wire       [4:0]    _zz_early0_BarrelShifterPlugin_logic_shift_amplitude;
  wire       [31:0]   _zz_early0_BarrelShifterPlugin_logic_shift_reversed;
  wire                _zz_early0_BarrelShifterPlugin_logic_shift_reversed_1;
  wire       [0:0]    _zz_early0_BarrelShifterPlugin_logic_shift_reversed_2;
  wire       [20:0]   _zz_early0_BarrelShifterPlugin_logic_shift_reversed_3;
  wire                _zz_early0_BarrelShifterPlugin_logic_shift_reversed_4;
  wire       [0:0]    _zz_early0_BarrelShifterPlugin_logic_shift_reversed_5;
  wire       [9:0]    _zz_early0_BarrelShifterPlugin_logic_shift_reversed_6;
  wire       [32:0]   _zz_early0_BarrelShifterPlugin_logic_shift_shifted;
  wire       [32:0]   _zz_early0_BarrelShifterPlugin_logic_shift_shifted_1;
  wire       [31:0]   _zz_early0_BarrelShifterPlugin_logic_shift_patched;
  wire                _zz_early0_BarrelShifterPlugin_logic_shift_patched_1;
  wire       [0:0]    _zz_early0_BarrelShifterPlugin_logic_shift_patched_2;
  wire       [20:0]   _zz_early0_BarrelShifterPlugin_logic_shift_patched_3;
  wire                _zz_early0_BarrelShifterPlugin_logic_shift_patched_4;
  wire       [0:0]    _zz_early0_BarrelShifterPlugin_logic_shift_patched_5;
  wire       [9:0]    _zz_early0_BarrelShifterPlugin_logic_shift_patched_6;
  wire       [32:0]   _zz_toplevel_execute_ctrl2_down_MUL_SRC1_lane0;
  wire       [32:0]   _zz_toplevel_execute_ctrl2_down_MUL_SRC2_lane0;
  wire       [46:0]   _zz_toplevel_execute_ctrl3_down_early0_MulPlugin_logic_mul_VALUES_1_lane0;
  wire       [33:0]   _zz_toplevel_execute_ctrl3_down_early0_MulPlugin_logic_mul_VALUES_1_lane0_1;
  wire       [17:0]   _zz_toplevel_execute_ctrl3_down_early0_MulPlugin_logic_mul_VALUES_1_lane0_2;
  wire       [15:0]   _zz_toplevel_execute_ctrl3_down_early0_MulPlugin_logic_mul_VALUES_1_lane0_3;
  wire       [46:0]   _zz_toplevel_execute_ctrl3_down_early0_MulPlugin_logic_mul_VALUES_2_lane0;
  wire       [33:0]   _zz_toplevel_execute_ctrl3_down_early0_MulPlugin_logic_mul_VALUES_2_lane0_1;
  wire       [15:0]   _zz_toplevel_execute_ctrl3_down_early0_MulPlugin_logic_mul_VALUES_2_lane0_2;
  wire       [17:0]   _zz_toplevel_execute_ctrl3_down_early0_MulPlugin_logic_mul_VALUES_2_lane0_3;
  wire       [29:0]   _zz_toplevel_execute_ctrl3_down_early0_MulPlugin_logic_mul_VALUES_3_lane0;
  wire       [31:0]   _zz_toplevel_execute_ctrl3_down_early0_MulPlugin_logic_mul_VALUES_3_lane0_1;
  wire       [15:0]   _zz_toplevel_execute_ctrl3_down_early0_MulPlugin_logic_mul_VALUES_3_lane0_2;
  wire       [15:0]   _zz_toplevel_execute_ctrl3_down_early0_MulPlugin_logic_mul_VALUES_3_lane0_3;
  wire       [62:0]   _zz_toplevel_execute_ctrl3_down_early0_MulPlugin_logic_steps_0_adders_0_lane0_3;
  wire       [62:0]   _zz_toplevel_execute_ctrl3_down_early0_MulPlugin_logic_steps_0_adders_0_lane0_4;
  wire       [62:0]   _zz_toplevel_execute_ctrl3_down_early0_MulPlugin_logic_steps_0_adders_0_lane0_5;
  wire       [62:0]   _zz_toplevel_execute_ctrl3_down_early0_MulPlugin_logic_steps_0_adders_0_lane0_6;
  wire       [4:0]    _zz_toplevel_execute_ctrl3_down_early0_MulPlugin_logic_steps_0_adders_1_lane0_3;
  wire       [4:0]    _zz_toplevel_execute_ctrl3_down_early0_MulPlugin_logic_steps_0_adders_1_lane0_4;
  wire       [4:0]    _zz_toplevel_execute_ctrl3_down_early0_MulPlugin_logic_steps_0_adders_1_lane0_5;
  wire       [4:0]    _zz_toplevel_execute_ctrl3_down_early0_MulPlugin_logic_steps_0_adders_1_lane0_6;
  wire       [31:0]   _zz_toplevel_execute_ctrl2_down_RsUnsignedPlugin_RS1_UNSIGNED_lane0;
  wire       [0:0]    _zz_toplevel_execute_ctrl2_down_RsUnsignedPlugin_RS1_UNSIGNED_lane0_1;
  wire       [31:0]   _zz_toplevel_execute_ctrl2_down_RsUnsignedPlugin_RS2_UNSIGNED_lane0;
  wire       [0:0]    _zz_toplevel_execute_ctrl2_down_RsUnsignedPlugin_RS2_UNSIGNED_lane0_1;
  wire       [31:0]   _zz_toplevel_execute_ctrl2_down_DivPlugin_DIV_RESULT_lane0_1;
  wire       [31:0]   _zz_toplevel_execute_ctrl2_down_DivPlugin_DIV_RESULT_lane0_2;
  wire       [0:0]    _zz_toplevel_execute_ctrl2_down_DivPlugin_DIV_RESULT_lane0_3;
  wire       [31:0]   _zz_late0_IntAluPlugin_logic_alu_result;
  wire       [31:0]   _zz_late0_IntAluPlugin_logic_alu_result_1;
  wire       [31:0]   _zz_late0_IntAluPlugin_logic_alu_result_2;
  wire       [31:0]   _zz_late0_IntAluPlugin_logic_alu_result_3;
  wire       [31:0]   _zz_late0_IntAluPlugin_logic_alu_result_4;
  wire       [0:0]    _zz_late0_IntAluPlugin_logic_alu_result_5;
  wire       [4:0]    _zz_late0_BarrelShifterPlugin_logic_shift_amplitude;
  wire       [31:0]   _zz_late0_BarrelShifterPlugin_logic_shift_reversed;
  wire                _zz_late0_BarrelShifterPlugin_logic_shift_reversed_1;
  wire       [0:0]    _zz_late0_BarrelShifterPlugin_logic_shift_reversed_2;
  wire       [20:0]   _zz_late0_BarrelShifterPlugin_logic_shift_reversed_3;
  wire                _zz_late0_BarrelShifterPlugin_logic_shift_reversed_4;
  wire       [0:0]    _zz_late0_BarrelShifterPlugin_logic_shift_reversed_5;
  wire       [9:0]    _zz_late0_BarrelShifterPlugin_logic_shift_reversed_6;
  wire       [32:0]   _zz_late0_BarrelShifterPlugin_logic_shift_shifted;
  wire       [32:0]   _zz_late0_BarrelShifterPlugin_logic_shift_shifted_1;
  wire       [31:0]   _zz_late0_BarrelShifterPlugin_logic_shift_patched;
  wire                _zz_late0_BarrelShifterPlugin_logic_shift_patched_1;
  wire       [0:0]    _zz_late0_BarrelShifterPlugin_logic_shift_patched_2;
  wire       [20:0]   _zz_late0_BarrelShifterPlugin_logic_shift_patched_3;
  wire                _zz_late0_BarrelShifterPlugin_logic_shift_patched_4;
  wire       [0:0]    _zz_late0_BarrelShifterPlugin_logic_shift_patched_5;
  wire       [9:0]    _zz_late0_BarrelShifterPlugin_logic_shift_patched_6;
  wire       [31:0]   _zz_early1_IntAluPlugin_logic_alu_result;
  wire       [31:0]   _zz_early1_IntAluPlugin_logic_alu_result_1;
  wire       [31:0]   _zz_early1_IntAluPlugin_logic_alu_result_2;
  wire       [31:0]   _zz_early1_IntAluPlugin_logic_alu_result_3;
  wire       [31:0]   _zz_early1_IntAluPlugin_logic_alu_result_4;
  wire       [0:0]    _zz_early1_IntAluPlugin_logic_alu_result_5;
  wire       [4:0]    _zz_early1_BarrelShifterPlugin_logic_shift_amplitude;
  wire       [31:0]   _zz_early1_BarrelShifterPlugin_logic_shift_reversed;
  wire                _zz_early1_BarrelShifterPlugin_logic_shift_reversed_1;
  wire       [0:0]    _zz_early1_BarrelShifterPlugin_logic_shift_reversed_2;
  wire       [20:0]   _zz_early1_BarrelShifterPlugin_logic_shift_reversed_3;
  wire                _zz_early1_BarrelShifterPlugin_logic_shift_reversed_4;
  wire       [0:0]    _zz_early1_BarrelShifterPlugin_logic_shift_reversed_5;
  wire       [9:0]    _zz_early1_BarrelShifterPlugin_logic_shift_reversed_6;
  wire       [32:0]   _zz_early1_BarrelShifterPlugin_logic_shift_shifted;
  wire       [32:0]   _zz_early1_BarrelShifterPlugin_logic_shift_shifted_1;
  wire       [31:0]   _zz_early1_BarrelShifterPlugin_logic_shift_patched;
  wire                _zz_early1_BarrelShifterPlugin_logic_shift_patched_1;
  wire       [0:0]    _zz_early1_BarrelShifterPlugin_logic_shift_patched_2;
  wire       [20:0]   _zz_early1_BarrelShifterPlugin_logic_shift_patched_3;
  wire                _zz_early1_BarrelShifterPlugin_logic_shift_patched_4;
  wire       [0:0]    _zz_early1_BarrelShifterPlugin_logic_shift_patched_5;
  wire       [9:0]    _zz_early1_BarrelShifterPlugin_logic_shift_patched_6;
  wire       [31:0]   _zz_late1_IntAluPlugin_logic_alu_result;
  wire       [31:0]   _zz_late1_IntAluPlugin_logic_alu_result_1;
  wire       [31:0]   _zz_late1_IntAluPlugin_logic_alu_result_2;
  wire       [31:0]   _zz_late1_IntAluPlugin_logic_alu_result_3;
  wire       [31:0]   _zz_late1_IntAluPlugin_logic_alu_result_4;
  wire       [0:0]    _zz_late1_IntAluPlugin_logic_alu_result_5;
  wire       [4:0]    _zz_late1_BarrelShifterPlugin_logic_shift_amplitude;
  wire       [31:0]   _zz_late1_BarrelShifterPlugin_logic_shift_reversed;
  wire                _zz_late1_BarrelShifterPlugin_logic_shift_reversed_1;
  wire       [0:0]    _zz_late1_BarrelShifterPlugin_logic_shift_reversed_2;
  wire       [20:0]   _zz_late1_BarrelShifterPlugin_logic_shift_reversed_3;
  wire                _zz_late1_BarrelShifterPlugin_logic_shift_reversed_4;
  wire       [0:0]    _zz_late1_BarrelShifterPlugin_logic_shift_reversed_5;
  wire       [9:0]    _zz_late1_BarrelShifterPlugin_logic_shift_reversed_6;
  wire       [32:0]   _zz_late1_BarrelShifterPlugin_logic_shift_shifted;
  wire       [32:0]   _zz_late1_BarrelShifterPlugin_logic_shift_shifted_1;
  wire       [31:0]   _zz_late1_BarrelShifterPlugin_logic_shift_patched;
  wire                _zz_late1_BarrelShifterPlugin_logic_shift_patched_1;
  wire       [0:0]    _zz_late1_BarrelShifterPlugin_logic_shift_patched_2;
  wire       [20:0]   _zz_late1_BarrelShifterPlugin_logic_shift_patched_3;
  wire                _zz_late1_BarrelShifterPlugin_logic_shift_patched_4;
  wire       [0:0]    _zz_late1_BarrelShifterPlugin_logic_shift_patched_5;
  wire       [9:0]    _zz_late1_BarrelShifterPlugin_logic_shift_patched_6;
  wire       [20:0]   _zz_early0_BranchPlugin_pcCalc_target_b;
  wire       [11:0]   _zz_early0_BranchPlugin_pcCalc_target_b_1;
  wire       [12:0]   _zz_early0_BranchPlugin_pcCalc_target_b_2;
  wire       [31:0]   _zz_toplevel_execute_ctrl2_down_early0_BranchPlugin_pcCalc_PC_TRUE_lane0;
  wire       [31:0]   _zz_toplevel_execute_ctrl2_down_early0_BranchPlugin_pcCalc_PC_FALSE_lane0;
  wire       [2:0]    _zz_toplevel_execute_ctrl2_down_early0_BranchPlugin_pcCalc_PC_FALSE_lane0_1;
  wire       [31:0]   _zz_toplevel_execute_ctrl2_down_early0_BranchPlugin_pcCalc_PC_LAST_SLICE_lane0;
  wire       [1:0]    _zz_toplevel_execute_ctrl2_down_early0_BranchPlugin_pcCalc_PC_LAST_SLICE_lane0_1;
  wire       [20:0]   _zz_early1_BranchPlugin_pcCalc_target_b;
  wire       [11:0]   _zz_early1_BranchPlugin_pcCalc_target_b_1;
  wire       [12:0]   _zz_early1_BranchPlugin_pcCalc_target_b_2;
  wire       [31:0]   _zz_toplevel_execute_ctrl2_down_early1_BranchPlugin_pcCalc_PC_TRUE_lane1;
  wire       [31:0]   _zz_toplevel_execute_ctrl2_down_early1_BranchPlugin_pcCalc_PC_FALSE_lane1;
  wire       [2:0]    _zz_toplevel_execute_ctrl2_down_early1_BranchPlugin_pcCalc_PC_FALSE_lane1_1;
  wire       [31:0]   _zz_toplevel_execute_ctrl2_down_early1_BranchPlugin_pcCalc_PC_LAST_SLICE_lane1;
  wire       [1:0]    _zz_toplevel_execute_ctrl2_down_early1_BranchPlugin_pcCalc_PC_LAST_SLICE_lane1_1;
  reg        [3:0]    _zz_fetch_logic_ctrls_2_down_AlignerPlugin_logic_FETCH_MASK;
  wire       [1:0]    _zz_fetch_logic_ctrls_2_down_AlignerPlugin_logic_FETCH_MASK_1;
  reg        [3:0]    _zz_fetch_logic_ctrls_2_down_AlignerPlugin_logic_FETCH_MASK_2;
  wire       [3:0]    _zz_fetch_logic_ctrls_2_down_AlignerPlugin_logic_FETCH_LAST;
  wire                _zz_AlignerPlugin_logic_extractors_0_usableMask;
  wire                _zz_AlignerPlugin_logic_extractors_0_usableMask_1;
  wire                _zz_AlignerPlugin_logic_extractors_0_usableMask_2;
  wire       [0:0]    _zz_AlignerPlugin_logic_extractors_0_usableMask_3;
  wire       [0:0]    _zz_AlignerPlugin_logic_extractors_0_usableMask_4;
  wire       [0:0]    _zz_AlignerPlugin_logic_extractors_0_redo_8;
  wire       [0:0]    _zz_AlignerPlugin_logic_extractors_0_redo_9;
  wire       [0:0]    _zz_AlignerPlugin_logic_extractors_0_redo_10;
  wire       [0:0]    _zz_AlignerPlugin_logic_extractors_0_redo_11;
  wire       [0:0]    _zz_AlignerPlugin_logic_extractors_0_redo_12;
  wire       [0:0]    _zz_AlignerPlugin_logic_extractors_0_redo_13;
  wire       [0:0]    _zz_AlignerPlugin_logic_extractors_0_redo_14;
  wire       [0:0]    _zz_AlignerPlugin_logic_extractors_0_redo_15;
  wire       [0:0]    _zz_AlignerPlugin_logic_extractors_0_redo_16;
  wire       [0:0]    _zz_AlignerPlugin_logic_extractors_0_redo_17;
  wire       [0:0]    _zz_AlignerPlugin_logic_extractors_0_redo_18;
  wire       [0:0]    _zz_AlignerPlugin_logic_extractors_0_redo_19;
  wire       [0:0]    _zz_AlignerPlugin_logic_extractors_0_redo_20;
  wire       [0:0]    _zz_AlignerPlugin_logic_extractors_0_redo_21;
  wire       [0:0]    _zz_AlignerPlugin_logic_extractors_0_redo_22;
  wire       [0:0]    _zz_AlignerPlugin_logic_extractors_0_redo_23;
  wire       [0:0]    _zz_AlignerPlugin_logic_extractors_0_redo_24;
  wire       [0:0]    _zz_AlignerPlugin_logic_extractors_0_localMask;
  wire       [0:0]    _zz_AlignerPlugin_logic_extractors_0_localMask_1;
  wire       [0:0]    _zz_AlignerPlugin_logic_extractors_0_localMask_2;
  wire       [0:0]    _zz_AlignerPlugin_logic_extractors_0_localMask_3;
  wire       [0:0]    _zz_AlignerPlugin_logic_extractors_0_localMask_4;
  wire       [0:0]    _zz_AlignerPlugin_logic_extractors_0_localMask_5;
  wire       [0:0]    _zz_AlignerPlugin_logic_extractors_0_localMask_6;
  wire       [0:0]    _zz_AlignerPlugin_logic_extractors_0_localMask_7;
  wire       [0:0]    _zz_AlignerPlugin_logic_extractors_0_localMask_8;
  wire       [0:0]    _zz_AlignerPlugin_logic_extractors_0_localMask_9;
  wire       [0:0]    _zz_AlignerPlugin_logic_extractors_0_localMask_10;
  wire       [0:0]    _zz_AlignerPlugin_logic_extractors_0_localMask_11;
  wire       [0:0]    _zz_AlignerPlugin_logic_extractors_0_localMask_12;
  wire       [0:0]    _zz_AlignerPlugin_logic_extractors_0_localMask_13;
  wire       [0:0]    _zz_AlignerPlugin_logic_extractors_0_localMask_14;
  wire       [0:0]    _zz_AlignerPlugin_logic_extractors_0_localMask_15;
  wire                _zz_AlignerPlugin_logic_extractors_1_usableMask;
  wire                _zz_AlignerPlugin_logic_extractors_1_usableMask_1;
  wire                _zz_AlignerPlugin_logic_extractors_1_usableMask_2;
  wire                _zz_AlignerPlugin_logic_extractors_1_usableMask_3;
  wire       [0:0]    _zz_AlignerPlugin_logic_extractors_1_redo_7;
  wire       [0:0]    _zz_AlignerPlugin_logic_extractors_1_redo_8;
  wire       [0:0]    _zz_AlignerPlugin_logic_extractors_1_redo_9;
  wire       [0:0]    _zz_AlignerPlugin_logic_extractors_1_redo_10;
  wire       [0:0]    _zz_AlignerPlugin_logic_extractors_1_redo_11;
  wire       [0:0]    _zz_AlignerPlugin_logic_extractors_1_redo_12;
  wire       [0:0]    _zz_AlignerPlugin_logic_extractors_1_redo_13;
  wire       [0:0]    _zz_AlignerPlugin_logic_extractors_1_redo_14;
  wire       [0:0]    _zz_AlignerPlugin_logic_extractors_1_redo_15;
  wire       [0:0]    _zz_AlignerPlugin_logic_extractors_1_redo_16;
  wire       [0:0]    _zz_AlignerPlugin_logic_extractors_1_redo_17;
  wire       [0:0]    _zz_AlignerPlugin_logic_extractors_1_redo_18;
  wire       [0:0]    _zz_AlignerPlugin_logic_extractors_1_redo_19;
  wire       [0:0]    _zz_AlignerPlugin_logic_extractors_1_localMask;
  wire       [0:0]    _zz_AlignerPlugin_logic_extractors_1_localMask_1;
  wire       [0:0]    _zz_AlignerPlugin_logic_extractors_1_localMask_2;
  wire       [0:0]    _zz_AlignerPlugin_logic_extractors_1_localMask_3;
  wire       [0:0]    _zz_AlignerPlugin_logic_extractors_1_localMask_4;
  wire       [0:0]    _zz_AlignerPlugin_logic_extractors_1_localMask_5;
  wire       [0:0]    _zz_AlignerPlugin_logic_extractors_1_localMask_6;
  wire       [0:0]    _zz_AlignerPlugin_logic_extractors_1_localMask_7;
  wire       [0:0]    _zz_AlignerPlugin_logic_extractors_1_localMask_8;
  wire       [0:0]    _zz_AlignerPlugin_logic_extractors_1_localMask_9;
  wire       [0:0]    _zz_AlignerPlugin_logic_extractors_1_localMask_10;
  wire       [0:0]    _zz_AlignerPlugin_logic_extractors_1_localMask_11;
  wire       [4:0]    _zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_23;
  wire       [0:0]    _zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_24;
  wire                _zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_25;
  wire       [31:0]   _zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_26;
  wire       [11:0]   _zz__zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_22;
  wire       [5:0]    _zz__zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_22_1;
  reg        [31:0]   _zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_27;
  wire       [1:0]    _zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_28;
  reg        [2:0]    _zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_29;
  wire       [2:0]    _zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_30;
  wire       [6:0]    _zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_31;
  wire       [4:0]    _zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_32;
  wire                _zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_33;
  wire       [4:0]    _zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_34;
  wire       [11:0]   _zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_35;
  wire       [11:0]   _zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_36;
  wire       [1:0]    _zz__zz_toplevel_decode_ctrls_0_up_Decode_INSTRUCTION_SLICE_COUNT_0_5;
  wire       [1:0]    _zz_AlignerPlugin_logic_feeder_lanes_0_onBtb_pcLastSlice;
  wire       [4:0]    _zz_AlignerPlugin_logic_feeder_lanes_1_withRvc_dec_inst_23;
  wire       [0:0]    _zz_AlignerPlugin_logic_feeder_lanes_1_withRvc_dec_inst_24;
  wire                _zz_AlignerPlugin_logic_feeder_lanes_1_withRvc_dec_inst_25;
  wire       [31:0]   _zz_AlignerPlugin_logic_feeder_lanes_1_withRvc_dec_inst_26;
  wire       [11:0]   _zz__zz_AlignerPlugin_logic_feeder_lanes_1_withRvc_dec_inst_22;
  wire       [5:0]    _zz__zz_AlignerPlugin_logic_feeder_lanes_1_withRvc_dec_inst_22_1;
  reg        [31:0]   _zz_AlignerPlugin_logic_feeder_lanes_1_withRvc_dec_inst_27;
  wire       [1:0]    _zz_AlignerPlugin_logic_feeder_lanes_1_withRvc_dec_inst_28;
  reg        [2:0]    _zz_AlignerPlugin_logic_feeder_lanes_1_withRvc_dec_inst_29;
  wire       [2:0]    _zz_AlignerPlugin_logic_feeder_lanes_1_withRvc_dec_inst_30;
  wire       [6:0]    _zz_AlignerPlugin_logic_feeder_lanes_1_withRvc_dec_inst_31;
  wire       [4:0]    _zz_AlignerPlugin_logic_feeder_lanes_1_withRvc_dec_inst_32;
  wire                _zz_AlignerPlugin_logic_feeder_lanes_1_withRvc_dec_inst_33;
  wire       [4:0]    _zz_AlignerPlugin_logic_feeder_lanes_1_withRvc_dec_inst_34;
  wire       [11:0]   _zz_AlignerPlugin_logic_feeder_lanes_1_withRvc_dec_inst_35;
  wire       [11:0]   _zz_AlignerPlugin_logic_feeder_lanes_1_withRvc_dec_inst_36;
  wire       [1:0]    _zz__zz_toplevel_decode_ctrls_0_up_Decode_INSTRUCTION_SLICE_COUNT_1_5;
  wire       [9:0]    _zz_toplevel_decode_ctrls_0_up_Decode_DOP_ID_1;
  wire       [0:0]    _zz_toplevel_decode_ctrls_0_up_Decode_DOP_ID_1_1;
  wire       [1:0]    _zz_AlignerPlugin_logic_feeder_lanes_1_onBtb_pcLastSlice;
  wire       [21:0]   _zz_FetchL1Plugin_logic_ways_0_mem_port;
  wire                _zz_FetchL1Plugin_logic_ways_0_mem_port_1;
  wire       [21:0]   _zz_FetchL1Plugin_logic_ways_1_mem_port;
  wire                _zz_FetchL1Plugin_logic_ways_1_mem_port_1;
  wire                _zz_when;
  wire       [19:0]   _zz_FetchL1Plugin_logic_hits_w_0_indirect_bypassHits;
  wire       [19:0]   _zz_FetchL1Plugin_logic_hits_w_1_indirect_bypassHits;
  wire       [0:0]    _zz_FetchL1Plugin_logic_ctrl_dataAccessFault;
  wire       [0:0]    _zz_FetchL1Plugin_logic_plru_write_payload_data_0;
  wire       [7:0]    _zz_GSharePlugin_logic_mem_counter_port;
  wire                _zz_fetch_logic_ctrls_0_down_GSharePlugin_logic_HASH_1;
  wire       [0:0]    _zz_fetch_logic_ctrls_0_down_GSharePlugin_logic_HASH_2;
  wire       [3:0]    _zz_fetch_logic_ctrls_0_down_GSharePlugin_logic_HASH_3;
  wire       [1:0]    _zz_BtbPlugin_logic_ras_ptr_push;
  wire       [1:0]    _zz_BtbPlugin_logic_ras_ptr_push_1;
  wire       [0:0]    _zz_BtbPlugin_logic_ras_ptr_push_2;
  wire       [1:0]    _zz_BtbPlugin_logic_ras_ptr_push_3;
  wire       [0:0]    _zz_BtbPlugin_logic_ras_ptr_push_4;
  wire       [1:0]    _zz_BtbPlugin_logic_ras_ptr_pop_aheadValue;
  wire       [1:0]    _zz_BtbPlugin_logic_ras_ptr_pop_aheadValue_1;
  wire       [0:0]    _zz_BtbPlugin_logic_ras_ptr_pop_aheadValue_2;
  wire       [1:0]    _zz_BtbPlugin_logic_ras_ptr_pop_aheadValue_3;
  wire       [0:0]    _zz_BtbPlugin_logic_ras_ptr_pop_aheadValue_4;
  wire       [30:0]   _zz_BtbPlugin_logic_ras_mem_stack_port;
  wire       [63:0]   _zz_WhiteboxerPlugin_logic_decodes_0_pc;
  wire       [63:0]   _zz_WhiteboxerPlugin_logic_decodes_1_pc;
  wire       [31:0]   _zz_early0_BranchPlugin_logic_alu_expectedMsb;
  wire       [12:0]   _zz_early0_BranchPlugin_logic_jumpLogic_history_fromFetch_shifter_1;
  wire       [12:0]   _zz_early0_BranchPlugin_logic_jumpLogic_history_fromFetch_shifter_2;
  wire       [12:0]   _zz_early0_BranchPlugin_logic_jumpLogic_history_fromFetch_shifter_3;
  wire       [12:0]   _zz_early0_BranchPlugin_logic_jumpLogic_history_fromFetch_shifter_4;
  wire       [3:0]    _zz_early0_EnvPlugin_logic_trapPort_payload_code;
  wire       [31:0]   _zz_early1_BranchPlugin_logic_alu_expectedMsb;
  wire       [12:0]   _zz_early1_BranchPlugin_logic_jumpLogic_history_fromFetch_shifter_1;
  wire       [12:0]   _zz_early1_BranchPlugin_logic_jumpLogic_history_fromFetch_shifter_2;
  wire       [12:0]   _zz_early1_BranchPlugin_logic_jumpLogic_history_fromFetch_shifter_3;
  wire       [12:0]   _zz_early1_BranchPlugin_logic_jumpLogic_history_fromFetch_shifter_4;
  wire       [11:0]   _zz__zz_toplevel_execute_ctrl1_down_early0_SrcPlugin_SRC2_lane0;
  wire       [11:0]   _zz__zz_toplevel_execute_ctrl1_down_early0_SrcPlugin_SRC2_lane0_1;
  wire       [31:0]   _zz_toplevel_execute_ctrl2_down_early0_SrcPlugin_ADD_SUB_lane0;
  wire       [31:0]   _zz_toplevel_execute_ctrl2_down_early0_SrcPlugin_ADD_SUB_lane0_1;
  wire       [31:0]   _zz_toplevel_execute_ctrl2_down_early0_SrcPlugin_ADD_SUB_lane0_2;
  wire       [0:0]    _zz_toplevel_execute_ctrl2_down_early0_SrcPlugin_ADD_SUB_lane0_3;
  wire       [11:0]   _zz__zz_toplevel_execute_ctrl3_down_late0_SrcPlugin_SRC2_lane0;
  wire       [31:0]   _zz_toplevel_execute_ctrl4_down_late0_SrcPlugin_ADD_SUB_lane0;
  wire       [31:0]   _zz_toplevel_execute_ctrl4_down_late0_SrcPlugin_ADD_SUB_lane0_1;
  wire       [31:0]   _zz_toplevel_execute_ctrl4_down_late0_SrcPlugin_ADD_SUB_lane0_2;
  wire       [0:0]    _zz_toplevel_execute_ctrl4_down_late0_SrcPlugin_ADD_SUB_lane0_3;
  wire       [11:0]   _zz__zz_toplevel_execute_ctrl1_down_early1_SrcPlugin_SRC2_lane1;
  wire       [31:0]   _zz_toplevel_execute_ctrl2_down_early1_SrcPlugin_ADD_SUB_lane1;
  wire       [31:0]   _zz_toplevel_execute_ctrl2_down_early1_SrcPlugin_ADD_SUB_lane1_1;
  wire       [31:0]   _zz_toplevel_execute_ctrl2_down_early1_SrcPlugin_ADD_SUB_lane1_2;
  wire       [0:0]    _zz_toplevel_execute_ctrl2_down_early1_SrcPlugin_ADD_SUB_lane1_3;
  wire       [11:0]   _zz__zz_toplevel_execute_ctrl3_down_late1_SrcPlugin_SRC2_lane1;
  wire       [31:0]   _zz_toplevel_execute_ctrl4_down_late1_SrcPlugin_ADD_SUB_lane1;
  wire       [31:0]   _zz_toplevel_execute_ctrl4_down_late1_SrcPlugin_ADD_SUB_lane1_1;
  wire       [31:0]   _zz_toplevel_execute_ctrl4_down_late1_SrcPlugin_ADD_SUB_lane1_2;
  wire       [0:0]    _zz_toplevel_execute_ctrl4_down_late1_SrcPlugin_ADD_SUB_lane1_3;
  wire       [31:0]   _zz_late0_BranchPlugin_logic_alu_expectedMsb;
  wire       [12:0]   _zz_late0_BranchPlugin_logic_jumpLogic_history_fromFetch_shifter_1;
  wire       [12:0]   _zz_late0_BranchPlugin_logic_jumpLogic_history_fromFetch_shifter_2;
  wire       [12:0]   _zz_late0_BranchPlugin_logic_jumpLogic_history_fromFetch_shifter_3;
  wire       [12:0]   _zz_late0_BranchPlugin_logic_jumpLogic_history_fromFetch_shifter_4;
  wire       [31:0]   _zz_late1_BranchPlugin_logic_alu_expectedMsb;
  wire       [12:0]   _zz_late1_BranchPlugin_logic_jumpLogic_history_fromFetch_shifter_1;
  wire       [12:0]   _zz_late1_BranchPlugin_logic_jumpLogic_history_fromFetch_shifter_2;
  wire       [12:0]   _zz_late1_BranchPlugin_logic_jumpLogic_history_fromFetch_shifter_3;
  wire       [12:0]   _zz_late1_BranchPlugin_logic_jumpLogic_history_fromFetch_shifter_4;
  wire                _zz_GSharePlugin_logic_onLearn_hash_1;
  wire       [0:0]    _zz_GSharePlugin_logic_onLearn_hash_2;
  wire       [3:0]    _zz_GSharePlugin_logic_onLearn_hash_3;
  wire       [101:0]  _zz_BtbPlugin_logic_mem_port;
  wire       [28:0]   _zz_BtbPlugin_logic_onLearn_port_payload_address;
  wire       [0:0]    _zz_toplevel_decode_ctrls_1_down_RS1_ENABLE_0;
  wire       [0:0]    _zz_toplevel_decode_ctrls_1_down_RS2_ENABLE_0;
  wire       [0:0]    _zz_toplevel_decode_ctrls_1_down_RD_ENABLE_0;
  wire       [31:0]   _zz_toplevel_decode_ctrls_1_down_RD_ENABLE_0_1;
  wire       [31:0]   _zz_toplevel_decode_ctrls_1_down_RD_ENABLE_0_2;
  wire       [31:0]   _zz_toplevel_decode_ctrls_1_down_RD_ENABLE_0_3;
  wire                _zz_toplevel_decode_ctrls_1_down_RD_ENABLE_0_4;
  wire       [31:0]   _zz_toplevel_decode_ctrls_1_down_Decode_LEGAL_0;
  wire       [31:0]   _zz_toplevel_decode_ctrls_1_down_Decode_LEGAL_0_1;
  wire       [31:0]   _zz_toplevel_decode_ctrls_1_down_Decode_LEGAL_0_2;
  wire                _zz_toplevel_decode_ctrls_1_down_Decode_LEGAL_0_3;
  wire       [0:0]    _zz_toplevel_decode_ctrls_1_down_Decode_LEGAL_0_4;
  wire       [17:0]   _zz_toplevel_decode_ctrls_1_down_Decode_LEGAL_0_5;
  wire       [31:0]   _zz_toplevel_decode_ctrls_1_down_Decode_LEGAL_0_6;
  wire       [31:0]   _zz_toplevel_decode_ctrls_1_down_Decode_LEGAL_0_7;
  wire       [31:0]   _zz_toplevel_decode_ctrls_1_down_Decode_LEGAL_0_8;
  wire                _zz_toplevel_decode_ctrls_1_down_Decode_LEGAL_0_9;
  wire       [0:0]    _zz_toplevel_decode_ctrls_1_down_Decode_LEGAL_0_10;
  wire       [11:0]   _zz_toplevel_decode_ctrls_1_down_Decode_LEGAL_0_11;
  wire       [31:0]   _zz_toplevel_decode_ctrls_1_down_Decode_LEGAL_0_12;
  wire       [31:0]   _zz_toplevel_decode_ctrls_1_down_Decode_LEGAL_0_13;
  wire       [31:0]   _zz_toplevel_decode_ctrls_1_down_Decode_LEGAL_0_14;
  wire                _zz_toplevel_decode_ctrls_1_down_Decode_LEGAL_0_15;
  wire       [0:0]    _zz_toplevel_decode_ctrls_1_down_Decode_LEGAL_0_16;
  wire       [5:0]    _zz_toplevel_decode_ctrls_1_down_Decode_LEGAL_0_17;
  wire       [31:0]   _zz_toplevel_decode_ctrls_1_down_Decode_LEGAL_0_18;
  wire       [31:0]   _zz_toplevel_decode_ctrls_1_down_Decode_LEGAL_0_19;
  wire       [31:0]   _zz_toplevel_decode_ctrls_1_down_Decode_LEGAL_0_20;
  wire                _zz_toplevel_decode_ctrls_1_down_Decode_LEGAL_0_21;
  wire                _zz_toplevel_decode_ctrls_1_down_Decode_LEGAL_0_22;
  wire       [0:0]    _zz_DecoderPlugin_logic_laneLogic_0_fixer_isJb;
  wire       [31:0]   _zz_DecoderPlugin_logic_forgetPort_payload_pcOnLastSlice;
  wire       [1:0]    _zz_DecoderPlugin_logic_forgetPort_payload_pcOnLastSlice_1;
  wire       [1:0]    _zz_DecoderPlugin_logic_forgetPort_payload_pcOnLastSlice_2;
  wire       [0:0]    _zz_toplevel_decode_ctrls_1_down_RS1_ENABLE_1;
  wire       [0:0]    _zz_toplevel_decode_ctrls_1_down_RS2_ENABLE_1;
  wire       [0:0]    _zz_toplevel_decode_ctrls_1_down_RD_ENABLE_1;
  wire       [31:0]   _zz_toplevel_decode_ctrls_1_down_RD_ENABLE_1_1;
  wire       [31:0]   _zz_toplevel_decode_ctrls_1_down_RD_ENABLE_1_2;
  wire       [31:0]   _zz_toplevel_decode_ctrls_1_down_RD_ENABLE_1_3;
  wire                _zz_toplevel_decode_ctrls_1_down_RD_ENABLE_1_4;
  wire       [31:0]   _zz_toplevel_decode_ctrls_1_down_Decode_LEGAL_1;
  wire       [31:0]   _zz_toplevel_decode_ctrls_1_down_Decode_LEGAL_1_1;
  wire       [31:0]   _zz_toplevel_decode_ctrls_1_down_Decode_LEGAL_1_2;
  wire                _zz_toplevel_decode_ctrls_1_down_Decode_LEGAL_1_3;
  wire       [0:0]    _zz_toplevel_decode_ctrls_1_down_Decode_LEGAL_1_4;
  wire       [17:0]   _zz_toplevel_decode_ctrls_1_down_Decode_LEGAL_1_5;
  wire       [31:0]   _zz_toplevel_decode_ctrls_1_down_Decode_LEGAL_1_6;
  wire       [31:0]   _zz_toplevel_decode_ctrls_1_down_Decode_LEGAL_1_7;
  wire       [31:0]   _zz_toplevel_decode_ctrls_1_down_Decode_LEGAL_1_8;
  wire                _zz_toplevel_decode_ctrls_1_down_Decode_LEGAL_1_9;
  wire       [0:0]    _zz_toplevel_decode_ctrls_1_down_Decode_LEGAL_1_10;
  wire       [11:0]   _zz_toplevel_decode_ctrls_1_down_Decode_LEGAL_1_11;
  wire       [31:0]   _zz_toplevel_decode_ctrls_1_down_Decode_LEGAL_1_12;
  wire       [31:0]   _zz_toplevel_decode_ctrls_1_down_Decode_LEGAL_1_13;
  wire       [31:0]   _zz_toplevel_decode_ctrls_1_down_Decode_LEGAL_1_14;
  wire                _zz_toplevel_decode_ctrls_1_down_Decode_LEGAL_1_15;
  wire       [0:0]    _zz_toplevel_decode_ctrls_1_down_Decode_LEGAL_1_16;
  wire       [5:0]    _zz_toplevel_decode_ctrls_1_down_Decode_LEGAL_1_17;
  wire       [31:0]   _zz_toplevel_decode_ctrls_1_down_Decode_LEGAL_1_18;
  wire       [31:0]   _zz_toplevel_decode_ctrls_1_down_Decode_LEGAL_1_19;
  wire       [31:0]   _zz_toplevel_decode_ctrls_1_down_Decode_LEGAL_1_20;
  wire                _zz_toplevel_decode_ctrls_1_down_Decode_LEGAL_1_21;
  wire                _zz_toplevel_decode_ctrls_1_down_Decode_LEGAL_1_22;
  wire       [0:0]    _zz_DecoderPlugin_logic_laneLogic_1_fixer_isJb;
  wire       [31:0]   _zz_DecoderPlugin_logic_forgetPort_payload_pcOnLastSlice_3;
  wire       [1:0]    _zz_DecoderPlugin_logic_forgetPort_payload_pcOnLastSlice_4;
  wire       [1:0]    _zz_DecoderPlugin_logic_forgetPort_payload_pcOnLastSlice_5;
  wire       [11:0]   _zz_CsrRamPlugin_csrMapper_ramAddress_1;
  wire       [11:0]   _zz_CsrRamPlugin_csrMapper_ramAddress_2;
  reg        [0:0]    _zz_DispatchPlugin_logic_candidates_1_age;
  wire       [0:0]    _zz_DispatchPlugin_logic_candidates_1_age_1;
  reg        [1:0]    _zz_DispatchPlugin_logic_candidates_2_age;
  wire       [1:0]    _zz_DispatchPlugin_logic_candidates_2_age_1;
  wire                _zz_DispatchPlugin_logic_rsHazardChecker_0_onLl_0_onRs_0_hazard;
  wire                _zz_DispatchPlugin_logic_rsHazardChecker_0_onLl_0_onRs_0_hazard_1;
  wire                _zz_DispatchPlugin_logic_rsHazardChecker_0_onLl_0_onRs_0_hazard_2;
  wire                _zz_DispatchPlugin_logic_rsHazardChecker_0_onLl_0_onRs_0_hazard_3;
  wire                _zz_DispatchPlugin_logic_rsHazardChecker_0_onLl_0_onRs_0_hazard_4;
  wire                _zz_DispatchPlugin_logic_rsHazardChecker_0_onLl_0_onRs_0_hazard_5;
  wire                _zz_DispatchPlugin_logic_rsHazardChecker_0_onLl_0_onRs_1_hazard;
  wire                _zz_DispatchPlugin_logic_rsHazardChecker_0_onLl_0_onRs_1_hazard_1;
  wire                _zz_DispatchPlugin_logic_rsHazardChecker_0_onLl_0_onRs_1_hazard_2;
  wire                _zz_DispatchPlugin_logic_rsHazardChecker_0_onLl_0_onRs_1_hazard_3;
  wire                _zz_DispatchPlugin_logic_rsHazardChecker_0_onLl_0_onRs_1_hazard_4;
  wire                _zz_DispatchPlugin_logic_rsHazardChecker_0_onLl_0_onRs_1_hazard_5;
  wire                _zz_DispatchPlugin_logic_rsHazardChecker_0_onLl_1_onRs_0_hazard;
  wire                _zz_DispatchPlugin_logic_rsHazardChecker_0_onLl_1_onRs_0_hazard_1;
  wire                _zz_DispatchPlugin_logic_rsHazardChecker_0_onLl_1_onRs_0_hazard_2;
  wire                _zz_DispatchPlugin_logic_rsHazardChecker_0_onLl_1_onRs_0_hazard_3;
  wire                _zz_DispatchPlugin_logic_rsHazardChecker_0_onLl_1_onRs_0_hazard_4;
  wire                _zz_DispatchPlugin_logic_rsHazardChecker_0_onLl_1_onRs_0_hazard_5;
  wire                _zz_DispatchPlugin_logic_rsHazardChecker_0_onLl_1_onRs_1_hazard;
  wire                _zz_DispatchPlugin_logic_rsHazardChecker_0_onLl_1_onRs_1_hazard_1;
  wire                _zz_DispatchPlugin_logic_rsHazardChecker_0_onLl_1_onRs_1_hazard_2;
  wire                _zz_DispatchPlugin_logic_rsHazardChecker_0_onLl_1_onRs_1_hazard_3;
  wire                _zz_DispatchPlugin_logic_rsHazardChecker_0_onLl_1_onRs_1_hazard_4;
  wire                _zz_DispatchPlugin_logic_rsHazardChecker_0_onLl_1_onRs_1_hazard_5;
  wire                _zz_DispatchPlugin_logic_rsHazardChecker_1_onLl_0_onRs_0_hazard;
  wire                _zz_DispatchPlugin_logic_rsHazardChecker_1_onLl_0_onRs_0_hazard_1;
  wire                _zz_DispatchPlugin_logic_rsHazardChecker_1_onLl_0_onRs_0_hazard_2;
  wire                _zz_DispatchPlugin_logic_rsHazardChecker_1_onLl_0_onRs_0_hazard_3;
  wire                _zz_DispatchPlugin_logic_rsHazardChecker_1_onLl_0_onRs_0_hazard_4;
  wire                _zz_DispatchPlugin_logic_rsHazardChecker_1_onLl_0_onRs_0_hazard_5;
  wire                _zz_DispatchPlugin_logic_rsHazardChecker_1_onLl_0_onRs_1_hazard;
  wire                _zz_DispatchPlugin_logic_rsHazardChecker_1_onLl_0_onRs_1_hazard_1;
  wire                _zz_DispatchPlugin_logic_rsHazardChecker_1_onLl_0_onRs_1_hazard_2;
  wire                _zz_DispatchPlugin_logic_rsHazardChecker_1_onLl_0_onRs_1_hazard_3;
  wire                _zz_DispatchPlugin_logic_rsHazardChecker_1_onLl_0_onRs_1_hazard_4;
  wire                _zz_DispatchPlugin_logic_rsHazardChecker_1_onLl_0_onRs_1_hazard_5;
  wire                _zz_DispatchPlugin_logic_rsHazardChecker_1_onLl_1_onRs_0_hazard;
  wire                _zz_DispatchPlugin_logic_rsHazardChecker_1_onLl_1_onRs_0_hazard_1;
  wire                _zz_DispatchPlugin_logic_rsHazardChecker_1_onLl_1_onRs_0_hazard_2;
  wire                _zz_DispatchPlugin_logic_rsHazardChecker_1_onLl_1_onRs_0_hazard_3;
  wire                _zz_DispatchPlugin_logic_rsHazardChecker_1_onLl_1_onRs_0_hazard_4;
  wire                _zz_DispatchPlugin_logic_rsHazardChecker_1_onLl_1_onRs_0_hazard_5;
  wire                _zz_DispatchPlugin_logic_rsHazardChecker_1_onLl_1_onRs_1_hazard;
  wire                _zz_DispatchPlugin_logic_rsHazardChecker_1_onLl_1_onRs_1_hazard_1;
  wire                _zz_DispatchPlugin_logic_rsHazardChecker_1_onLl_1_onRs_1_hazard_2;
  wire                _zz_DispatchPlugin_logic_rsHazardChecker_1_onLl_1_onRs_1_hazard_3;
  wire                _zz_DispatchPlugin_logic_rsHazardChecker_1_onLl_1_onRs_1_hazard_4;
  wire                _zz_DispatchPlugin_logic_rsHazardChecker_1_onLl_1_onRs_1_hazard_5;
  wire                _zz_DispatchPlugin_logic_rsHazardChecker_2_onLl_0_onRs_0_hazard;
  wire                _zz_DispatchPlugin_logic_rsHazardChecker_2_onLl_0_onRs_0_hazard_1;
  wire                _zz_DispatchPlugin_logic_rsHazardChecker_2_onLl_0_onRs_0_hazard_2;
  wire                _zz_DispatchPlugin_logic_rsHazardChecker_2_onLl_0_onRs_0_hazard_3;
  wire                _zz_DispatchPlugin_logic_rsHazardChecker_2_onLl_0_onRs_0_hazard_4;
  wire                _zz_DispatchPlugin_logic_rsHazardChecker_2_onLl_0_onRs_0_hazard_5;
  wire                _zz_DispatchPlugin_logic_rsHazardChecker_2_onLl_0_onRs_1_hazard;
  wire                _zz_DispatchPlugin_logic_rsHazardChecker_2_onLl_0_onRs_1_hazard_1;
  wire                _zz_DispatchPlugin_logic_rsHazardChecker_2_onLl_0_onRs_1_hazard_2;
  wire                _zz_DispatchPlugin_logic_rsHazardChecker_2_onLl_0_onRs_1_hazard_3;
  wire                _zz_DispatchPlugin_logic_rsHazardChecker_2_onLl_0_onRs_1_hazard_4;
  wire                _zz_DispatchPlugin_logic_rsHazardChecker_2_onLl_0_onRs_1_hazard_5;
  wire                _zz_DispatchPlugin_logic_rsHazardChecker_2_onLl_1_onRs_0_hazard;
  wire                _zz_DispatchPlugin_logic_rsHazardChecker_2_onLl_1_onRs_0_hazard_1;
  wire                _zz_DispatchPlugin_logic_rsHazardChecker_2_onLl_1_onRs_0_hazard_2;
  wire                _zz_DispatchPlugin_logic_rsHazardChecker_2_onLl_1_onRs_0_hazard_3;
  wire                _zz_DispatchPlugin_logic_rsHazardChecker_2_onLl_1_onRs_0_hazard_4;
  wire                _zz_DispatchPlugin_logic_rsHazardChecker_2_onLl_1_onRs_0_hazard_5;
  wire                _zz_DispatchPlugin_logic_rsHazardChecker_2_onLl_1_onRs_1_hazard;
  wire                _zz_DispatchPlugin_logic_rsHazardChecker_2_onLl_1_onRs_1_hazard_1;
  wire                _zz_DispatchPlugin_logic_rsHazardChecker_2_onLl_1_onRs_1_hazard_2;
  wire                _zz_DispatchPlugin_logic_rsHazardChecker_2_onLl_1_onRs_1_hazard_3;
  wire                _zz_DispatchPlugin_logic_rsHazardChecker_2_onLl_1_onRs_1_hazard_4;
  wire                _zz_DispatchPlugin_logic_rsHazardChecker_2_onLl_1_onRs_1_hazard_5;
  wire       [0:0]    _zz_toplevel_decode_ctrls_1_down_DispatchPlugin_logic_LANES_LAYER_HIT_0_0_2;
  wire       [0:0]    _zz_toplevel_decode_ctrls_1_down_DispatchPlugin_logic_LANES_LAYER_HIT_0_0_3;
  wire       [0:0]    _zz_toplevel_decode_ctrls_1_down_DispatchPlugin_logic_LANES_LAYER_HIT_1_0;
  wire       [0:0]    _zz_toplevel_decode_ctrls_1_down_DispatchPlugin_logic_LANES_LAYER_HIT_1_0_1;
  wire       [0:0]    _zz_toplevel_decode_ctrls_1_down_DispatchPlugin_logic_LANES_LAYER_HIT_2_0;
  wire       [0:0]    _zz_toplevel_decode_ctrls_1_down_DispatchPlugin_logic_LANES_LAYER_HIT_2_0_1;
  wire       [0:0]    _zz_toplevel_decode_ctrls_1_down_DispatchPlugin_logic_LANES_LAYER_HIT_3_0_5;
  wire       [0:0]    _zz_toplevel_decode_ctrls_1_down_DispatchPlugin_logic_LANES_LAYER_HIT_3_0_6;
  wire       [0:0]    _zz_toplevel_decode_ctrls_1_down_DispatchPlugin_MAY_FLUSH_0_1;
  wire       [0:0]    _zz_toplevel_decode_ctrls_1_down_DispatchPlugin_MAY_FLUSH_0_2;
  wire       [0:0]    _zz_toplevel_decode_ctrls_1_down_DispatchPlugin_DONT_FLUSH_0;
  wire       [0:0]    _zz_toplevel_decode_ctrls_1_down_DispatchPlugin_DONT_FLUSH_0_1;
  wire       [0:0]    _zz_toplevel_decode_ctrls_1_down_DispatchPlugin_DONT_FLUSH_FROM_LANES_0;
  wire       [0:0]    _zz_toplevel_decode_ctrls_1_down_DispatchPlugin_DONT_FLUSH_FROM_LANES_0_1;
  wire       [0:0]    _zz_toplevel_decode_ctrls_1_down_DispatchPlugin_FENCE_OLDER_0;
  wire       [0:0]    _zz_toplevel_decode_ctrls_1_down_DispatchPlugin_FENCE_OLDER_0_1;
  wire       [0:0]    _zz_toplevel_decode_ctrls_1_down_DONT_FLUSH_PRECISE_3_0;
  wire       [0:0]    _zz_toplevel_decode_ctrls_1_down_DONT_FLUSH_PRECISE_3_0_1;
  wire       [0:0]    _zz_toplevel_decode_ctrls_1_down_DONT_FLUSH_PRECISE_4_0_2;
  wire       [0:0]    _zz_toplevel_decode_ctrls_1_down_DONT_FLUSH_PRECISE_4_0_3;
  wire       [0:0]    _zz_toplevel_decode_ctrls_1_down_DecoderPlugin_logic_NEED_FPU_0;
  wire       [0:0]    _zz_toplevel_decode_ctrls_1_down_DecoderPlugin_logic_NEED_FPU_0_1;
  wire       [0:0]    _zz_toplevel_decode_ctrls_1_down_DecoderPlugin_logic_NEED_RM_0;
  wire       [0:0]    _zz_toplevel_decode_ctrls_1_down_DecoderPlugin_logic_NEED_RM_0_1;
  wire       [0:0]    _zz_toplevel_decode_ctrls_1_down_DispatchPlugin_logic_hcs_0_onRs_0_ENABLES_0_0;
  wire       [0:0]    _zz_toplevel_decode_ctrls_1_down_DispatchPlugin_logic_hcs_0_onRs_0_ENABLES_0_0_1;
  wire       [0:0]    _zz_toplevel_decode_ctrls_1_down_DispatchPlugin_logic_hcs_0_onRs_1_ENABLES_0_0;
  wire       [0:0]    _zz_toplevel_decode_ctrls_1_down_DispatchPlugin_logic_hcs_0_onRs_1_ENABLES_0_0_1;
  wire       [0:0]    _zz_toplevel_decode_ctrls_1_down_DispatchPlugin_logic_hcs_1_onRs_0_ENABLES_0_0;
  wire       [0:0]    _zz_toplevel_decode_ctrls_1_down_DispatchPlugin_logic_hcs_1_onRs_0_ENABLES_0_0_1;
  wire       [0:0]    _zz_toplevel_decode_ctrls_1_down_DispatchPlugin_logic_hcs_1_onRs_1_ENABLES_0_0_1;
  wire       [0:0]    _zz_toplevel_decode_ctrls_1_down_DispatchPlugin_logic_hcs_1_onRs_1_ENABLES_0_0_2;
  wire       [0:0]    _zz_toplevel_decode_ctrls_1_down_DispatchPlugin_logic_hcs_1_onRs_1_ENABLES_1_0;
  wire       [0:0]    _zz_toplevel_decode_ctrls_1_down_DispatchPlugin_logic_hcs_1_onRs_1_ENABLES_1_0_1;
  wire       [0:0]    _zz_toplevel_decode_ctrls_1_down_DispatchPlugin_logic_hcs_2_onRs_0_ENABLES_0_0;
  wire       [0:0]    _zz_toplevel_decode_ctrls_1_down_DispatchPlugin_logic_hcs_2_onRs_0_ENABLES_0_0_1;
  wire       [0:0]    _zz_toplevel_decode_ctrls_1_down_DispatchPlugin_logic_hcs_2_onRs_1_ENABLES_0_0;
  wire       [0:0]    _zz_toplevel_decode_ctrls_1_down_DispatchPlugin_logic_hcs_2_onRs_1_ENABLES_0_0_1;
  wire       [0:0]    _zz_toplevel_decode_ctrls_1_down_DispatchPlugin_logic_hcs_3_onRs_0_ENABLES_0_0;
  wire       [0:0]    _zz_toplevel_decode_ctrls_1_down_DispatchPlugin_logic_hcs_3_onRs_0_ENABLES_0_0_1;
  wire       [0:0]    _zz_toplevel_decode_ctrls_1_down_DispatchPlugin_logic_hcs_3_onRs_1_ENABLES_0_0_1;
  wire       [0:0]    _zz_toplevel_decode_ctrls_1_down_DispatchPlugin_logic_hcs_3_onRs_1_ENABLES_0_0_2;
  wire       [0:0]    _zz_toplevel_decode_ctrls_1_down_DispatchPlugin_logic_LANES_LAYER_HIT_0_1_2;
  wire       [0:0]    _zz_toplevel_decode_ctrls_1_down_DispatchPlugin_logic_LANES_LAYER_HIT_0_1_3;
  wire       [0:0]    _zz_toplevel_decode_ctrls_1_down_DispatchPlugin_logic_LANES_LAYER_HIT_1_1;
  wire       [0:0]    _zz_toplevel_decode_ctrls_1_down_DispatchPlugin_logic_LANES_LAYER_HIT_1_1_1;
  wire       [0:0]    _zz_toplevel_decode_ctrls_1_down_DispatchPlugin_logic_LANES_LAYER_HIT_2_1;
  wire       [0:0]    _zz_toplevel_decode_ctrls_1_down_DispatchPlugin_logic_LANES_LAYER_HIT_2_1_1;
  wire       [0:0]    _zz_toplevel_decode_ctrls_1_down_DispatchPlugin_logic_LANES_LAYER_HIT_3_1_5;
  wire       [0:0]    _zz_toplevel_decode_ctrls_1_down_DispatchPlugin_logic_LANES_LAYER_HIT_3_1_6;
  wire       [0:0]    _zz_toplevel_decode_ctrls_1_down_DispatchPlugin_MAY_FLUSH_1_1;
  wire       [0:0]    _zz_toplevel_decode_ctrls_1_down_DispatchPlugin_MAY_FLUSH_1_2;
  wire       [0:0]    _zz_toplevel_decode_ctrls_1_down_DispatchPlugin_DONT_FLUSH_1;
  wire       [0:0]    _zz_toplevel_decode_ctrls_1_down_DispatchPlugin_DONT_FLUSH_1_1;
  wire       [0:0]    _zz_toplevel_decode_ctrls_1_down_DispatchPlugin_DONT_FLUSH_FROM_LANES_1;
  wire       [0:0]    _zz_toplevel_decode_ctrls_1_down_DispatchPlugin_DONT_FLUSH_FROM_LANES_1_1;
  wire       [0:0]    _zz_toplevel_decode_ctrls_1_down_DispatchPlugin_FENCE_OLDER_1;
  wire       [0:0]    _zz_toplevel_decode_ctrls_1_down_DispatchPlugin_FENCE_OLDER_1_1;
  wire       [0:0]    _zz_toplevel_decode_ctrls_1_down_DONT_FLUSH_PRECISE_3_1;
  wire       [0:0]    _zz_toplevel_decode_ctrls_1_down_DONT_FLUSH_PRECISE_3_1_1;
  wire       [0:0]    _zz_toplevel_decode_ctrls_1_down_DONT_FLUSH_PRECISE_4_1_2;
  wire       [0:0]    _zz_toplevel_decode_ctrls_1_down_DONT_FLUSH_PRECISE_4_1_3;
  wire       [0:0]    _zz_toplevel_decode_ctrls_1_down_DecoderPlugin_logic_NEED_FPU_1;
  wire       [0:0]    _zz_toplevel_decode_ctrls_1_down_DecoderPlugin_logic_NEED_FPU_1_1;
  wire       [0:0]    _zz_toplevel_decode_ctrls_1_down_DecoderPlugin_logic_NEED_RM_1;
  wire       [0:0]    _zz_toplevel_decode_ctrls_1_down_DecoderPlugin_logic_NEED_RM_1_1;
  wire       [0:0]    _zz_toplevel_decode_ctrls_1_down_DispatchPlugin_logic_hcs_0_onRs_0_ENABLES_0_1;
  wire       [0:0]    _zz_toplevel_decode_ctrls_1_down_DispatchPlugin_logic_hcs_0_onRs_0_ENABLES_0_1_1;
  wire       [0:0]    _zz_toplevel_decode_ctrls_1_down_DispatchPlugin_logic_hcs_0_onRs_1_ENABLES_0_1;
  wire       [0:0]    _zz_toplevel_decode_ctrls_1_down_DispatchPlugin_logic_hcs_0_onRs_1_ENABLES_0_1_1;
  wire       [0:0]    _zz_toplevel_decode_ctrls_1_down_DispatchPlugin_logic_hcs_1_onRs_0_ENABLES_0_1;
  wire       [0:0]    _zz_toplevel_decode_ctrls_1_down_DispatchPlugin_logic_hcs_1_onRs_0_ENABLES_0_1_1;
  wire       [0:0]    _zz_toplevel_decode_ctrls_1_down_DispatchPlugin_logic_hcs_1_onRs_1_ENABLES_0_1_1;
  wire       [0:0]    _zz_toplevel_decode_ctrls_1_down_DispatchPlugin_logic_hcs_1_onRs_1_ENABLES_0_1_2;
  wire       [0:0]    _zz_toplevel_decode_ctrls_1_down_DispatchPlugin_logic_hcs_1_onRs_1_ENABLES_1_1;
  wire       [0:0]    _zz_toplevel_decode_ctrls_1_down_DispatchPlugin_logic_hcs_1_onRs_1_ENABLES_1_1_1;
  wire       [0:0]    _zz_toplevel_decode_ctrls_1_down_DispatchPlugin_logic_hcs_2_onRs_0_ENABLES_0_1;
  wire       [0:0]    _zz_toplevel_decode_ctrls_1_down_DispatchPlugin_logic_hcs_2_onRs_0_ENABLES_0_1_1;
  wire       [0:0]    _zz_toplevel_decode_ctrls_1_down_DispatchPlugin_logic_hcs_2_onRs_1_ENABLES_0_1;
  wire       [0:0]    _zz_toplevel_decode_ctrls_1_down_DispatchPlugin_logic_hcs_2_onRs_1_ENABLES_0_1_1;
  wire       [0:0]    _zz_toplevel_decode_ctrls_1_down_DispatchPlugin_logic_hcs_3_onRs_0_ENABLES_0_1;
  wire       [0:0]    _zz_toplevel_decode_ctrls_1_down_DispatchPlugin_logic_hcs_3_onRs_0_ENABLES_0_1_1;
  wire       [0:0]    _zz_toplevel_decode_ctrls_1_down_DispatchPlugin_logic_hcs_3_onRs_1_ENABLES_0_1_1;
  wire       [0:0]    _zz_toplevel_decode_ctrls_1_down_DispatchPlugin_logic_hcs_3_onRs_1_ENABLES_0_1_2;
  wire       [28:0]   _zz_BtbPlugin_logic_onLearn_port_payload_address_1;
  wire       [28:0]   _zz_BtbPlugin_logic_readPort_cmd_payload;
  wire       [30:0]   _zz__zz_BtbPlugin_logic_applyIt_entry_hash;
  wire       [16:0]   _zz__zz_BtbPlugin_logic_applyIt_entry_hash_1;
  wire       [30:0]   _zz__zz_BtbPlugin_logic_applyIt_entry_hash_2;
  wire       [16:0]   _zz__zz_BtbPlugin_logic_applyIt_entry_hash_3;
  wire       [31:0]   _zz_BtbPlugin_logic_ras_write_payload_data;
  wire                _zz_AlignerPlugin_logic_buffer_flushIt;
  wire                _zz_AlignerPlugin_logic_buffer_flushIt_1;
  wire       [0:0]    _zz_AlignerPlugin_logic_buffer_flushIt_2;
  wire       [1:0]    _zz_AlignerPlugin_logic_buffer_flushIt_3;
  wire                _zz_AlignerPlugin_logic_extractors_0_ctx_instruction_1;
  wire       [31:0]   _zz_AlignerPlugin_logic_extractors_0_ctx_instruction_2;
  wire                _zz_AlignerPlugin_logic_extractors_0_ctx_instruction_3;
  wire       [31:0]   _zz_AlignerPlugin_logic_extractors_0_ctx_instruction_4;
  wire                _zz_AlignerPlugin_logic_extractors_0_ctx_instruction_5;
  wire       [31:0]   _zz_AlignerPlugin_logic_extractors_0_ctx_instruction_6;
  wire                _zz_AlignerPlugin_logic_extractors_0_ctx_instruction_7;
  wire       [31:0]   _zz_AlignerPlugin_logic_extractors_0_ctx_instruction_8;
  wire                _zz_AlignerPlugin_logic_extractors_0_ctx_instruction_9;
  wire       [31:0]   _zz_AlignerPlugin_logic_extractors_0_ctx_instruction_10;
  wire                _zz_AlignerPlugin_logic_extractors_0_ctx_instruction_11;
  wire       [31:0]   _zz_AlignerPlugin_logic_extractors_0_ctx_instruction_12;
  wire                _zz_AlignerPlugin_logic_extractors_0_ctx_instruction_13;
  wire       [31:0]   _zz_AlignerPlugin_logic_extractors_0_ctx_instruction_14;
  wire                _zz_AlignerPlugin_logic_extractors_0_ctx_instruction_15;
  wire       [31:0]   _zz_AlignerPlugin_logic_extractors_0_ctx_instruction_16;
  wire                _zz_DispatchPlugin_logic_candidates_0_cancel;
  wire                _zz_DispatchPlugin_logic_candidates_0_cancel_1;
  reg        [1:0]    _zz_DispatchPlugin_logic_slotsFeeds_fit;
  wire       [1:0]    _zz_DispatchPlugin_logic_slotsFeeds_fit_1;
  wire       [0:0]    _zz__zz_DispatchPlugin_logic_slots_0_ctx_valid_4;
  wire       [141:0]  _zz__zz_DispatchPlugin_logic_slots_0_ctx_valid_4_1;
  wire       [0:0]    _zz__zz_DispatchPlugin_logic_slots_0_ctx_valid_4_2;
  wire       [135:0]  _zz__zz_DispatchPlugin_logic_slots_0_ctx_valid_4_3;
  wire       [0:0]    _zz__zz_DispatchPlugin_logic_slots_0_ctx_valid_4_4;
  wire       [116:0]  _zz__zz_DispatchPlugin_logic_slots_0_ctx_valid_4_5;
  wire       [0:0]    _zz__zz_DispatchPlugin_logic_slots_0_ctx_valid_4_6;
  wire       [64:0]   _zz__zz_DispatchPlugin_logic_slots_0_ctx_valid_4_7;
  wire       [7:0]    _zz__zz_DispatchPlugin_logic_slots_0_ctx_valid_4_8;
  wire       [40:0]   _zz__zz_DispatchPlugin_logic_slots_0_ctx_valid_4_9;
  wire       [0:0]    _zz__zz_DispatchPlugin_logic_slots_0_ctx_valid_4_10;
  wire       [0:0]    _zz__zz_DispatchPlugin_logic_slots_0_ctx_valid_4_11;
  wire       [141:0]  _zz__zz_DispatchPlugin_logic_slots_0_ctx_valid_4_12;
  wire       [0:0]    _zz__zz_DispatchPlugin_logic_slots_0_ctx_valid_4_13;
  wire       [135:0]  _zz__zz_DispatchPlugin_logic_slots_0_ctx_valid_4_14;
  wire       [0:0]    _zz__zz_DispatchPlugin_logic_slots_0_ctx_valid_4_15;
  wire       [116:0]  _zz__zz_DispatchPlugin_logic_slots_0_ctx_valid_4_16;
  wire       [0:0]    _zz__zz_DispatchPlugin_logic_slots_0_ctx_valid_4_17;
  wire       [64:0]   _zz__zz_DispatchPlugin_logic_slots_0_ctx_valid_4_18;
  wire       [7:0]    _zz__zz_DispatchPlugin_logic_slots_0_ctx_valid_4_19;
  wire       [40:0]   _zz__zz_DispatchPlugin_logic_slots_0_ctx_valid_4_20;
  wire       [0:0]    _zz__zz_DispatchPlugin_logic_slots_0_ctx_valid_4_21;
  wire       [0:0]    _zz_DispatchPlugin_logic_inserter_0_trap;
  wire       [0:0]    _zz_toplevel_execute_ctrl0_up_LANE_SEL_lane0;
  wire       [0:0]    _zz_toplevel_execute_ctrl0_up_Prediction_ALIGNED_JUMPED_lane0;
  wire       [1:0]    _zz__zz_toplevel_execute_ctrl0_up_GSharePlugin_GSHARE_COUNTER_lane0_0;
  wire       [3:0]    _zz__zz_toplevel_execute_ctrl0_up_GSharePlugin_GSHARE_COUNTER_lane0_0_1;
  wire       [1:0]    _zz__zz_toplevel_execute_ctrl0_up_GSharePlugin_GSHARE_COUNTER_lane0_0_2;
  wire       [3:0]    _zz__zz_toplevel_execute_ctrl0_up_GSharePlugin_GSHARE_COUNTER_lane0_0_3;
  wire       [1:0]    _zz__zz_toplevel_execute_ctrl0_up_GSharePlugin_GSHARE_COUNTER_lane0_0_4;
  wire       [1:0]    _zz__zz_toplevel_execute_ctrl0_up_GSharePlugin_GSHARE_COUNTER_lane0_0_5;
  wire       [0:0]    _zz_toplevel_execute_ctrl0_up_DispatchPlugin_FENCE_OLDER_lane0;
  wire       [0:0]    _zz_toplevel_execute_ctrl0_up_DispatchPlugin_MAY_FLUSH_lane0;
  wire       [0:0]    _zz_toplevel_execute_ctrl0_up_DispatchPlugin_DONT_FLUSH_lane0;
  wire       [0:0]    _zz_toplevel_execute_ctrl0_up_DispatchPlugin_DONT_FLUSH_FROM_LANES_lane0;
  wire       [0:0]    _zz_toplevel_execute_ctrl0_up_DONT_FLUSH_PRECISE_3_lane0;
  wire       [0:0]    _zz_toplevel_execute_ctrl0_up_DONT_FLUSH_PRECISE_4_lane0;
  wire       [0:0]    _zz_toplevel_execute_ctrl0_up_TRAP_lane0;
  wire       [0:0]    _zz_toplevel_execute_ctrl0_up_RS1_ENABLE_lane0;
  wire       [0:0]    _zz_toplevel_execute_ctrl0_up_RS2_ENABLE_lane0;
  wire       [0:0]    _zz_toplevel_execute_ctrl0_up_RD_ENABLE_lane0;
  wire       [0:0]    _zz_toplevel_execute_ctrl0_up_DispatchPlugin_logic_hcs_0_onRs_0_ENABLES_0_lane0;
  wire       [0:0]    _zz_toplevel_execute_ctrl0_up_DispatchPlugin_logic_hcs_0_onRs_1_ENABLES_0_lane0;
  wire       [0:0]    _zz_toplevel_execute_ctrl0_up_DispatchPlugin_logic_hcs_1_onRs_0_ENABLES_0_lane0;
  wire       [0:0]    _zz_toplevel_execute_ctrl0_up_DispatchPlugin_logic_hcs_1_onRs_1_ENABLES_0_lane0;
  wire       [0:0]    _zz_toplevel_execute_ctrl0_up_DispatchPlugin_logic_hcs_1_onRs_1_ENABLES_1_lane0;
  wire       [0:0]    _zz_toplevel_execute_ctrl0_up_DispatchPlugin_logic_hcs_2_onRs_0_ENABLES_0_lane0;
  wire       [0:0]    _zz_toplevel_execute_ctrl0_up_DispatchPlugin_logic_hcs_2_onRs_1_ENABLES_0_lane0;
  wire       [0:0]    _zz_toplevel_execute_ctrl0_up_DispatchPlugin_logic_hcs_3_onRs_0_ENABLES_0_lane0;
  wire       [0:0]    _zz_toplevel_execute_ctrl0_up_DispatchPlugin_logic_hcs_3_onRs_1_ENABLES_0_lane0;
  wire       [0:0]    _zz_DispatchPlugin_logic_inserter_1_trap;
  wire       [0:0]    _zz_toplevel_execute_ctrl0_up_LANE_SEL_lane1;
  wire       [0:0]    _zz_toplevel_execute_ctrl0_up_Prediction_ALIGNED_JUMPED_lane1;
  wire       [1:0]    _zz__zz_toplevel_execute_ctrl0_up_GSharePlugin_GSHARE_COUNTER_lane1_0;
  wire       [1:0]    _zz__zz_toplevel_execute_ctrl0_up_GSharePlugin_GSHARE_COUNTER_lane1_0_1;
  wire       [1:0]    _zz__zz_toplevel_execute_ctrl0_up_GSharePlugin_GSHARE_COUNTER_lane1_0_2;
  wire       [1:0]    _zz__zz_toplevel_execute_ctrl0_up_GSharePlugin_GSHARE_COUNTER_lane1_0_3;
  wire       [0:0]    _zz_toplevel_execute_ctrl0_up_DispatchPlugin_FENCE_OLDER_lane1;
  wire       [0:0]    _zz_toplevel_execute_ctrl0_up_DispatchPlugin_MAY_FLUSH_lane1;
  wire       [0:0]    _zz_toplevel_execute_ctrl0_up_DispatchPlugin_DONT_FLUSH_lane1;
  wire       [0:0]    _zz_toplevel_execute_ctrl0_up_DispatchPlugin_DONT_FLUSH_FROM_LANES_lane1;
  wire       [0:0]    _zz_toplevel_execute_ctrl0_up_DONT_FLUSH_PRECISE_3_lane1;
  wire       [0:0]    _zz_toplevel_execute_ctrl0_up_DONT_FLUSH_PRECISE_4_lane1;
  wire       [0:0]    _zz_toplevel_execute_ctrl0_up_TRAP_lane1;
  wire       [0:0]    _zz_toplevel_execute_ctrl0_up_RS1_ENABLE_lane1;
  wire       [0:0]    _zz_toplevel_execute_ctrl0_up_RS2_ENABLE_lane1;
  wire       [0:0]    _zz_toplevel_execute_ctrl0_up_RD_ENABLE_lane1;
  wire       [0:0]    _zz_toplevel_execute_ctrl0_up_DispatchPlugin_logic_hcs_0_onRs_0_ENABLES_0_lane1;
  wire       [0:0]    _zz_toplevel_execute_ctrl0_up_DispatchPlugin_logic_hcs_0_onRs_1_ENABLES_0_lane1;
  wire       [0:0]    _zz_toplevel_execute_ctrl0_up_DispatchPlugin_logic_hcs_1_onRs_0_ENABLES_0_lane1;
  wire       [0:0]    _zz_toplevel_execute_ctrl0_up_DispatchPlugin_logic_hcs_1_onRs_1_ENABLES_0_lane1;
  wire       [0:0]    _zz_toplevel_execute_ctrl0_up_DispatchPlugin_logic_hcs_1_onRs_1_ENABLES_1_lane1;
  wire       [0:0]    _zz_toplevel_execute_ctrl0_up_DispatchPlugin_logic_hcs_2_onRs_0_ENABLES_0_lane1;
  wire       [0:0]    _zz_toplevel_execute_ctrl0_up_DispatchPlugin_logic_hcs_2_onRs_1_ENABLES_0_lane1;
  wire       [0:0]    _zz_toplevel_execute_ctrl0_up_DispatchPlugin_logic_hcs_3_onRs_0_ENABLES_0_lane1;
  wire       [0:0]    _zz_toplevel_execute_ctrl0_up_DispatchPlugin_logic_hcs_3_onRs_1_ENABLES_0_lane1;
  wire                _zz_decode_logic_flushes_0_onLanes_0_doIt;
  wire                _zz_decode_logic_flushes_0_onLanes_0_doIt_1;
  wire       [0:0]    _zz_decode_logic_flushes_0_onLanes_0_doIt_2;
  wire       [0:0]    _zz_decode_logic_flushes_0_onLanes_0_doIt_3;
  wire                _zz_decode_logic_flushes_0_onLanes_1_doIt;
  wire                _zz_decode_logic_flushes_0_onLanes_1_doIt_1;
  wire       [0:0]    _zz_decode_logic_flushes_0_onLanes_1_doIt_2;
  wire       [0:0]    _zz_decode_logic_flushes_0_onLanes_1_doIt_3;
  wire       [0:0]    _zz_decode_logic_flushes_1_onLanes_0_doIt;
  wire                _zz_decode_logic_flushes_1_onLanes_0_doIt_1;
  wire                _zz_decode_logic_flushes_1_onLanes_0_doIt_2;
  wire                _zz_decode_logic_flushes_1_onLanes_0_doIt_3;
  wire                _zz_decode_logic_flushes_1_onLanes_0_doIt_4;
  wire                _zz_decode_logic_flushes_1_onLanes_0_doIt_5;
  wire                _zz_decode_logic_flushes_1_onLanes_0_doIt_6;
  wire       [0:0]    _zz_decode_logic_flushes_1_onLanes_0_doIt_7;
  wire       [3:0]    _zz_decode_logic_flushes_1_onLanes_0_doIt_8;
  wire                _zz_decode_logic_flushes_1_onLanes_1_doIt_1;
  wire                _zz_decode_logic_flushes_1_onLanes_1_doIt_2;
  wire                _zz_decode_logic_flushes_1_onLanes_1_doIt_3;
  wire       [0:0]    _zz_decode_logic_flushes_1_onLanes_1_doIt_4;
  wire       [2:0]    _zz_decode_logic_flushes_1_onLanes_1_doIt_5;
  wire       [21:0]   _zz_LsuL1Plugin_logic_ways_0_mem_port;
  wire                _zz_LsuL1Plugin_logic_ways_0_mem_port_1;
  wire       [21:0]   _zz_LsuL1Plugin_logic_ways_1_mem_port;
  wire                _zz_LsuL1Plugin_logic_ways_1_mem_port_1;
  wire       [2:0]    _zz_LsuL1Plugin_logic_shared_mem_port;
  wire       [0:0]    _zz_LsuL1Plugin_logic_shared_lsuRead_rsp_plru_0_1;
  wire       [2:0]    _zz_LsuL1Plugin_logic_writeback_read_wordIndex;
  wire       [0:0]    _zz_LsuL1Plugin_logic_writeback_read_wordIndex_1;
  reg        [63:0]   _zz_LsuL1Plugin_logic_writeback_read_readedData;
  wire       [2:0]    _zz_LsuL1Plugin_logic_writeback_victimBuffer_port;
  wire       [2:0]    _zz_LsuL1Plugin_logic_writeback_write_wordIndex;
  wire       [0:0]    _zz_LsuL1Plugin_logic_writeback_write_wordIndex_1;
  reg        [31:0]   _zz_toplevel_execute_ctrl3_down_LsuL1Plugin_logic_BANKS_MUXES_lane0_0;
  wire       [0:0]    _zz_toplevel_execute_ctrl3_down_LsuL1Plugin_logic_BANKS_MUXES_lane0_0_1;
  reg        [31:0]   _zz_toplevel_execute_ctrl3_down_LsuL1Plugin_logic_BANKS_MUXES_lane0_1;
  wire       [0:0]    _zz_toplevel_execute_ctrl3_down_LsuL1Plugin_logic_BANKS_MUXES_lane0_1_1;
  wire       [1:0]    _zz_LsuL1Plugin_logic_ls_ctrl_refillWayNeedWriteback;
  wire       [0:0]    _zz_LsuL1Plugin_logic_ls_ctrl_doWrite;
  reg        [1:0]    _zz_55;
  wire       [1:0]    _zz_56;
  reg        [1:0]    _zz_57;
  wire       [2:0]    _zz_58;
  wire       [1:0]    _zz_LsuL1Plugin_logic_shared_write_payload_data_dirty;
  reg        [19:0]   _zz__zz_LsuL1Plugin_logic_waysWrite_tag_address;
  reg                 _zz_LsuL1Plugin_logic_waysWrite_tag_fault;
  reg        [19:0]   _zz_LsuL1Plugin_logic_writeback_push_payload_address;
  wire       [0:0]    _zz_LsuL1Plugin_logic_shared_write_payload_data_plru_0_1;
  wire       [11:0]   _zz_LsuPlugin_logic_onAddress0_ls_storeId;
  wire       [0:0]    _zz_LsuPlugin_logic_onAddress0_ls_storeId_1;
  wire       [12:0]   _zz_LsuPlugin_logic_onAddress0_flush_port_payload_address;
  wire       [31:0]   _zz_LsuPlugin_logic_onPma_addressExtension;
  reg        [7:0]    _zz_LsuPlugin_logic_onCtrl_loadData_shited;
  wire       [1:0]    _zz_LsuPlugin_logic_onCtrl_loadData_shited_1;
  reg        [7:0]    _zz_LsuPlugin_logic_onCtrl_loadData_shited_2;
  wire       [0:0]    _zz_LsuPlugin_logic_onCtrl_loadData_shited_3;
  wire       [31:0]   _zz_LsuPlugin_logic_onCtrl_rva_alu_addSub;
  wire       [31:0]   _zz_LsuPlugin_logic_onCtrl_rva_alu_addSub_1;
  wire       [31:0]   _zz_LsuPlugin_logic_onCtrl_rva_alu_addSub_2;
  wire       [31:0]   _zz_LsuPlugin_logic_onCtrl_rva_alu_addSub_3;
  wire       [31:0]   _zz_LsuPlugin_logic_onCtrl_rva_alu_addSub_4;
  wire       [1:0]    _zz_LsuPlugin_logic_onCtrl_rva_alu_addSub_5;
  wire       [5:0]    _zz_LsuPlugin_logic_onCtrl_rva_nc_age;
  wire       [0:0]    _zz_LsuPlugin_logic_onCtrl_rva_nc_age_1;
  wire       [2:0]    _zz_LsuPlugin_logic_trapPort_payload_code;
  wire       [5:0]    _zz_LsuPlugin_logic_flusher_cmdCounter;
  reg        [2:0]    _zz_LsuL1TileLinkPlugin_logic_down_a_tracker_last;
  wire       [32:0]   _zz__zz_TrapPlugin_logic_harts_0_trap_pending_arbiter_down_payload_exception;
  wire       [32:0]   _zz__zz_TrapPlugin_logic_harts_0_trap_pending_arbiter_down_payload_exception_1;
  wire       [32:0]   _zz__zz_TrapPlugin_logic_harts_0_trap_pending_arbiter_down_payload_exception_2;
  wire       [32:0]   _zz__zz_TrapPlugin_logic_harts_0_trap_pending_arbiter_down_payload_exception_3;
  wire       [1:0]    _zz_TrapPlugin_logic_harts_0_trap_pending_slices;
  wire       [0:0]    _zz_TrapPlugin_logic_harts_0_trap_pending_slices_1;
  wire       [31:0]   _zz_TrapPlugin_logic_harts_0_trap_fsm_jumpTarget;
  wire       [2:0]    _zz_TrapPlugin_logic_harts_0_trap_fsm_jumpTarget_1;
  wire       [38:0]   _zz_FetchL1Plugin_logic_translationStorage_logic_sl_0_ways_0_port;
  wire                _zz_FetchL1Plugin_logic_translationStorage_logic_sl_0_ways_0_port_1;
  wire       [38:0]   _zz_FetchL1Plugin_logic_translationStorage_logic_sl_0_ways_1_port;
  wire                _zz_FetchL1Plugin_logic_translationStorage_logic_sl_0_ways_1_port_1;
  wire       [18:0]   _zz_FetchL1Plugin_logic_translationStorage_logic_sl_1_ways_0_port;
  wire                _zz_FetchL1Plugin_logic_translationStorage_logic_sl_1_ways_0_port_1;
  wire       [38:0]   _zz_LsuPlugin_logic_translationStorage_logic_sl_0_ways_0_port;
  wire                _zz_LsuPlugin_logic_translationStorage_logic_sl_0_ways_0_port_1;
  wire       [38:0]   _zz_LsuPlugin_logic_translationStorage_logic_sl_0_ways_1_port;
  wire                _zz_LsuPlugin_logic_translationStorage_logic_sl_0_ways_1_port_1;
  wire       [18:0]   _zz_LsuPlugin_logic_translationStorage_logic_sl_1_ways_0_port;
  wire                _zz_LsuPlugin_logic_translationStorage_logic_sl_1_ways_0_port_1;
  wire       [0:0]    _zz_LsuPlugin_logic_onAddress0_translationPort_logic_ctrl_lineAllowExecute_3;
  wire       [0:0]    _zz_LsuPlugin_logic_onAddress0_translationPort_logic_ctrl_lineAllowRead;
  wire       [0:0]    _zz_LsuPlugin_logic_onAddress0_translationPort_logic_ctrl_lineAllowWrite;
  wire       [0:0]    _zz_LsuPlugin_logic_onAddress0_translationPort_logic_ctrl_lineAllowUser;
  wire       [11:0]   _zz_LsuPlugin_logic_onAddress0_translationPort_logic_ctrl_lineTranslated;
  wire       [11:0]   _zz_LsuPlugin_logic_onAddress0_translationPort_logic_ctrl_lineTranslated_1;
  wire       [0:0]    _zz_FetchL1Plugin_logic_translationPort_logic_ctrl_lineAllowExecute_3;
  wire       [0:0]    _zz_FetchL1Plugin_logic_translationPort_logic_ctrl_lineAllowRead;
  wire       [0:0]    _zz_FetchL1Plugin_logic_translationPort_logic_ctrl_lineAllowWrite;
  wire       [0:0]    _zz_FetchL1Plugin_logic_translationPort_logic_ctrl_lineAllowUser;
  wire       [11:0]   _zz_FetchL1Plugin_logic_translationPort_logic_ctrl_lineTranslated;
  wire       [11:0]   _zz_FetchL1Plugin_logic_translationPort_logic_ctrl_lineTranslated_1;
  wire       [31:0]   _zz_PcPlugin_logic_harts_0_self_pc;
  wire       [3:0]    _zz_PcPlugin_logic_harts_0_self_pc_1;
  wire       [31:0]   _zz_PcPlugin_logic_harts_0_aggregator_target_7;
  wire       [31:0]   _zz_PcPlugin_logic_harts_0_aggregator_target_8;
  wire       [31:0]   _zz_PcPlugin_logic_harts_0_aggregator_target_9;
  wire       [31:0]   _zz_PcPlugin_logic_harts_0_aggregator_target_10;
  wire       [31:0]   _zz_PcPlugin_logic_harts_0_aggregator_target_11;
  wire       [31:0]   _zz_PcPlugin_logic_harts_0_aggregator_target_12;
  wire       [31:0]   _zz_PcPlugin_logic_harts_0_aggregator_target_13;
  wire       [31:0]   _zz_PcPlugin_logic_harts_0_aggregator_target_14;
  wire       [31:0]   _zz_PcPlugin_logic_harts_0_aggregator_target_15;
  wire       [31:0]   _zz_PcPlugin_logic_harts_0_aggregator_target_16;
  wire       [31:0]   _zz_PcPlugin_logic_harts_0_aggregator_target_17;
  wire       [31:0]   _zz_PcPlugin_logic_harts_0_aggregator_target_18;
  wire       [0:0]    _zz_PcPlugin_logic_harts_0_aggregator_fault;
  wire       [11:0]   _zz_COMB_CSR_CsrRamPlugin_csrMapper_selFilter;
  wire                _zz_COMB_CSR_CsrRamPlugin_csrMapper_selFilter_1;
  wire       [0:0]    _zz_COMB_CSR_CsrRamPlugin_csrMapper_selFilter_2;
  wire       [0:0]    _zz_COMB_CSR_CsrRamPlugin_csrMapper_selFilter_3;
  wire       [0:0]    _zz_CsrAccessPlugin_logic_fsm_inject_implemented;
  wire       [13:0]   _zz_CsrAccessPlugin_logic_fsm_inject_implemented_1;
  wire       [0:0]    _zz_CsrAccessPlugin_logic_fsm_inject_implemented_2;
  wire       [2:0]    _zz_CsrAccessPlugin_logic_fsm_inject_implemented_3;
  wire       [31:0]   _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_13;
  wire       [31:0]   _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_14;
  wire       [5:0]    _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_15;
  wire       [31:0]   _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_16;
  wire       [31:0]   _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_17;
  wire       [31:0]   _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_18;
  wire       [7:0]    _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_19;
  wire       [31:0]   _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_20;
  wire       [31:0]   _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_21;
  wire       [3:0]    _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_22;
  wire       [31:0]   _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_23;
  wire       [12:0]   _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_24;
  wire       [31:0]   _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_25;
  wire       [31:0]   _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_26;
  wire       [31:0]   _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_27;
  wire       [14:0]   _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_28;
  wire       [31:0]   _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_29;
  wire       [31:0]   _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_30;
  wire       [22:0]   _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_31;
  wire       [31:0]   _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_32;
  wire       [20:0]   _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_33;
  wire       [31:0]   _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_34;
  wire       [31:0]   _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_35;
  wire       [21:0]   _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_36;
  wire       [31:0]   _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_37;
  wire       [31:0]   _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_38;
  wire       [31:0]   _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_39;
  wire       [3:0]    _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_40;
  wire       [31:0]   _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_41;
  wire       [11:0]   _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_42;
  wire       [31:0]   _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_43;
  wire       [31:0]   _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_44;
  wire       [7:0]    _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_45;
  wire       [31:0]   _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_46;
  wire       [3:0]    _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_47;
  wire       [31:0]   _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_48;
  wire       [31:0]   _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_49;
  wire       [11:0]   _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_50;
  wire       [31:0]   _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_51;
  wire       [7:0]    _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_52;
  wire       [31:0]   _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_53;
  wire       [31:0]   _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_54;
  wire       [3:0]    _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_55;
  wire       [31:0]   _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_56;
  wire       [0:0]    _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_57;
  wire       [31:0]   _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_58;
  wire       [31:0]   _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_59;
  wire       [3:0]    _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_60;
  wire       [31:0]   _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_61;
  wire       [8:0]    _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_62;
  wire       [31:0]   _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_63;
  wire       [31:0]   _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_64;
  wire       [9:0]    _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_65;
  wire       [31:0]   _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_66;
  wire       [12:0]   _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_67;
  wire       [31:0]   _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_68;
  wire       [31:0]   _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_69;
  wire       [13:0]   _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_70;
  wire       [31:0]   _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_71;
  wire       [15:0]   _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_72;
  wire       [31:0]   _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_73;
  wire       [31:0]   _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_74;
  wire       [9:0]    _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_75;
  wire       [31:0]   _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_76;
  wire       [5:0]    _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_77;
  wire       [31:0]   _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_78;
  wire       [31:0]   _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_79;
  wire       [1:0]    _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_80;
  wire       [31:0]   _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_81;
  wire       [31:0]   _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_82;
  wire       [31:0]   _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_83;
  wire       [3:0]    _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_84;
  wire       [31:0]   _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_85;
  wire       [31:0]   _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_86;
  wire       [31:0]   _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_87;
  wire       [8:0]    _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_88;
  wire       [31:0]   _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_89;
  wire       [5:0]    _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_90;
  wire       [31:0]   _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_91;
  wire       [31:0]   _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_92;
  wire       [1:0]    _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_93;
  wire       [31:0]   _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_94;
  wire       [8:0]    _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_95;
  wire       [31:0]   _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_96;
  wire       [31:0]   _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_97;
  wire       [5:0]    _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_98;
  wire       [31:0]   _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_99;
  wire       [1:0]    _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_100;
  wire       [31:0]   _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_101;
  wire       [31:0]   _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_102;
  wire       [14:0]   _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_103;
  wire       [31:0]   _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_104;
  wire       [9:0]    _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_105;
  wire       [31:0]   _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_106;
  wire       [31:0]   _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_107;
  wire       [9:0]    _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_108;
  wire       [31:0]   _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_109;
  wire       [5:0]    _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_110;
  wire       [31:0]   _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_111;
  wire       [31:0]   _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_112;
  wire       [5:0]    _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_113;
  wire       [31:0]   _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_114;
  wire       [1:0]    _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_115;
  wire       [31:0]   _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_116;
  wire       [31:0]   _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_117;
  wire       [1:0]    _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_118;
  wire       [31:0]   _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_119;
  wire       [9:0]    _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_120;
  wire       [31:0]   _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_121;
  wire       [31:0]   _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_122;
  wire       [9:0]    _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_123;
  wire       [31:0]   _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_124;
  wire       [5:0]    _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_125;
  wire       [31:0]   _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_126;
  wire       [31:0]   _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_127;
  wire       [5:0]    _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_128;
  wire       [31:0]   _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_129;
  wire       [1:0]    _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_130;
  wire       [31:0]   _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_131;
  wire       [31:0]   _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_132;
  wire       [1:0]    _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_133;
  wire       [31:0]   _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_134;
  wire       [31:0]   _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_135;
  wire       [19:0]   _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_136;
  wire       [31:0]   _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_137;
  wire       [31:0]   _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_138;
  wire       [18:0]   _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_139;
  wire       [31:0]   _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_140;
  wire       [19:0]   _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_141;
  wire       [31:0]   _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_142;
  wire       [31:0]   _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_143;
  wire       [18:0]   _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_144;
  wire       [31:0]   _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_145;
  wire       [17:0]   _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_146;
  wire       [31:0]   _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_147;
  wire       [31:0]   _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_148;
  wire       [31:0]   _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_149;
  wire       [19:0]   _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_150;
  wire       [31:0]   _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_151;
  wire       [31:0]   _zz_CsrAccessPlugin_logic_fsm_writeLogic_alu_mask;
  wire       [4:0]    _zz_CsrAccessPlugin_logic_fsm_writeLogic_alu_mask_1;
  wire       [2:0]    _zz_CsrRamPlugin_logic_writeLogic_hits_ohFirst_masked;
  wire       [1:0]    _zz_CsrRamPlugin_logic_readLogic_hits_ohFirst_masked;
  reg        [2:0]    _zz_CsrRamPlugin_logic_readLogic_port_cmd_payload;
  wire       [3:0]    _zz_CsrRamPlugin_logic_flush_counter;
  wire       [0:0]    _zz_CsrRamPlugin_logic_flush_counter_1;
  wire                _zz__zz_toplevel_execute_ctrl1_down_integer_RS1_lane0_1;
  wire       [31:0]   _zz__zz_toplevel_execute_ctrl1_down_integer_RS1_lane0_1_1;
  wire                _zz__zz_toplevel_execute_ctrl1_down_integer_RS1_lane0_1_2;
  wire       [31:0]   _zz__zz_toplevel_execute_ctrl1_down_integer_RS1_lane0_1_3;
  wire                _zz__zz_toplevel_execute_ctrl1_down_integer_RS1_lane0_1_4;
  wire       [31:0]   _zz__zz_toplevel_execute_ctrl1_down_integer_RS1_lane0_1_5;
  wire                _zz__zz_toplevel_execute_ctrl1_down_integer_RS1_lane0_1_6;
  wire       [31:0]   _zz__zz_toplevel_execute_ctrl1_down_integer_RS1_lane0_1_7;
  wire                _zz__zz_toplevel_execute_ctrl1_down_integer_RS1_lane0_1_8;
  wire       [31:0]   _zz__zz_toplevel_execute_ctrl1_down_integer_RS1_lane0_1_9;
  wire                _zz__zz_toplevel_execute_ctrl1_down_integer_RS1_lane0_1_10;
  wire       [31:0]   _zz__zz_toplevel_execute_ctrl1_down_integer_RS1_lane0_1_11;
  wire                _zz__zz_toplevel_execute_ctrl1_down_integer_RS1_lane0_1_12;
  wire       [31:0]   _zz__zz_toplevel_execute_ctrl1_down_integer_RS1_lane0_1_13;
  wire                _zz__zz_toplevel_execute_ctrl1_down_integer_RS1_lane0_1_14;
  wire       [31:0]   _zz__zz_toplevel_execute_ctrl1_down_integer_RS1_lane0_1_15;
  wire                _zz__zz_toplevel_execute_ctrl1_down_integer_RS2_lane0_1;
  wire       [31:0]   _zz__zz_toplevel_execute_ctrl1_down_integer_RS2_lane0_1_1;
  wire                _zz__zz_toplevel_execute_ctrl1_down_integer_RS2_lane0_1_2;
  wire       [31:0]   _zz__zz_toplevel_execute_ctrl1_down_integer_RS2_lane0_1_3;
  wire                _zz__zz_toplevel_execute_ctrl1_down_integer_RS2_lane0_1_4;
  wire       [31:0]   _zz__zz_toplevel_execute_ctrl1_down_integer_RS2_lane0_1_5;
  wire                _zz__zz_toplevel_execute_ctrl1_down_integer_RS2_lane0_1_6;
  wire       [31:0]   _zz__zz_toplevel_execute_ctrl1_down_integer_RS2_lane0_1_7;
  wire                _zz__zz_toplevel_execute_ctrl1_down_integer_RS2_lane0_1_8;
  wire       [31:0]   _zz__zz_toplevel_execute_ctrl1_down_integer_RS2_lane0_1_9;
  wire                _zz__zz_toplevel_execute_ctrl1_down_integer_RS2_lane0_1_10;
  wire       [31:0]   _zz__zz_toplevel_execute_ctrl1_down_integer_RS2_lane0_1_11;
  wire                _zz__zz_toplevel_execute_ctrl1_down_integer_RS2_lane0_1_12;
  wire       [31:0]   _zz__zz_toplevel_execute_ctrl1_down_integer_RS2_lane0_1_13;
  wire                _zz__zz_toplevel_execute_ctrl1_down_integer_RS2_lane0_1_14;
  wire       [31:0]   _zz__zz_toplevel_execute_ctrl1_down_integer_RS2_lane0_1_15;
  wire       [0:0]    _zz_toplevel_execute_ctrl1_down_early0_IntAluPlugin_SEL_lane0;
  wire       [0:0]    _zz_toplevel_execute_ctrl1_down_early0_IntAluPlugin_SEL_lane0_1;
  wire       [0:0]    _zz_toplevel_execute_ctrl1_down_early0_BarrelShifterPlugin_SEL_lane0;
  wire       [0:0]    _zz_toplevel_execute_ctrl1_down_early0_BarrelShifterPlugin_SEL_lane0_1;
  wire       [0:0]    _zz_toplevel_execute_ctrl1_down_early0_BranchPlugin_SEL_lane0;
  wire       [0:0]    _zz_toplevel_execute_ctrl1_down_early0_BranchPlugin_SEL_lane0_1;
  wire       [0:0]    _zz_toplevel_execute_ctrl1_down_early0_MulPlugin_SEL_lane0;
  wire       [0:0]    _zz_toplevel_execute_ctrl1_down_early0_MulPlugin_SEL_lane0_1;
  wire       [0:0]    _zz_toplevel_execute_ctrl1_down_early0_DivPlugin_SEL_lane0;
  wire       [0:0]    _zz_toplevel_execute_ctrl1_down_early0_DivPlugin_SEL_lane0_1;
  wire       [0:0]    _zz_toplevel_execute_ctrl1_down_early0_EnvPlugin_SEL_lane0;
  wire       [0:0]    _zz_toplevel_execute_ctrl1_down_early0_EnvPlugin_SEL_lane0_1;
  wire       [0:0]    _zz_toplevel_execute_ctrl1_down_late0_IntAluPlugin_SEL_lane0;
  wire       [0:0]    _zz_toplevel_execute_ctrl1_down_late0_IntAluPlugin_SEL_lane0_1;
  wire       [0:0]    _zz_toplevel_execute_ctrl1_down_late0_BarrelShifterPlugin_SEL_lane0;
  wire       [0:0]    _zz_toplevel_execute_ctrl1_down_late0_BarrelShifterPlugin_SEL_lane0_1;
  wire       [0:0]    _zz_toplevel_execute_ctrl1_down_late0_BranchPlugin_SEL_lane0_1;
  wire       [0:0]    _zz_toplevel_execute_ctrl1_down_late0_BranchPlugin_SEL_lane0_2;
  wire       [0:0]    _zz_toplevel_execute_ctrl1_down_MulPlugin_HIGH_lane0;
  wire       [0:0]    _zz_toplevel_execute_ctrl1_down_MulPlugin_HIGH_lane0_1;
  wire       [0:0]    _zz_toplevel_execute_ctrl1_down_CsrAccessPlugin_SEL_lane0;
  wire       [0:0]    _zz_toplevel_execute_ctrl1_down_CsrAccessPlugin_SEL_lane0_1;
  wire       [0:0]    _zz_toplevel_execute_ctrl1_down_AguPlugin_SEL_lane0;
  wire       [0:0]    _zz_toplevel_execute_ctrl1_down_AguPlugin_SEL_lane0_1;
  wire       [0:0]    _zz_toplevel_execute_ctrl1_down_LsuPlugin_logic_FENCE_lane0;
  wire       [0:0]    _zz_toplevel_execute_ctrl1_down_LsuPlugin_logic_FENCE_lane0_1;
  wire       [0:0]    _zz_toplevel_execute_ctrl1_down_lane0_integer_WriteBackPlugin_SEL_lane0_1;
  wire       [0:0]    _zz_toplevel_execute_ctrl1_down_lane0_integer_WriteBackPlugin_SEL_lane0_2;
  wire       [32:0]   _zz_toplevel_execute_ctrl1_down_lane0_integer_WriteBackPlugin_SEL_lane0_3;
  wire       [32:0]   _zz_toplevel_execute_ctrl1_down_lane0_integer_WriteBackPlugin_SEL_lane0_4;
  wire       [0:0]    _zz_toplevel_execute_ctrl1_down_COMPLETION_AT_2_lane0;
  wire       [0:0]    _zz_toplevel_execute_ctrl1_down_COMPLETION_AT_2_lane0_1;
  wire       [0:0]    _zz_toplevel_execute_ctrl1_down_COMPLETION_AT_3_lane0;
  wire       [0:0]    _zz_toplevel_execute_ctrl1_down_COMPLETION_AT_3_lane0_1;
  wire       [0:0]    _zz_toplevel_execute_ctrl1_down_COMPLETION_AT_4_lane0;
  wire       [0:0]    _zz_toplevel_execute_ctrl1_down_COMPLETION_AT_4_lane0_1;
  wire       [0:0]    _zz_toplevel_execute_ctrl1_down_execute_lane0_logic_completions_onCtrl_0_ENABLE_lane0_7;
  wire       [0:0]    _zz_toplevel_execute_ctrl1_down_execute_lane0_logic_completions_onCtrl_0_ENABLE_lane0_8;
  wire       [0:0]    _zz_toplevel_execute_ctrl1_down_execute_lane0_logic_completions_onCtrl_1_ENABLE_lane0_6;
  wire       [0:0]    _zz_toplevel_execute_ctrl1_down_execute_lane0_logic_completions_onCtrl_1_ENABLE_lane0_7;
  wire       [0:0]    _zz_toplevel_execute_ctrl1_down_execute_lane0_logic_completions_onCtrl_2_ENABLE_lane0_4;
  wire       [0:0]    _zz_toplevel_execute_ctrl1_down_execute_lane0_logic_completions_onCtrl_2_ENABLE_lane0_5;
  wire       [0:0]    _zz_toplevel_execute_ctrl1_down_early0_IntAluPlugin_ALU_ADD_SUB_lane0;
  wire       [0:0]    _zz_toplevel_execute_ctrl1_down_early0_IntAluPlugin_ALU_ADD_SUB_lane0_1;
  wire       [0:0]    _zz_toplevel_execute_ctrl1_down_early0_IntAluPlugin_ALU_SLTX_lane0;
  wire       [0:0]    _zz_toplevel_execute_ctrl1_down_early0_IntAluPlugin_ALU_SLTX_lane0_1;
  wire       [0:0]    _zz_toplevel_execute_ctrl1_down_SrcStageables_REVERT_lane0;
  wire       [0:0]    _zz_toplevel_execute_ctrl1_down_SrcStageables_REVERT_lane0_1;
  wire       [0:0]    _zz_toplevel_execute_ctrl1_down_SrcStageables_ZERO_lane0;
  wire       [0:0]    _zz_toplevel_execute_ctrl1_down_SrcStageables_ZERO_lane0_1;
  wire       [0:0]    _zz_toplevel_execute_ctrl1_down_lane0_IntFormatPlugin_logic_SIGNED_lane0;
  wire       [0:0]    _zz_toplevel_execute_ctrl1_down_lane0_IntFormatPlugin_logic_SIGNED_lane0_1;
  wire       [32:0]   _zz_toplevel_execute_ctrl1_down_lane0_IntFormatPlugin_logic_WIDTH_ID_lane0;
  wire       [32:0]   _zz_toplevel_execute_ctrl1_down_lane0_IntFormatPlugin_logic_WIDTH_ID_lane0_1;
  wire       [32:0]   _zz_toplevel_execute_ctrl1_down_lane0_IntFormatPlugin_logic_WIDTH_ID_lane0_2;
  wire       [0:0]    _zz_toplevel_execute_ctrl1_down_BYPASSED_AT_2_lane0;
  wire       [0:0]    _zz_toplevel_execute_ctrl1_down_BYPASSED_AT_2_lane0_1;
  wire       [0:0]    _zz_toplevel_execute_ctrl1_down_BYPASSED_AT_3_lane0_1;
  wire       [0:0]    _zz_toplevel_execute_ctrl1_down_BYPASSED_AT_3_lane0_2;
  wire       [0:0]    _zz_toplevel_execute_ctrl1_down_MAY_FLUSH_PRECISE_3_lane0;
  wire       [0:0]    _zz_toplevel_execute_ctrl1_down_MAY_FLUSH_PRECISE_3_lane0_1;
  wire       [0:0]    _zz_toplevel_execute_ctrl1_down_MAY_FLUSH_PRECISE_4_lane0;
  wire       [0:0]    _zz_toplevel_execute_ctrl1_down_MAY_FLUSH_PRECISE_4_lane0_1;
  wire       [0:0]    _zz_toplevel_execute_ctrl1_down_SrcStageables_UNSIGNED_lane0_1;
  wire       [0:0]    _zz_toplevel_execute_ctrl1_down_SrcStageables_UNSIGNED_lane0_2;
  wire       [0:0]    _zz_toplevel_execute_ctrl1_down_BarrelShifterPlugin_LEFT_lane0_1;
  wire       [0:0]    _zz_toplevel_execute_ctrl1_down_BarrelShifterPlugin_LEFT_lane0_2;
  wire       [0:0]    _zz_toplevel_execute_ctrl1_down_BarrelShifterPlugin_SIGNED_lane0;
  wire       [0:0]    _zz_toplevel_execute_ctrl1_down_BarrelShifterPlugin_SIGNED_lane0_1;
  wire       [0:0]    _zz_toplevel_execute_ctrl1_down_RsUnsignedPlugin_RS1_SIGNED_lane0;
  wire       [0:0]    _zz_toplevel_execute_ctrl1_down_RsUnsignedPlugin_RS1_SIGNED_lane0_1;
  wire       [0:0]    _zz_toplevel_execute_ctrl1_down_RsUnsignedPlugin_RS2_SIGNED_lane0;
  wire       [0:0]    _zz_toplevel_execute_ctrl1_down_RsUnsignedPlugin_RS2_SIGNED_lane0_1;
  wire       [0:0]    _zz_toplevel_execute_ctrl1_down_DivPlugin_REM_lane0;
  wire       [0:0]    _zz_toplevel_execute_ctrl1_down_DivPlugin_REM_lane0_1;
  wire       [0:0]    _zz_toplevel_execute_ctrl1_down_CsrAccessPlugin_CSR_IMM_lane0;
  wire       [0:0]    _zz_toplevel_execute_ctrl1_down_CsrAccessPlugin_CSR_IMM_lane0_1;
  wire       [0:0]    _zz_toplevel_execute_ctrl1_down_CsrAccessPlugin_CSR_MASK_lane0_1;
  wire       [0:0]    _zz_toplevel_execute_ctrl1_down_CsrAccessPlugin_CSR_MASK_lane0_2;
  wire       [0:0]    _zz_toplevel_execute_ctrl1_down_CsrAccessPlugin_CSR_CLEAR_lane0_1;
  wire       [0:0]    _zz_toplevel_execute_ctrl1_down_CsrAccessPlugin_CSR_CLEAR_lane0_2;
  wire       [0:0]    _zz_toplevel_execute_ctrl1_down_AguPlugin_LOAD_lane0_1;
  wire       [0:0]    _zz_toplevel_execute_ctrl1_down_AguPlugin_LOAD_lane0_2;
  wire       [0:0]    _zz_toplevel_execute_ctrl1_down_AguPlugin_STORE_lane0_1;
  wire       [0:0]    _zz_toplevel_execute_ctrl1_down_AguPlugin_STORE_lane0_2;
  wire       [0:0]    _zz_toplevel_execute_ctrl1_down_AguPlugin_ATOMIC_lane0_1;
  wire       [0:0]    _zz_toplevel_execute_ctrl1_down_AguPlugin_ATOMIC_lane0_2;
  wire       [0:0]    _zz_toplevel_execute_ctrl1_down_AguPlugin_FLOAT_lane0;
  wire       [0:0]    _zz_toplevel_execute_ctrl1_down_AguPlugin_FLOAT_lane0_1;
  wire       [0:0]    _zz_toplevel_execute_ctrl1_down_LsuPlugin_logic_LSU_PREFETCH_lane0;
  wire       [0:0]    _zz_toplevel_execute_ctrl1_down_LsuPlugin_logic_LSU_PREFETCH_lane0_1;
  wire       [32:0]   _zz__zz_toplevel_execute_ctrl1_down_early0_EnvPlugin_OP_lane0_2;
  wire       [32:0]   _zz__zz_toplevel_execute_ctrl1_down_early0_EnvPlugin_OP_lane0_2_1;
  wire       [32:0]   _zz__zz_toplevel_execute_ctrl1_down_early0_EnvPlugin_OP_lane0_2_2;
  wire       [32:0]   _zz__zz_toplevel_execute_ctrl1_down_early0_EnvPlugin_OP_lane0_2_3;
  wire                _zz__zz_toplevel_execute_ctrl1_down_early0_EnvPlugin_OP_lane0_2_4;
  wire                _zz__zz_toplevel_execute_ctrl1_down_early0_EnvPlugin_OP_lane0_2_5;
  wire       [0:0]    _zz_toplevel_execute_ctrl1_down_late0_IntAluPlugin_ALU_ADD_SUB_lane0_1;
  wire       [0:0]    _zz_toplevel_execute_ctrl1_down_late0_IntAluPlugin_ALU_ADD_SUB_lane0_2;
  wire       [0:0]    _zz_toplevel_execute_ctrl1_down_late0_IntAluPlugin_ALU_SLTX_lane0_1;
  wire       [0:0]    _zz_toplevel_execute_ctrl1_down_late0_IntAluPlugin_ALU_SLTX_lane0_2;
  wire                _zz_when_ExecuteLanePlugin_l300_2;
  wire                _zz_when_ExecuteLanePlugin_l300_2_1;
  wire                _zz_when_ExecuteLanePlugin_l300_2_2;
  wire                _zz_when_ExecuteLanePlugin_l300_2_3;
  wire                _zz_when_ExecuteLanePlugin_l300_2_4;
  wire                _zz_when_ExecuteLanePlugin_l300_2_5;
  wire                _zz_when_ExecuteLanePlugin_l300_3;
  wire                _zz_when_ExecuteLanePlugin_l300_3_1;
  wire                _zz_when_ExecuteLanePlugin_l300_3_2;
  wire                _zz_when_ExecuteLanePlugin_l300_4;
  wire                _zz_when_ExecuteLanePlugin_l300_4_1;
  wire       [31:0]   _zz_WhiteboxerPlugin_logic_csr_access_payload_address;
  wire                _zz_fetch_logic_flushes_0_doIt;
  wire                _zz_fetch_logic_flushes_0_doIt_1;
  wire       [0:0]    _zz_fetch_logic_flushes_0_doIt_2;
  wire       [1:0]    _zz_fetch_logic_flushes_0_doIt_3;
  wire                _zz_fetch_logic_flushes_1_doIt;
  wire                _zz_fetch_logic_flushes_1_doIt_1;
  wire       [0:0]    _zz_fetch_logic_flushes_1_doIt_2;
  wire       [1:0]    _zz_fetch_logic_flushes_1_doIt_3;
  wire                _zz__zz_toplevel_execute_ctrl1_down_integer_RS1_lane1_1;
  wire       [31:0]   _zz__zz_toplevel_execute_ctrl1_down_integer_RS1_lane1_1_1;
  wire                _zz__zz_toplevel_execute_ctrl1_down_integer_RS1_lane1_1_2;
  wire       [31:0]   _zz__zz_toplevel_execute_ctrl1_down_integer_RS1_lane1_1_3;
  wire                _zz__zz_toplevel_execute_ctrl1_down_integer_RS1_lane1_1_4;
  wire       [31:0]   _zz__zz_toplevel_execute_ctrl1_down_integer_RS1_lane1_1_5;
  wire                _zz__zz_toplevel_execute_ctrl1_down_integer_RS1_lane1_1_6;
  wire       [31:0]   _zz__zz_toplevel_execute_ctrl1_down_integer_RS1_lane1_1_7;
  wire                _zz__zz_toplevel_execute_ctrl1_down_integer_RS1_lane1_1_8;
  wire       [31:0]   _zz__zz_toplevel_execute_ctrl1_down_integer_RS1_lane1_1_9;
  wire                _zz__zz_toplevel_execute_ctrl1_down_integer_RS1_lane1_1_10;
  wire       [31:0]   _zz__zz_toplevel_execute_ctrl1_down_integer_RS1_lane1_1_11;
  wire                _zz__zz_toplevel_execute_ctrl1_down_integer_RS1_lane1_1_12;
  wire       [31:0]   _zz__zz_toplevel_execute_ctrl1_down_integer_RS1_lane1_1_13;
  wire                _zz__zz_toplevel_execute_ctrl1_down_integer_RS1_lane1_1_14;
  wire       [31:0]   _zz__zz_toplevel_execute_ctrl1_down_integer_RS1_lane1_1_15;
  wire                _zz__zz_toplevel_execute_ctrl1_down_integer_RS2_lane1_1;
  wire       [31:0]   _zz__zz_toplevel_execute_ctrl1_down_integer_RS2_lane1_1_1;
  wire                _zz__zz_toplevel_execute_ctrl1_down_integer_RS2_lane1_1_2;
  wire       [31:0]   _zz__zz_toplevel_execute_ctrl1_down_integer_RS2_lane1_1_3;
  wire                _zz__zz_toplevel_execute_ctrl1_down_integer_RS2_lane1_1_4;
  wire       [31:0]   _zz__zz_toplevel_execute_ctrl1_down_integer_RS2_lane1_1_5;
  wire                _zz__zz_toplevel_execute_ctrl1_down_integer_RS2_lane1_1_6;
  wire       [31:0]   _zz__zz_toplevel_execute_ctrl1_down_integer_RS2_lane1_1_7;
  wire                _zz__zz_toplevel_execute_ctrl1_down_integer_RS2_lane1_1_8;
  wire       [31:0]   _zz__zz_toplevel_execute_ctrl1_down_integer_RS2_lane1_1_9;
  wire                _zz__zz_toplevel_execute_ctrl1_down_integer_RS2_lane1_1_10;
  wire       [31:0]   _zz__zz_toplevel_execute_ctrl1_down_integer_RS2_lane1_1_11;
  wire                _zz__zz_toplevel_execute_ctrl1_down_integer_RS2_lane1_1_12;
  wire       [31:0]   _zz__zz_toplevel_execute_ctrl1_down_integer_RS2_lane1_1_13;
  wire                _zz__zz_toplevel_execute_ctrl1_down_integer_RS2_lane1_1_14;
  wire       [31:0]   _zz__zz_toplevel_execute_ctrl1_down_integer_RS2_lane1_1_15;
  wire       [0:0]    _zz_toplevel_execute_ctrl1_down_early1_IntAluPlugin_SEL_lane1;
  wire       [0:0]    _zz_toplevel_execute_ctrl1_down_early1_IntAluPlugin_SEL_lane1_1;
  wire       [0:0]    _zz_toplevel_execute_ctrl1_down_early1_BarrelShifterPlugin_SEL_lane1;
  wire       [0:0]    _zz_toplevel_execute_ctrl1_down_early1_BarrelShifterPlugin_SEL_lane1_1;
  wire       [0:0]    _zz_toplevel_execute_ctrl1_down_early1_BranchPlugin_SEL_lane1;
  wire       [0:0]    _zz_toplevel_execute_ctrl1_down_early1_BranchPlugin_SEL_lane1_1;
  wire       [0:0]    _zz_toplevel_execute_ctrl1_down_late1_IntAluPlugin_SEL_lane1;
  wire       [0:0]    _zz_toplevel_execute_ctrl1_down_late1_IntAluPlugin_SEL_lane1_1;
  wire       [0:0]    _zz_toplevel_execute_ctrl1_down_late1_BarrelShifterPlugin_SEL_lane1;
  wire       [0:0]    _zz_toplevel_execute_ctrl1_down_late1_BarrelShifterPlugin_SEL_lane1_1;
  wire       [0:0]    _zz_toplevel_execute_ctrl1_down_late1_BranchPlugin_SEL_lane1_1;
  wire       [0:0]    _zz_toplevel_execute_ctrl1_down_late1_BranchPlugin_SEL_lane1_2;
  wire       [0:0]    _zz_toplevel_execute_ctrl1_down_lane1_integer_WriteBackPlugin_SEL_lane1;
  wire       [0:0]    _zz_toplevel_execute_ctrl1_down_lane1_integer_WriteBackPlugin_SEL_lane1_1;
  wire       [0:0]    _zz_toplevel_execute_ctrl1_down_COMPLETION_AT_2_lane1;
  wire       [0:0]    _zz_toplevel_execute_ctrl1_down_COMPLETION_AT_2_lane1_1;
  wire       [0:0]    _zz_toplevel_execute_ctrl1_down_COMPLETION_AT_3_lane1;
  wire       [0:0]    _zz_toplevel_execute_ctrl1_down_COMPLETION_AT_3_lane1_1;
  wire       [0:0]    _zz_toplevel_execute_ctrl1_down_COMPLETION_AT_4_lane1;
  wire       [0:0]    _zz_toplevel_execute_ctrl1_down_COMPLETION_AT_4_lane1_1;
  wire       [0:0]    _zz_toplevel_execute_ctrl1_down_execute_lane1_logic_completions_onCtrl_0_ENABLE_lane1_3;
  wire       [0:0]    _zz_toplevel_execute_ctrl1_down_execute_lane1_logic_completions_onCtrl_0_ENABLE_lane1_4;
  wire       [0:0]    _zz_toplevel_execute_ctrl1_down_execute_lane1_logic_completions_onCtrl_1_ENABLE_lane1_2;
  wire       [0:0]    _zz_toplevel_execute_ctrl1_down_execute_lane1_logic_completions_onCtrl_1_ENABLE_lane1_3;
  wire       [0:0]    _zz_toplevel_execute_ctrl1_down_execute_lane1_logic_completions_onCtrl_2_ENABLE_lane1_1;
  wire       [0:0]    _zz_toplevel_execute_ctrl1_down_execute_lane1_logic_completions_onCtrl_2_ENABLE_lane1_2;
  wire       [0:0]    _zz_toplevel_execute_ctrl1_down_early1_IntAluPlugin_ALU_ADD_SUB_lane1;
  wire       [0:0]    _zz_toplevel_execute_ctrl1_down_early1_IntAluPlugin_ALU_ADD_SUB_lane1_1;
  wire       [0:0]    _zz_toplevel_execute_ctrl1_down_early1_IntAluPlugin_ALU_SLTX_lane1;
  wire       [0:0]    _zz_toplevel_execute_ctrl1_down_early1_IntAluPlugin_ALU_SLTX_lane1_1;
  wire       [0:0]    _zz_toplevel_execute_ctrl1_down_SrcStageables_REVERT_lane1_1;
  wire       [0:0]    _zz_toplevel_execute_ctrl1_down_SrcStageables_REVERT_lane1_2;
  wire       [0:0]    _zz_toplevel_execute_ctrl1_down_SrcStageables_ZERO_lane1;
  wire       [0:0]    _zz_toplevel_execute_ctrl1_down_SrcStageables_ZERO_lane1_1;
  wire       [0:0]    _zz_toplevel_execute_ctrl1_down_lane1_IntFormatPlugin_logic_SIGNED_lane1;
  wire       [0:0]    _zz_toplevel_execute_ctrl1_down_lane1_IntFormatPlugin_logic_SIGNED_lane1_1;
  wire       [0:0]    _zz_toplevel_execute_ctrl1_down_BYPASSED_AT_2_lane1;
  wire       [0:0]    _zz_toplevel_execute_ctrl1_down_BYPASSED_AT_2_lane1_1;
  wire       [0:0]    _zz_toplevel_execute_ctrl1_down_BYPASSED_AT_3_lane1;
  wire       [0:0]    _zz_toplevel_execute_ctrl1_down_BYPASSED_AT_3_lane1_1;
  wire       [0:0]    _zz_toplevel_execute_ctrl1_down_MAY_FLUSH_PRECISE_3_lane1;
  wire       [0:0]    _zz_toplevel_execute_ctrl1_down_MAY_FLUSH_PRECISE_3_lane1_1;
  wire       [0:0]    _zz_toplevel_execute_ctrl1_down_MAY_FLUSH_PRECISE_4_lane1;
  wire       [0:0]    _zz_toplevel_execute_ctrl1_down_MAY_FLUSH_PRECISE_4_lane1_1;
  wire       [0:0]    _zz_toplevel_execute_ctrl1_down_SrcStageables_UNSIGNED_lane1;
  wire       [0:0]    _zz_toplevel_execute_ctrl1_down_SrcStageables_UNSIGNED_lane1_1;
  wire       [0:0]    _zz_toplevel_execute_ctrl1_down_BarrelShifterPlugin_LEFT_lane1_1;
  wire       [0:0]    _zz_toplevel_execute_ctrl1_down_BarrelShifterPlugin_LEFT_lane1_2;
  wire       [0:0]    _zz_toplevel_execute_ctrl1_down_BarrelShifterPlugin_SIGNED_lane1;
  wire       [0:0]    _zz_toplevel_execute_ctrl1_down_BarrelShifterPlugin_SIGNED_lane1_1;
  wire       [0:0]    _zz_toplevel_execute_ctrl1_down_late1_IntAluPlugin_ALU_ADD_SUB_lane1_1;
  wire       [0:0]    _zz_toplevel_execute_ctrl1_down_late1_IntAluPlugin_ALU_ADD_SUB_lane1_2;
  wire       [0:0]    _zz_toplevel_execute_ctrl1_down_late1_IntAluPlugin_ALU_SLTX_lane1_1;
  wire       [0:0]    _zz_toplevel_execute_ctrl1_down_late1_IntAluPlugin_ALU_SLTX_lane1_2;
  wire                _zz_when_ExecuteLanePlugin_l300_7;
  wire                _zz_when_ExecuteLanePlugin_l300_7_1;
  wire                _zz_when_ExecuteLanePlugin_l300_7_2;
  wire                _zz_when_ExecuteLanePlugin_l300_7_3;
  wire                _zz_when_ExecuteLanePlugin_l300_7_4;
  wire                _zz_when_ExecuteLanePlugin_l300_7_5;
  wire                _zz_when_ExecuteLanePlugin_l300_8;
  wire                _zz_when_ExecuteLanePlugin_l300_8_1;
  wire                _zz_when_ExecuteLanePlugin_l300_8_2;
  wire                _zz_when_ExecuteLanePlugin_l300_9;
  wire                _zz_when_ExecuteLanePlugin_l300_9_1;
  wire       [0:0]    _zz_FetchL1Plugin_pmaBuilder_onTransfers_0_addressHit;
  wire       [0:0]    _zz_FetchL1Plugin_logic_ctrl_pmaPort_rsp_io_1;
  wire       [0:0]    _zz_LsuPlugin_pmaBuilder_l1_onTransfers_0_addressHit;
  wire       [0:0]    _zz_LsuPlugin_logic_onPma_cached_rsp_io_1;
  wire       [0:0]    _zz_LsuPlugin_pmaBuilder_io_onTransfers_0_addressHit;
  wire       [0:0]    _zz_LsuPlugin_pmaBuilder_io_onTransfers_1_addressHit;
  wire       [0:0]    _zz_LsuPlugin_logic_onPma_io_rsp_io_2;
  reg        [1:0]    _zz_WhiteboxerPlugin_logic_perf_candidatesCount;
  wire       [2:0]    _zz_WhiteboxerPlugin_logic_perf_candidatesCount_1;
  reg        [1:0]    _zz_WhiteboxerPlugin_logic_perf_dispatchFeedCount;
  wire       [1:0]    _zz_WhiteboxerPlugin_logic_perf_dispatchFeedCount_1;
  wire       [59:0]   _zz__zz_WhiteboxerPlugin_logic_perf_executeFreezedCounter_1;
  wire       [0:0]    _zz__zz_WhiteboxerPlugin_logic_perf_executeFreezedCounter_1_1;
  wire       [59:0]   _zz__zz_WhiteboxerPlugin_logic_perf_dispatchHazardsCounter_1;
  wire       [0:0]    _zz__zz_WhiteboxerPlugin_logic_perf_dispatchHazardsCounter_1_1;
  wire       [59:0]   _zz__zz_WhiteboxerPlugin_logic_perf_candidatesCountCounters_0_1;
  wire       [0:0]    _zz__zz_WhiteboxerPlugin_logic_perf_candidatesCountCounters_0_1_1;
  wire       [59:0]   _zz__zz_WhiteboxerPlugin_logic_perf_candidatesCountCounters_1_1;
  wire       [0:0]    _zz__zz_WhiteboxerPlugin_logic_perf_candidatesCountCounters_1_1_1;
  wire       [59:0]   _zz__zz_WhiteboxerPlugin_logic_perf_candidatesCountCounters_2_1;
  wire       [0:0]    _zz__zz_WhiteboxerPlugin_logic_perf_candidatesCountCounters_2_1_1;
  wire       [59:0]   _zz__zz_WhiteboxerPlugin_logic_perf_candidatesCountCounters_3_1;
  wire       [0:0]    _zz__zz_WhiteboxerPlugin_logic_perf_candidatesCountCounters_3_1_1;
  wire       [59:0]   _zz__zz_WhiteboxerPlugin_logic_perf_dispatchFeedCounters_0_1;
  wire       [0:0]    _zz__zz_WhiteboxerPlugin_logic_perf_dispatchFeedCounters_0_1_1;
  wire       [59:0]   _zz__zz_WhiteboxerPlugin_logic_perf_dispatchFeedCounters_1_1;
  wire       [0:0]    _zz__zz_WhiteboxerPlugin_logic_perf_dispatchFeedCounters_1_1_1;
  wire       [59:0]   _zz__zz_WhiteboxerPlugin_logic_perf_dispatchFeedCounters_2_1;
  wire       [0:0]    _zz__zz_WhiteboxerPlugin_logic_perf_dispatchFeedCounters_2_1_1;
  wire       [1:0]    _zz_FetchL1Plugin_logic_translationStorage_logic_sl_0_write_mask;
  wire       [1:0]    _zz_LsuPlugin_logic_translationStorage_logic_sl_0_write_mask;
  wire                toplevel_decode_ctrls_0_up_isValid;
  wire                fetch_logic_ctrls_0_up_isReady;
  wire                fetch_logic_ctrls_0_up_isValid;
  reg        [31:0]   toplevel_execute_ctrl5_up_lane1_integer_WriteBackPlugin_logic_DATA_lane1;
  reg        [31:0]   toplevel_execute_ctrl5_up_lane0_integer_WriteBackPlugin_logic_DATA_lane0;
  reg                 toplevel_execute_ctrl5_up_COMMIT_lane1;
  reg                 toplevel_execute_ctrl5_up_COMMIT_lane0;
  reg        [0:0]    toplevel_execute_ctrl5_up_LANE_AGE_lane1;
  reg        [4:0]    toplevel_execute_ctrl5_up_RD_PHYS_lane1;
  reg        [0:0]    toplevel_execute_ctrl5_up_LANE_AGE_lane0;
  reg        [4:0]    toplevel_execute_ctrl5_up_RD_PHYS_lane0;
  wire       [11:0]   toplevel_execute_ctrl3_down_Decode_STORE_ID_lane0;
  wire                toplevel_execute_ctrl3_down_LsuL1_PREFETCH_lane0;
  wire       [3:0]    toplevel_execute_ctrl3_down_LsuL1_MASK_lane0;
  wire                toplevel_execute_ctrl3_down_LsuPlugin_logic_FROM_ACCESS_lane0;
  wire       [31:0]   toplevel_execute_ctrl3_down_early1_BranchPlugin_pcCalc_PC_LAST_SLICE_lane1;
  wire       [31:0]   toplevel_execute_ctrl3_down_early0_BranchPlugin_pcCalc_PC_LAST_SLICE_lane0;
  wire       [1:0]    toplevel_execute_ctrl3_down_late1_IntAluPlugin_ALU_BITWISE_CTRL_lane1;
  wire                toplevel_execute_ctrl3_down_late1_IntAluPlugin_ALU_SLTX_lane1;
  wire                toplevel_execute_ctrl3_down_late1_IntAluPlugin_ALU_ADD_SUB_lane1;
  wire                toplevel_execute_ctrl3_down_BarrelShifterPlugin_SIGNED_lane1;
  wire                toplevel_execute_ctrl3_down_BarrelShifterPlugin_LEFT_lane1;
  wire                toplevel_execute_ctrl3_down_SrcStageables_UNSIGNED_lane1;
  wire                toplevel_execute_ctrl3_down_SrcStageables_ZERO_lane1;
  wire                toplevel_execute_ctrl3_down_SrcStageables_REVERT_lane1;
  wire                toplevel_execute_ctrl3_down_execute_lane1_logic_completions_onCtrl_2_ENABLE_lane1;
  wire                toplevel_execute_ctrl3_down_COMPLETION_AT_4_lane1;
  wire                toplevel_execute_ctrl3_down_lane1_integer_WriteBackPlugin_SEL_lane1;
  wire                toplevel_execute_ctrl3_down_late1_BranchPlugin_SEL_lane1;
  wire                toplevel_execute_ctrl3_down_late1_BarrelShifterPlugin_SEL_lane1;
  wire                toplevel_execute_ctrl3_down_late1_IntAluPlugin_SEL_lane1;
  wire       [1:0]    toplevel_execute_ctrl3_down_late0_IntAluPlugin_ALU_BITWISE_CTRL_lane0;
  wire                toplevel_execute_ctrl3_down_late0_IntAluPlugin_ALU_SLTX_lane0;
  wire                toplevel_execute_ctrl3_down_late0_IntAluPlugin_ALU_ADD_SUB_lane0;
  wire                toplevel_execute_ctrl3_down_LsuPlugin_logic_LSU_PREFETCH_lane0;
  wire                toplevel_execute_ctrl3_down_AguPlugin_FLOAT_lane0;
  wire                toplevel_execute_ctrl3_down_AguPlugin_ATOMIC_lane0;
  wire                toplevel_execute_ctrl3_down_AguPlugin_LOAD_lane0;
  wire                toplevel_execute_ctrl3_down_BarrelShifterPlugin_SIGNED_lane0;
  wire                toplevel_execute_ctrl3_down_BarrelShifterPlugin_LEFT_lane0;
  wire                toplevel_execute_ctrl3_down_SrcStageables_UNSIGNED_lane0;
  wire       [1:0]    toplevel_execute_ctrl3_down_lane0_IntFormatPlugin_logic_WIDTH_ID_lane0;
  wire                toplevel_execute_ctrl3_down_lane0_IntFormatPlugin_logic_SIGNED_lane0;
  wire                toplevel_execute_ctrl3_down_SrcStageables_ZERO_lane0;
  wire                toplevel_execute_ctrl3_down_SrcStageables_REVERT_lane0;
  wire                toplevel_execute_ctrl3_down_execute_lane0_logic_completions_onCtrl_2_ENABLE_lane0;
  wire                toplevel_execute_ctrl3_down_COMPLETION_AT_4_lane0;
  wire                toplevel_execute_ctrl3_down_lane0_integer_WriteBackPlugin_SEL_lane0;
  wire                toplevel_execute_ctrl3_down_MulPlugin_HIGH_lane0;
  wire                toplevel_execute_ctrl3_down_late0_BranchPlugin_SEL_lane0;
  wire                toplevel_execute_ctrl3_down_late0_BarrelShifterPlugin_SEL_lane0;
  wire                toplevel_execute_ctrl3_down_late0_IntAluPlugin_SEL_lane0;
  wire                toplevel_execute_ctrl3_down_early0_MulPlugin_SEL_lane0;
  wire       [1:0]    toplevel_execute_ctrl3_down_AguPlugin_SIZE_lane0;
  wire       [0:0]    toplevel_execute_ctrl3_down_Decode_INSTRUCTION_SLICE_COUNT_lane1;
  wire       [1:0]    toplevel_execute_ctrl3_down_GSharePlugin_GSHARE_COUNTER_lane1_0;
  wire       [1:0]    toplevel_execute_ctrl3_down_GSharePlugin_GSHARE_COUNTER_lane1_1;
  wire       [1:0]    toplevel_execute_ctrl3_down_GSharePlugin_GSHARE_COUNTER_lane1_2;
  wire       [1:0]    toplevel_execute_ctrl3_down_GSharePlugin_GSHARE_COUNTER_lane1_3;
  wire       [31:0]   toplevel_execute_ctrl3_down_Prediction_ALIGNED_JUMPED_PC_lane1;
  wire       [0:0]    toplevel_execute_ctrl3_down_Decode_INSTRUCTION_SLICE_COUNT_lane0;
  wire       [1:0]    toplevel_execute_ctrl3_down_GSharePlugin_GSHARE_COUNTER_lane0_0;
  wire       [1:0]    toplevel_execute_ctrl3_down_GSharePlugin_GSHARE_COUNTER_lane0_1;
  wire       [1:0]    toplevel_execute_ctrl3_down_GSharePlugin_GSHARE_COUNTER_lane0_2;
  wire       [1:0]    toplevel_execute_ctrl3_down_GSharePlugin_GSHARE_COUNTER_lane0_3;
  wire       [31:0]   toplevel_execute_ctrl3_down_Prediction_ALIGNED_JUMPED_PC_lane0;
  reg                 toplevel_execute_ctrl4_up_MMU_BYPASS_TRANSLATION_lane0;
  reg                 toplevel_execute_ctrl4_up_MMU_HAZARD_lane0;
  reg                 toplevel_execute_ctrl4_up_MMU_REFILL_lane0;
  reg                 toplevel_execute_ctrl4_up_MMU_ACCESS_FAULT_lane0;
  reg                 toplevel_execute_ctrl4_up_LsuPlugin_logic_MMU_FAILURE_lane0;
  reg                 toplevel_execute_ctrl4_up_LsuPlugin_logic_MMU_PAGE_FAULT_lane0;
  reg                 toplevel_execute_ctrl4_up_LsuPlugin_logic_onPma_FROM_LSU_MSB_FAILED_lane0;
  reg                 toplevel_execute_ctrl4_up_LsuPlugin_logic_onPma_IO_lane0;
  reg                 toplevel_execute_ctrl4_up_LsuPlugin_logic_onPma_IO_RSP_lane0_fault;
  reg                 toplevel_execute_ctrl4_up_LsuPlugin_logic_onPma_IO_RSP_lane0_io;
  reg                 toplevel_execute_ctrl4_up_LsuPlugin_logic_onPma_CACHED_RSP_lane0_fault;
  reg                 toplevel_execute_ctrl4_up_LsuPlugin_logic_onPma_CACHED_RSP_lane0_io;
  reg                 toplevel_execute_ctrl4_up_LsuPlugin_logic_preCtrl_IS_AMO_lane0;
  reg                 toplevel_execute_ctrl4_up_LsuPlugin_logic_preCtrl_MISS_ALIGNED_lane0;
  reg        [31:0]   toplevel_execute_ctrl4_up_MMU_TRANSLATED_lane0;
  reg                 toplevel_execute_ctrl4_up_LsuPlugin_logic_onTrigger_HIT_lane0;
  reg        [1:0]    toplevel_execute_ctrl4_up_LsuL1Plugin_logic_WAYS_HITS_lane0;
  reg                 toplevel_execute_ctrl4_up_LsuL1Plugin_logic_WAYS_TAGS_lane0_0_loaded;
  reg        [19:0]   toplevel_execute_ctrl4_up_LsuL1Plugin_logic_WAYS_TAGS_lane0_0_address;
  reg                 toplevel_execute_ctrl4_up_LsuL1Plugin_logic_WAYS_TAGS_lane0_0_fault;
  reg                 toplevel_execute_ctrl4_up_LsuL1Plugin_logic_WAYS_TAGS_lane0_1_loaded;
  reg        [19:0]   toplevel_execute_ctrl4_up_LsuL1Plugin_logic_WAYS_TAGS_lane0_1_address;
  reg                 toplevel_execute_ctrl4_up_LsuL1Plugin_logic_WAYS_TAGS_lane0_1_fault;
  reg        [31:0]   toplevel_execute_ctrl4_up_LsuL1_PHYSICAL_ADDRESS_lane0;
  reg        [1:0]    toplevel_execute_ctrl4_up_LsuL1Plugin_logic_WRITE_TO_READ_HAZARDS_lane0;
  reg        [31:0]   toplevel_execute_ctrl4_up_LsuL1Plugin_logic_BANKS_MUXES_lane0_0;
  reg        [31:0]   toplevel_execute_ctrl4_up_LsuL1Plugin_logic_BANKS_MUXES_lane0_1;
  reg        [1:0]    toplevel_execute_ctrl4_up_LsuL1Plugin_logic_BANK_BUSY_REMAPPED_lane0;
  reg        [31:0]   toplevel_execute_ctrl4_up_late1_SrcPlugin_SRC2_lane1;
  reg        [31:0]   toplevel_execute_ctrl4_up_late1_SrcPlugin_SRC1_lane1;
  reg        [31:0]   toplevel_execute_ctrl4_up_late0_SrcPlugin_SRC2_lane0;
  reg        [31:0]   toplevel_execute_ctrl4_up_late0_SrcPlugin_SRC1_lane0;
  reg        [4:0]    toplevel_execute_ctrl4_up_early0_MulPlugin_logic_steps_0_adders_1_lane0;
  reg        [62:0]   toplevel_execute_ctrl4_up_early0_MulPlugin_logic_steps_0_adders_0_lane0;
  reg        [0:0]    toplevel_execute_ctrl4_up_LsuL1Plugin_logic_SHARED_lane0_plru_0;
  reg        [1:0]    toplevel_execute_ctrl4_up_LsuL1Plugin_logic_SHARED_lane0_dirty;
  reg                 toplevel_execute_ctrl4_up_LsuPlugin_logic_FROM_PREFETCH_lane0;
  reg                 toplevel_execute_ctrl4_up_LsuPlugin_logic_FROM_LSU_lane0;
  reg        [11:0]   toplevel_execute_ctrl4_up_Decode_STORE_ID_lane0;
  reg                 toplevel_execute_ctrl4_up_LsuL1_FLUSH_lane0;
  reg                 toplevel_execute_ctrl4_up_LsuL1_PREFETCH_lane0;
  reg                 toplevel_execute_ctrl4_up_LsuL1_STORE_lane0;
  reg                 toplevel_execute_ctrl4_up_LsuL1_ATOMIC_lane0;
  reg                 toplevel_execute_ctrl4_up_LsuL1_LOAD_lane0;
  reg        [1:0]    toplevel_execute_ctrl4_up_LsuL1_SIZE_lane0;
  reg        [3:0]    toplevel_execute_ctrl4_up_LsuL1_MASK_lane0;
  reg                 toplevel_execute_ctrl4_up_LsuPlugin_logic_FROM_ACCESS_lane0;
  reg        [3:0]    toplevel_execute_ctrl4_up_LsuL1Plugin_logic_EVENT_WRITE_MASK_lane0;
  reg        [31:0]   toplevel_execute_ctrl4_up_LsuL1Plugin_logic_EVENT_WRITE_DATA_lane0;
  reg        [31:0]   toplevel_execute_ctrl4_up_LsuL1_MIXED_ADDRESS_lane0;
  reg        [31:0]   toplevel_execute_ctrl4_up_early1_BranchPlugin_pcCalc_PC_LAST_SLICE_lane1;
  reg        [31:0]   toplevel_execute_ctrl4_up_early1_BranchPlugin_pcCalc_PC_FALSE_lane1;
  reg        [31:0]   toplevel_execute_ctrl4_up_early1_BranchPlugin_pcCalc_PC_TRUE_lane1;
  reg        [31:0]   toplevel_execute_ctrl4_up_early0_BranchPlugin_pcCalc_PC_LAST_SLICE_lane0;
  reg        [31:0]   toplevel_execute_ctrl4_up_early0_BranchPlugin_pcCalc_PC_FALSE_lane0;
  reg        [31:0]   toplevel_execute_ctrl4_up_early0_BranchPlugin_pcCalc_PC_TRUE_lane0;
  reg                 toplevel_execute_ctrl4_up_COMMIT_lane1;
  reg        [1:0]    toplevel_execute_ctrl4_up_late1_IntAluPlugin_ALU_BITWISE_CTRL_lane1;
  reg                 toplevel_execute_ctrl4_up_late1_IntAluPlugin_ALU_SLTX_lane1;
  reg                 toplevel_execute_ctrl4_up_late1_IntAluPlugin_ALU_ADD_SUB_lane1;
  reg        [1:0]    toplevel_execute_ctrl4_up_BranchPlugin_BRANCH_CTRL_lane1;
  reg                 toplevel_execute_ctrl4_up_BarrelShifterPlugin_SIGNED_lane1;
  reg                 toplevel_execute_ctrl4_up_BarrelShifterPlugin_LEFT_lane1;
  reg                 toplevel_execute_ctrl4_up_SrcStageables_UNSIGNED_lane1;
  reg                 toplevel_execute_ctrl4_up_SrcStageables_ZERO_lane1;
  reg                 toplevel_execute_ctrl4_up_SrcStageables_REVERT_lane1;
  reg                 toplevel_execute_ctrl4_up_execute_lane1_logic_completions_onCtrl_2_ENABLE_lane1;
  reg                 toplevel_execute_ctrl4_up_COMPLETION_AT_4_lane1;
  reg                 toplevel_execute_ctrl4_up_lane1_integer_WriteBackPlugin_SEL_lane1;
  reg                 toplevel_execute_ctrl4_up_late1_BranchPlugin_SEL_lane1;
  reg                 toplevel_execute_ctrl4_up_late1_BarrelShifterPlugin_SEL_lane1;
  reg                 toplevel_execute_ctrl4_up_late1_IntAluPlugin_SEL_lane1;
  reg                 toplevel_execute_ctrl4_up_early1_BranchPlugin_SEL_lane1;
  reg        [1:0]    toplevel_execute_ctrl4_up_late0_IntAluPlugin_ALU_BITWISE_CTRL_lane0;
  reg                 toplevel_execute_ctrl4_up_late0_IntAluPlugin_ALU_SLTX_lane0;
  reg                 toplevel_execute_ctrl4_up_late0_IntAluPlugin_ALU_ADD_SUB_lane0;
  reg                 toplevel_execute_ctrl4_up_LsuPlugin_logic_LSU_PREFETCH_lane0;
  reg                 toplevel_execute_ctrl4_up_AguPlugin_FLOAT_lane0;
  reg                 toplevel_execute_ctrl4_up_AguPlugin_ATOMIC_lane0;
  reg                 toplevel_execute_ctrl4_up_AguPlugin_STORE_lane0;
  reg                 toplevel_execute_ctrl4_up_AguPlugin_LOAD_lane0;
  reg        [1:0]    toplevel_execute_ctrl4_up_BranchPlugin_BRANCH_CTRL_lane0;
  reg                 toplevel_execute_ctrl4_up_BarrelShifterPlugin_SIGNED_lane0;
  reg                 toplevel_execute_ctrl4_up_BarrelShifterPlugin_LEFT_lane0;
  reg                 toplevel_execute_ctrl4_up_SrcStageables_UNSIGNED_lane0;
  reg        [1:0]    toplevel_execute_ctrl4_up_lane0_IntFormatPlugin_logic_WIDTH_ID_lane0;
  reg                 toplevel_execute_ctrl4_up_lane0_IntFormatPlugin_logic_SIGNED_lane0;
  reg                 toplevel_execute_ctrl4_up_SrcStageables_ZERO_lane0;
  reg                 toplevel_execute_ctrl4_up_SrcStageables_REVERT_lane0;
  reg                 toplevel_execute_ctrl4_up_execute_lane0_logic_completions_onCtrl_2_ENABLE_lane0;
  reg                 toplevel_execute_ctrl4_up_COMPLETION_AT_4_lane0;
  reg                 toplevel_execute_ctrl4_up_lane0_integer_WriteBackPlugin_SEL_lane0;
  reg                 toplevel_execute_ctrl4_up_LsuPlugin_logic_FENCE_lane0;
  reg                 toplevel_execute_ctrl4_up_AguPlugin_SEL_lane0;
  reg                 toplevel_execute_ctrl4_up_MulPlugin_HIGH_lane0;
  reg                 toplevel_execute_ctrl4_up_late0_BranchPlugin_SEL_lane0;
  reg                 toplevel_execute_ctrl4_up_late0_BarrelShifterPlugin_SEL_lane0;
  reg                 toplevel_execute_ctrl4_up_late0_IntAluPlugin_SEL_lane0;
  reg                 toplevel_execute_ctrl4_up_early0_MulPlugin_SEL_lane0;
  reg                 toplevel_execute_ctrl4_up_early0_BranchPlugin_SEL_lane0;
  reg        [1:0]    toplevel_execute_ctrl4_up_AguPlugin_SIZE_lane0;
  reg        [0:0]    toplevel_execute_ctrl4_up_LANE_AGE_lane1;
  reg        [4:0]    toplevel_execute_ctrl4_up_RD_PHYS_lane1;
  reg        [15:0]   toplevel_execute_ctrl4_up_Decode_UOP_ID_lane1;
  reg                 toplevel_execute_ctrl4_up_TRAP_lane1;
  reg        [31:0]   toplevel_execute_ctrl4_up_PC_lane1;
  reg        [0:0]    toplevel_execute_ctrl4_up_Decode_INSTRUCTION_SLICE_COUNT_lane1;
  reg        [11:0]   toplevel_execute_ctrl4_up_Prediction_BRANCH_HISTORY_lane1;
  reg        [1:0]    toplevel_execute_ctrl4_up_GSharePlugin_GSHARE_COUNTER_lane1_0;
  reg        [1:0]    toplevel_execute_ctrl4_up_GSharePlugin_GSHARE_COUNTER_lane1_1;
  reg        [1:0]    toplevel_execute_ctrl4_up_GSharePlugin_GSHARE_COUNTER_lane1_2;
  reg        [1:0]    toplevel_execute_ctrl4_up_GSharePlugin_GSHARE_COUNTER_lane1_3;
  reg        [3:0]    toplevel_execute_ctrl4_up_Prediction_ALIGNED_SLICES_BRANCH_lane1;
  reg        [3:0]    toplevel_execute_ctrl4_up_Prediction_ALIGNED_SLICES_TAKEN_lane1;
  reg        [31:0]   toplevel_execute_ctrl4_up_Prediction_ALIGNED_JUMPED_PC_lane1;
  reg                 toplevel_execute_ctrl4_up_Prediction_ALIGNED_JUMPED_lane1;
  reg        [31:0]   toplevel_execute_ctrl4_up_Decode_UOP_lane1;
  reg        [0:0]    toplevel_execute_ctrl4_up_LANE_AGE_lane0;
  reg        [4:0]    toplevel_execute_ctrl4_up_RD_PHYS_lane0;
  reg        [15:0]   toplevel_execute_ctrl4_up_Decode_UOP_ID_lane0;
  reg        [31:0]   toplevel_execute_ctrl4_up_PC_lane0;
  reg        [0:0]    toplevel_execute_ctrl4_up_Decode_INSTRUCTION_SLICE_COUNT_lane0;
  reg        [11:0]   toplevel_execute_ctrl4_up_Prediction_BRANCH_HISTORY_lane0;
  reg        [1:0]    toplevel_execute_ctrl4_up_GSharePlugin_GSHARE_COUNTER_lane0_0;
  reg        [1:0]    toplevel_execute_ctrl4_up_GSharePlugin_GSHARE_COUNTER_lane0_1;
  reg        [1:0]    toplevel_execute_ctrl4_up_GSharePlugin_GSHARE_COUNTER_lane0_2;
  reg        [1:0]    toplevel_execute_ctrl4_up_GSharePlugin_GSHARE_COUNTER_lane0_3;
  reg        [3:0]    toplevel_execute_ctrl4_up_Prediction_ALIGNED_SLICES_BRANCH_lane0;
  reg        [3:0]    toplevel_execute_ctrl4_up_Prediction_ALIGNED_SLICES_TAKEN_lane0;
  reg        [31:0]   toplevel_execute_ctrl4_up_Prediction_ALIGNED_JUMPED_PC_lane0;
  reg                 toplevel_execute_ctrl4_up_Prediction_ALIGNED_JUMPED_lane0;
  reg        [31:0]   toplevel_execute_ctrl4_up_Decode_UOP_lane0;
  wire       [1:0]    toplevel_execute_ctrl2_down_late1_SrcPlugin_logic_SRC2_CTRL_lane1;
  wire       [0:0]    toplevel_execute_ctrl2_down_late1_SrcPlugin_logic_SRC1_CTRL_lane1;
  wire       [1:0]    toplevel_execute_ctrl2_down_late1_IntAluPlugin_ALU_BITWISE_CTRL_lane1;
  wire                toplevel_execute_ctrl2_down_late1_IntAluPlugin_ALU_SLTX_lane1;
  wire                toplevel_execute_ctrl2_down_late1_IntAluPlugin_ALU_ADD_SUB_lane1;
  wire                toplevel_execute_ctrl2_down_execute_lane1_logic_completions_onCtrl_2_ENABLE_lane1;
  wire                toplevel_execute_ctrl2_down_execute_lane1_logic_completions_onCtrl_1_ENABLE_lane1;
  wire                toplevel_execute_ctrl2_down_COMPLETION_AT_4_lane1;
  wire                toplevel_execute_ctrl2_down_COMPLETION_AT_3_lane1;
  wire                toplevel_execute_ctrl2_down_lane1_integer_WriteBackPlugin_SEL_lane1;
  wire                toplevel_execute_ctrl2_down_late1_BranchPlugin_SEL_lane1;
  wire                toplevel_execute_ctrl2_down_late1_BarrelShifterPlugin_SEL_lane1;
  wire                toplevel_execute_ctrl2_down_late1_IntAluPlugin_SEL_lane1;
  wire                toplevel_execute_ctrl2_down_early1_BarrelShifterPlugin_SEL_lane1;
  wire       [1:0]    toplevel_execute_ctrl2_down_late0_SrcPlugin_logic_SRC2_CTRL_lane0;
  wire       [0:0]    toplevel_execute_ctrl2_down_late0_SrcPlugin_logic_SRC1_CTRL_lane0;
  wire       [1:0]    toplevel_execute_ctrl2_down_late0_IntAluPlugin_ALU_BITWISE_CTRL_lane0;
  wire                toplevel_execute_ctrl2_down_late0_IntAluPlugin_ALU_SLTX_lane0;
  wire                toplevel_execute_ctrl2_down_late0_IntAluPlugin_ALU_ADD_SUB_lane0;
  wire                toplevel_execute_ctrl2_down_LsuPlugin_logic_LSU_PREFETCH_lane0;
  wire                toplevel_execute_ctrl2_down_AguPlugin_FLOAT_lane0;
  wire       [1:0]    toplevel_execute_ctrl2_down_lane0_IntFormatPlugin_logic_WIDTH_ID_lane0;
  wire                toplevel_execute_ctrl2_down_lane0_IntFormatPlugin_logic_SIGNED_lane0;
  wire                toplevel_execute_ctrl2_down_execute_lane0_logic_completions_onCtrl_2_ENABLE_lane0;
  wire                toplevel_execute_ctrl2_down_execute_lane0_logic_completions_onCtrl_1_ENABLE_lane0;
  wire                toplevel_execute_ctrl2_down_COMPLETION_AT_4_lane0;
  wire                toplevel_execute_ctrl2_down_COMPLETION_AT_3_lane0;
  wire                toplevel_execute_ctrl2_down_lane0_integer_WriteBackPlugin_SEL_lane0;
  wire                toplevel_execute_ctrl2_down_LsuPlugin_logic_FENCE_lane0;
  wire                toplevel_execute_ctrl2_down_MulPlugin_HIGH_lane0;
  wire                toplevel_execute_ctrl2_down_late0_BranchPlugin_SEL_lane0;
  wire                toplevel_execute_ctrl2_down_late0_BarrelShifterPlugin_SEL_lane0;
  wire                toplevel_execute_ctrl2_down_late0_IntAluPlugin_SEL_lane0;
  wire                toplevel_execute_ctrl2_down_early0_MulPlugin_SEL_lane0;
  wire                toplevel_execute_ctrl2_down_early0_BarrelShifterPlugin_SEL_lane0;
  wire       [11:0]   toplevel_execute_ctrl2_down_Prediction_BRANCH_HISTORY_lane1;
  wire       [1:0]    toplevel_execute_ctrl2_down_GSharePlugin_GSHARE_COUNTER_lane1_0;
  wire       [1:0]    toplevel_execute_ctrl2_down_GSharePlugin_GSHARE_COUNTER_lane1_1;
  wire       [1:0]    toplevel_execute_ctrl2_down_GSharePlugin_GSHARE_COUNTER_lane1_2;
  wire       [1:0]    toplevel_execute_ctrl2_down_GSharePlugin_GSHARE_COUNTER_lane1_3;
  wire       [3:0]    toplevel_execute_ctrl2_down_Prediction_ALIGNED_SLICES_BRANCH_lane1;
  wire       [3:0]    toplevel_execute_ctrl2_down_Prediction_ALIGNED_SLICES_TAKEN_lane1;
  wire                toplevel_execute_ctrl2_down_Prediction_ALIGNED_JUMPED_lane1;
  wire       [11:0]   toplevel_execute_ctrl2_down_Prediction_BRANCH_HISTORY_lane0;
  wire       [1:0]    toplevel_execute_ctrl2_down_GSharePlugin_GSHARE_COUNTER_lane0_0;
  wire       [1:0]    toplevel_execute_ctrl2_down_GSharePlugin_GSHARE_COUNTER_lane0_1;
  wire       [1:0]    toplevel_execute_ctrl2_down_GSharePlugin_GSHARE_COUNTER_lane0_2;
  wire       [1:0]    toplevel_execute_ctrl2_down_GSharePlugin_GSHARE_COUNTER_lane0_3;
  wire       [3:0]    toplevel_execute_ctrl2_down_Prediction_ALIGNED_SLICES_BRANCH_lane0;
  wire       [3:0]    toplevel_execute_ctrl2_down_Prediction_ALIGNED_SLICES_TAKEN_lane0;
  wire                toplevel_execute_ctrl2_down_Prediction_ALIGNED_JUMPED_lane0;
  reg                 toplevel_execute_ctrl3_up_LsuPlugin_logic_FROM_PREFETCH_lane0;
  reg                 toplevel_execute_ctrl3_up_LsuPlugin_logic_FROM_LSU_lane0;
  reg        [11:0]   toplevel_execute_ctrl3_up_Decode_STORE_ID_lane0;
  reg                 toplevel_execute_ctrl3_up_LsuL1_FLUSH_lane0;
  reg                 toplevel_execute_ctrl3_up_LsuL1_PREFETCH_lane0;
  reg                 toplevel_execute_ctrl3_up_LsuL1_STORE_lane0;
  reg                 toplevel_execute_ctrl3_up_LsuL1_ATOMIC_lane0;
  reg                 toplevel_execute_ctrl3_up_LsuL1_LOAD_lane0;
  reg        [1:0]    toplevel_execute_ctrl3_up_LsuL1_SIZE_lane0;
  reg        [3:0]    toplevel_execute_ctrl3_up_LsuL1_MASK_lane0;
  reg                 toplevel_execute_ctrl3_up_LsuPlugin_logic_FROM_ACCESS_lane0;
  reg                 toplevel_execute_ctrl3_up_LsuPlugin_logic_FORCE_PHYSICAL_lane0;
  reg        [3:0]    toplevel_execute_ctrl3_up_LsuL1Plugin_logic_EVENT_WRITE_MASK_lane0;
  reg        [31:0]   toplevel_execute_ctrl3_up_LsuL1Plugin_logic_EVENT_WRITE_DATA_lane0;
  reg        [0:0]    toplevel_execute_ctrl3_up_LsuL1Plugin_logic_ls_rt0_SHARED_BYPASS_VALUE_lane0_plru_0;
  reg        [1:0]    toplevel_execute_ctrl3_up_LsuL1Plugin_logic_ls_rt0_SHARED_BYPASS_VALUE_lane0_dirty;
  reg                 toplevel_execute_ctrl3_up_LsuL1Plugin_logic_ls_rt0_SHARED_BYPASS_VALID_lane0;
  reg        [31:0]   toplevel_execute_ctrl3_up_LsuL1Plugin_logic_EVENT_WRITE_ADDRESS_lane0;
  reg                 toplevel_execute_ctrl3_up_LsuL1Plugin_logic_EVENT_WRITE_VALID_lane0;
  reg        [1:0]    toplevel_execute_ctrl3_up_LsuL1Plugin_logic_BANK_BUSY_lane0;
  reg        [31:0]   toplevel_execute_ctrl3_up_LsuL1_MIXED_ADDRESS_lane0;
  reg                 toplevel_execute_ctrl3_up_early1_BranchPlugin_logic_alu_MSB_FAILED_lane1;
  reg                 toplevel_execute_ctrl3_up_early1_BranchPlugin_logic_alu_btb_BAD_TARGET_lane1;
  reg                 toplevel_execute_ctrl3_up_early1_BranchPlugin_logic_alu_EQ_lane1;
  reg                 toplevel_execute_ctrl3_up_early0_BranchPlugin_logic_alu_MSB_FAILED_lane0;
  reg                 toplevel_execute_ctrl3_up_early0_BranchPlugin_logic_alu_btb_BAD_TARGET_lane0;
  reg                 toplevel_execute_ctrl3_up_early0_BranchPlugin_logic_alu_EQ_lane0;
  reg        [31:0]   toplevel_execute_ctrl3_up_early1_BranchPlugin_pcCalc_PC_LAST_SLICE_lane1;
  reg        [31:0]   toplevel_execute_ctrl3_up_early1_BranchPlugin_pcCalc_PC_FALSE_lane1;
  reg        [31:0]   toplevel_execute_ctrl3_up_early1_BranchPlugin_pcCalc_PC_TRUE_lane1;
  reg        [31:0]   toplevel_execute_ctrl3_up_early0_BranchPlugin_pcCalc_PC_LAST_SLICE_lane0;
  reg        [31:0]   toplevel_execute_ctrl3_up_early0_BranchPlugin_pcCalc_PC_FALSE_lane0;
  reg        [31:0]   toplevel_execute_ctrl3_up_early0_BranchPlugin_pcCalc_PC_TRUE_lane0;
  reg        [31:0]   toplevel_execute_ctrl3_up_early1_BarrelShifterPlugin_SHIFT_RESULT_lane1;
  reg                 toplevel_execute_ctrl3_up_early1_SrcPlugin_LESS_lane1;
  reg        [31:0]   toplevel_execute_ctrl3_up_DivPlugin_DIV_RESULT_lane0;
  reg        [32:0]   toplevel_execute_ctrl3_up_MUL_SRC2_lane0;
  reg        [32:0]   toplevel_execute_ctrl3_up_MUL_SRC1_lane0;
  reg        [31:0]   toplevel_execute_ctrl3_up_early0_BarrelShifterPlugin_SHIFT_RESULT_lane0;
  reg                 toplevel_execute_ctrl3_up_early0_SrcPlugin_LESS_lane0;
  reg        [31:0]   toplevel_execute_ctrl3_up_early0_SrcPlugin_ADD_SUB_lane0;
  reg                 toplevel_execute_ctrl3_up_COMMIT_lane1;
  reg                 toplevel_execute_ctrl3_up_COMMIT_lane0;
  reg        [1:0]    toplevel_execute_ctrl3_up_late1_SrcPlugin_logic_SRC2_CTRL_lane1;
  reg        [0:0]    toplevel_execute_ctrl3_up_late1_SrcPlugin_logic_SRC1_CTRL_lane1;
  reg        [1:0]    toplevel_execute_ctrl3_up_late1_IntAluPlugin_ALU_BITWISE_CTRL_lane1;
  reg                 toplevel_execute_ctrl3_up_late1_IntAluPlugin_ALU_SLTX_lane1;
  reg                 toplevel_execute_ctrl3_up_late1_IntAluPlugin_ALU_ADD_SUB_lane1;
  reg        [1:0]    toplevel_execute_ctrl3_up_BranchPlugin_BRANCH_CTRL_lane1;
  reg                 toplevel_execute_ctrl3_up_BarrelShifterPlugin_SIGNED_lane1;
  reg                 toplevel_execute_ctrl3_up_BarrelShifterPlugin_LEFT_lane1;
  reg                 toplevel_execute_ctrl3_up_SrcStageables_UNSIGNED_lane1;
  reg                 toplevel_execute_ctrl3_up_SrcStageables_ZERO_lane1;
  reg                 toplevel_execute_ctrl3_up_SrcStageables_REVERT_lane1;
  reg                 toplevel_execute_ctrl3_up_execute_lane1_logic_completions_onCtrl_2_ENABLE_lane1;
  reg                 toplevel_execute_ctrl3_up_execute_lane1_logic_completions_onCtrl_1_ENABLE_lane1;
  reg                 toplevel_execute_ctrl3_up_COMPLETION_AT_4_lane1;
  reg                 toplevel_execute_ctrl3_up_COMPLETION_AT_3_lane1;
  reg                 toplevel_execute_ctrl3_up_lane1_integer_WriteBackPlugin_SEL_lane1;
  reg                 toplevel_execute_ctrl3_up_late1_BranchPlugin_SEL_lane1;
  reg                 toplevel_execute_ctrl3_up_late1_BarrelShifterPlugin_SEL_lane1;
  reg                 toplevel_execute_ctrl3_up_late1_IntAluPlugin_SEL_lane1;
  reg                 toplevel_execute_ctrl3_up_early1_BranchPlugin_SEL_lane1;
  reg                 toplevel_execute_ctrl3_up_early1_BarrelShifterPlugin_SEL_lane1;
  reg        [1:0]    toplevel_execute_ctrl3_up_late0_SrcPlugin_logic_SRC2_CTRL_lane0;
  reg        [0:0]    toplevel_execute_ctrl3_up_late0_SrcPlugin_logic_SRC1_CTRL_lane0;
  reg        [1:0]    toplevel_execute_ctrl3_up_late0_IntAluPlugin_ALU_BITWISE_CTRL_lane0;
  reg                 toplevel_execute_ctrl3_up_late0_IntAluPlugin_ALU_SLTX_lane0;
  reg                 toplevel_execute_ctrl3_up_late0_IntAluPlugin_ALU_ADD_SUB_lane0;
  reg                 toplevel_execute_ctrl3_up_LsuPlugin_logic_LSU_PREFETCH_lane0;
  reg                 toplevel_execute_ctrl3_up_AguPlugin_FLOAT_lane0;
  reg                 toplevel_execute_ctrl3_up_AguPlugin_ATOMIC_lane0;
  reg                 toplevel_execute_ctrl3_up_AguPlugin_STORE_lane0;
  reg                 toplevel_execute_ctrl3_up_AguPlugin_LOAD_lane0;
  reg        [1:0]    toplevel_execute_ctrl3_up_BranchPlugin_BRANCH_CTRL_lane0;
  reg                 toplevel_execute_ctrl3_up_BarrelShifterPlugin_SIGNED_lane0;
  reg                 toplevel_execute_ctrl3_up_BarrelShifterPlugin_LEFT_lane0;
  reg                 toplevel_execute_ctrl3_up_SrcStageables_UNSIGNED_lane0;
  reg        [1:0]    toplevel_execute_ctrl3_up_lane0_IntFormatPlugin_logic_WIDTH_ID_lane0;
  reg                 toplevel_execute_ctrl3_up_lane0_IntFormatPlugin_logic_SIGNED_lane0;
  reg                 toplevel_execute_ctrl3_up_SrcStageables_ZERO_lane0;
  reg                 toplevel_execute_ctrl3_up_SrcStageables_REVERT_lane0;
  reg                 toplevel_execute_ctrl3_up_execute_lane0_logic_completions_onCtrl_2_ENABLE_lane0;
  reg                 toplevel_execute_ctrl3_up_execute_lane0_logic_completions_onCtrl_1_ENABLE_lane0;
  reg                 toplevel_execute_ctrl3_up_COMPLETION_AT_4_lane0;
  reg                 toplevel_execute_ctrl3_up_COMPLETION_AT_3_lane0;
  reg                 toplevel_execute_ctrl3_up_lane0_integer_WriteBackPlugin_SEL_lane0;
  reg                 toplevel_execute_ctrl3_up_LsuPlugin_logic_FENCE_lane0;
  reg                 toplevel_execute_ctrl3_up_AguPlugin_SEL_lane0;
  reg                 toplevel_execute_ctrl3_up_CsrAccessPlugin_SEL_lane0;
  reg                 toplevel_execute_ctrl3_up_MulPlugin_HIGH_lane0;
  reg                 toplevel_execute_ctrl3_up_late0_BranchPlugin_SEL_lane0;
  reg                 toplevel_execute_ctrl3_up_late0_BarrelShifterPlugin_SEL_lane0;
  reg                 toplevel_execute_ctrl3_up_late0_IntAluPlugin_SEL_lane0;
  reg                 toplevel_execute_ctrl3_up_early0_DivPlugin_SEL_lane0;
  reg                 toplevel_execute_ctrl3_up_early0_MulPlugin_SEL_lane0;
  reg                 toplevel_execute_ctrl3_up_early0_BranchPlugin_SEL_lane0;
  reg                 toplevel_execute_ctrl3_up_early0_BarrelShifterPlugin_SEL_lane0;
  reg        [1:0]    toplevel_execute_ctrl3_up_AguPlugin_SIZE_lane0;
  reg        [0:0]    toplevel_execute_ctrl3_up_LANE_AGE_lane1;
  reg        [4:0]    toplevel_execute_ctrl3_up_RD_PHYS_lane1;
  reg        [4:0]    toplevel_execute_ctrl3_up_RS2_PHYS_lane1;
  reg        [4:0]    toplevel_execute_ctrl3_up_RS1_PHYS_lane1;
  reg        [15:0]   toplevel_execute_ctrl3_up_Decode_UOP_ID_lane1;
  reg                 toplevel_execute_ctrl3_up_TRAP_lane1;
  reg        [31:0]   toplevel_execute_ctrl3_up_PC_lane1;
  reg        [0:0]    toplevel_execute_ctrl3_up_Decode_INSTRUCTION_SLICE_COUNT_lane1;
  reg        [11:0]   toplevel_execute_ctrl3_up_Prediction_BRANCH_HISTORY_lane1;
  reg        [1:0]    toplevel_execute_ctrl3_up_GSharePlugin_GSHARE_COUNTER_lane1_0;
  reg        [1:0]    toplevel_execute_ctrl3_up_GSharePlugin_GSHARE_COUNTER_lane1_1;
  reg        [1:0]    toplevel_execute_ctrl3_up_GSharePlugin_GSHARE_COUNTER_lane1_2;
  reg        [1:0]    toplevel_execute_ctrl3_up_GSharePlugin_GSHARE_COUNTER_lane1_3;
  reg        [3:0]    toplevel_execute_ctrl3_up_Prediction_ALIGNED_SLICES_BRANCH_lane1;
  reg        [3:0]    toplevel_execute_ctrl3_up_Prediction_ALIGNED_SLICES_TAKEN_lane1;
  reg        [31:0]   toplevel_execute_ctrl3_up_Prediction_ALIGNED_JUMPED_PC_lane1;
  reg                 toplevel_execute_ctrl3_up_Prediction_ALIGNED_JUMPED_lane1;
  reg        [31:0]   toplevel_execute_ctrl3_up_Decode_UOP_lane1;
  reg        [0:0]    toplevel_execute_ctrl3_up_LANE_AGE_lane0;
  reg        [4:0]    toplevel_execute_ctrl3_up_RD_PHYS_lane0;
  reg        [4:0]    toplevel_execute_ctrl3_up_RS2_PHYS_lane0;
  reg        [4:0]    toplevel_execute_ctrl3_up_RS1_PHYS_lane0;
  reg        [15:0]   toplevel_execute_ctrl3_up_Decode_UOP_ID_lane0;
  reg                 toplevel_execute_ctrl3_up_TRAP_lane0;
  reg        [31:0]   toplevel_execute_ctrl3_up_PC_lane0;
  reg        [0:0]    toplevel_execute_ctrl3_up_Decode_INSTRUCTION_SLICE_COUNT_lane0;
  reg        [11:0]   toplevel_execute_ctrl3_up_Prediction_BRANCH_HISTORY_lane0;
  reg        [1:0]    toplevel_execute_ctrl3_up_GSharePlugin_GSHARE_COUNTER_lane0_0;
  reg        [1:0]    toplevel_execute_ctrl3_up_GSharePlugin_GSHARE_COUNTER_lane0_1;
  reg        [1:0]    toplevel_execute_ctrl3_up_GSharePlugin_GSHARE_COUNTER_lane0_2;
  reg        [1:0]    toplevel_execute_ctrl3_up_GSharePlugin_GSHARE_COUNTER_lane0_3;
  reg        [3:0]    toplevel_execute_ctrl3_up_Prediction_ALIGNED_SLICES_BRANCH_lane0;
  reg        [3:0]    toplevel_execute_ctrl3_up_Prediction_ALIGNED_SLICES_TAKEN_lane0;
  reg        [31:0]   toplevel_execute_ctrl3_up_Prediction_ALIGNED_JUMPED_PC_lane0;
  reg                 toplevel_execute_ctrl3_up_Prediction_ALIGNED_JUMPED_lane0;
  reg        [31:0]   toplevel_execute_ctrl3_up_Decode_UOP_lane0;
  wire       [1:0]    toplevel_execute_ctrl1_down_AguPlugin_SIZE_lane0;
  wire                toplevel_execute_ctrl1_down_COMPLETED_lane1;
  wire       [4:0]    toplevel_execute_ctrl1_down_RD_PHYS_lane1;
  wire       [15:0]   toplevel_execute_ctrl1_down_Decode_UOP_ID_lane1;
  wire       [0:0]    toplevel_execute_ctrl1_down_Decode_INSTRUCTION_SLICE_COUNT_lane1;
  wire       [11:0]   toplevel_execute_ctrl1_down_Prediction_BRANCH_HISTORY_lane1;
  wire       [1:0]    toplevel_execute_ctrl1_down_GSharePlugin_GSHARE_COUNTER_lane1_0;
  wire       [1:0]    toplevel_execute_ctrl1_down_GSharePlugin_GSHARE_COUNTER_lane1_1;
  wire       [1:0]    toplevel_execute_ctrl1_down_GSharePlugin_GSHARE_COUNTER_lane1_2;
  wire       [1:0]    toplevel_execute_ctrl1_down_GSharePlugin_GSHARE_COUNTER_lane1_3;
  wire       [3:0]    toplevel_execute_ctrl1_down_Prediction_ALIGNED_SLICES_BRANCH_lane1;
  wire       [3:0]    toplevel_execute_ctrl1_down_Prediction_ALIGNED_SLICES_TAKEN_lane1;
  wire       [31:0]   toplevel_execute_ctrl1_down_Prediction_ALIGNED_JUMPED_PC_lane1;
  wire                toplevel_execute_ctrl1_down_Prediction_ALIGNED_JUMPED_lane1;
  wire                toplevel_execute_ctrl1_down_COMPLETED_lane0;
  wire       [4:0]    toplevel_execute_ctrl1_down_RD_PHYS_lane0;
  wire       [15:0]   toplevel_execute_ctrl1_down_Decode_UOP_ID_lane0;
  wire       [0:0]    toplevel_execute_ctrl1_down_Decode_INSTRUCTION_SLICE_COUNT_lane0;
  wire       [11:0]   toplevel_execute_ctrl1_down_Prediction_BRANCH_HISTORY_lane0;
  wire       [1:0]    toplevel_execute_ctrl1_down_GSharePlugin_GSHARE_COUNTER_lane0_0;
  wire       [1:0]    toplevel_execute_ctrl1_down_GSharePlugin_GSHARE_COUNTER_lane0_1;
  wire       [1:0]    toplevel_execute_ctrl1_down_GSharePlugin_GSHARE_COUNTER_lane0_2;
  wire       [1:0]    toplevel_execute_ctrl1_down_GSharePlugin_GSHARE_COUNTER_lane0_3;
  wire       [3:0]    toplevel_execute_ctrl1_down_Prediction_ALIGNED_SLICES_BRANCH_lane0;
  wire       [3:0]    toplevel_execute_ctrl1_down_Prediction_ALIGNED_SLICES_TAKEN_lane0;
  wire       [31:0]   toplevel_execute_ctrl1_down_Prediction_ALIGNED_JUMPED_PC_lane0;
  wire                toplevel_execute_ctrl1_down_Prediction_ALIGNED_JUMPED_lane0;
  wire                toplevel_execute_ctrl1_down_isReady;
  reg        [1:0]    toplevel_execute_ctrl2_up_late1_SrcPlugin_logic_SRC2_CTRL_lane1;
  reg        [0:0]    toplevel_execute_ctrl2_up_late1_SrcPlugin_logic_SRC1_CTRL_lane1;
  reg        [1:0]    toplevel_execute_ctrl2_up_late1_IntAluPlugin_ALU_BITWISE_CTRL_lane1;
  reg                 toplevel_execute_ctrl2_up_late1_IntAluPlugin_ALU_SLTX_lane1;
  reg                 toplevel_execute_ctrl2_up_late1_IntAluPlugin_ALU_ADD_SUB_lane1;
  reg        [1:0]    toplevel_execute_ctrl2_up_BranchPlugin_BRANCH_CTRL_lane1;
  reg                 toplevel_execute_ctrl2_up_BarrelShifterPlugin_SIGNED_lane1;
  reg                 toplevel_execute_ctrl2_up_BarrelShifterPlugin_LEFT_lane1;
  reg                 toplevel_execute_ctrl2_up_SrcStageables_UNSIGNED_lane1;
  reg                 toplevel_execute_ctrl2_up_BYPASSED_AT_3_lane1;
  reg                 toplevel_execute_ctrl2_up_SrcStageables_ZERO_lane1;
  reg                 toplevel_execute_ctrl2_up_SrcStageables_REVERT_lane1;
  reg        [1:0]    toplevel_execute_ctrl2_up_early1_IntAluPlugin_ALU_BITWISE_CTRL_lane1;
  reg                 toplevel_execute_ctrl2_up_early1_IntAluPlugin_ALU_SLTX_lane1;
  reg                 toplevel_execute_ctrl2_up_early1_IntAluPlugin_ALU_ADD_SUB_lane1;
  reg                 toplevel_execute_ctrl2_up_execute_lane1_logic_completions_onCtrl_2_ENABLE_lane1;
  reg                 toplevel_execute_ctrl2_up_execute_lane1_logic_completions_onCtrl_1_ENABLE_lane1;
  reg                 toplevel_execute_ctrl2_up_execute_lane1_logic_completions_onCtrl_0_ENABLE_lane1;
  reg                 toplevel_execute_ctrl2_up_COMPLETION_AT_4_lane1;
  reg                 toplevel_execute_ctrl2_up_COMPLETION_AT_3_lane1;
  reg                 toplevel_execute_ctrl2_up_COMPLETION_AT_2_lane1;
  reg                 toplevel_execute_ctrl2_up_lane1_integer_WriteBackPlugin_SEL_lane1;
  reg                 toplevel_execute_ctrl2_up_late1_BranchPlugin_SEL_lane1;
  reg                 toplevel_execute_ctrl2_up_late1_BarrelShifterPlugin_SEL_lane1;
  reg                 toplevel_execute_ctrl2_up_late1_IntAluPlugin_SEL_lane1;
  reg                 toplevel_execute_ctrl2_up_early1_BranchPlugin_SEL_lane1;
  reg                 toplevel_execute_ctrl2_up_early1_BarrelShifterPlugin_SEL_lane1;
  reg                 toplevel_execute_ctrl2_up_early1_IntAluPlugin_SEL_lane1;
  reg        [1:0]    toplevel_execute_ctrl2_up_late0_SrcPlugin_logic_SRC2_CTRL_lane0;
  reg        [0:0]    toplevel_execute_ctrl2_up_late0_SrcPlugin_logic_SRC1_CTRL_lane0;
  reg        [1:0]    toplevel_execute_ctrl2_up_late0_IntAluPlugin_ALU_BITWISE_CTRL_lane0;
  reg                 toplevel_execute_ctrl2_up_late0_IntAluPlugin_ALU_SLTX_lane0;
  reg                 toplevel_execute_ctrl2_up_late0_IntAluPlugin_ALU_ADD_SUB_lane0;
  reg        [2:0]    toplevel_execute_ctrl2_up_early0_EnvPlugin_OP_lane0;
  reg                 toplevel_execute_ctrl2_up_LsuPlugin_logic_LSU_PREFETCH_lane0;
  reg                 toplevel_execute_ctrl2_up_AguPlugin_FLOAT_lane0;
  reg                 toplevel_execute_ctrl2_up_AguPlugin_ATOMIC_lane0;
  reg                 toplevel_execute_ctrl2_up_AguPlugin_STORE_lane0;
  reg                 toplevel_execute_ctrl2_up_AguPlugin_LOAD_lane0;
  reg                 toplevel_execute_ctrl2_up_CsrAccessPlugin_CSR_CLEAR_lane0;
  reg                 toplevel_execute_ctrl2_up_CsrAccessPlugin_CSR_MASK_lane0;
  reg                 toplevel_execute_ctrl2_up_CsrAccessPlugin_CSR_IMM_lane0;
  reg                 toplevel_execute_ctrl2_up_DivPlugin_REM_lane0;
  reg                 toplevel_execute_ctrl2_up_RsUnsignedPlugin_RS2_SIGNED_lane0;
  reg                 toplevel_execute_ctrl2_up_RsUnsignedPlugin_RS1_SIGNED_lane0;
  reg        [1:0]    toplevel_execute_ctrl2_up_BranchPlugin_BRANCH_CTRL_lane0;
  reg                 toplevel_execute_ctrl2_up_BarrelShifterPlugin_SIGNED_lane0;
  reg                 toplevel_execute_ctrl2_up_BarrelShifterPlugin_LEFT_lane0;
  reg                 toplevel_execute_ctrl2_up_SrcStageables_UNSIGNED_lane0;
  reg                 toplevel_execute_ctrl2_up_BYPASSED_AT_3_lane0;
  reg        [1:0]    toplevel_execute_ctrl2_up_lane0_IntFormatPlugin_logic_WIDTH_ID_lane0;
  reg                 toplevel_execute_ctrl2_up_lane0_IntFormatPlugin_logic_SIGNED_lane0;
  reg                 toplevel_execute_ctrl2_up_SrcStageables_ZERO_lane0;
  reg                 toplevel_execute_ctrl2_up_SrcStageables_REVERT_lane0;
  reg        [1:0]    toplevel_execute_ctrl2_up_early0_IntAluPlugin_ALU_BITWISE_CTRL_lane0;
  reg                 toplevel_execute_ctrl2_up_early0_IntAluPlugin_ALU_SLTX_lane0;
  reg                 toplevel_execute_ctrl2_up_early0_IntAluPlugin_ALU_ADD_SUB_lane0;
  reg                 toplevel_execute_ctrl2_up_execute_lane0_logic_completions_onCtrl_2_ENABLE_lane0;
  reg                 toplevel_execute_ctrl2_up_execute_lane0_logic_completions_onCtrl_1_ENABLE_lane0;
  reg                 toplevel_execute_ctrl2_up_execute_lane0_logic_completions_onCtrl_0_ENABLE_lane0;
  reg                 toplevel_execute_ctrl2_up_COMPLETION_AT_4_lane0;
  reg                 toplevel_execute_ctrl2_up_COMPLETION_AT_3_lane0;
  reg                 toplevel_execute_ctrl2_up_COMPLETION_AT_2_lane0;
  reg                 toplevel_execute_ctrl2_up_lane0_integer_WriteBackPlugin_SEL_lane0;
  reg                 toplevel_execute_ctrl2_up_LsuPlugin_logic_FENCE_lane0;
  reg                 toplevel_execute_ctrl2_up_AguPlugin_SEL_lane0;
  reg                 toplevel_execute_ctrl2_up_CsrAccessPlugin_SEL_lane0;
  reg                 toplevel_execute_ctrl2_up_MulPlugin_HIGH_lane0;
  reg                 toplevel_execute_ctrl2_up_late0_BranchPlugin_SEL_lane0;
  reg                 toplevel_execute_ctrl2_up_late0_BarrelShifterPlugin_SEL_lane0;
  reg                 toplevel_execute_ctrl2_up_late0_IntAluPlugin_SEL_lane0;
  reg                 toplevel_execute_ctrl2_up_early0_EnvPlugin_SEL_lane0;
  reg                 toplevel_execute_ctrl2_up_early0_DivPlugin_SEL_lane0;
  reg                 toplevel_execute_ctrl2_up_early0_MulPlugin_SEL_lane0;
  reg                 toplevel_execute_ctrl2_up_early0_BranchPlugin_SEL_lane0;
  reg                 toplevel_execute_ctrl2_up_early0_BarrelShifterPlugin_SEL_lane0;
  reg                 toplevel_execute_ctrl2_up_early0_IntAluPlugin_SEL_lane0;
  reg                 toplevel_execute_ctrl2_up_MAY_FLUSH_PRECISE_3_lane1;
  reg                 toplevel_execute_ctrl2_up_MAY_FLUSH_PRECISE_3_lane0;
  reg        [31:0]   toplevel_execute_ctrl2_up_early1_SrcPlugin_SRC2_lane1;
  reg        [31:0]   toplevel_execute_ctrl2_up_early1_SrcPlugin_SRC1_lane1;
  reg        [31:0]   toplevel_execute_ctrl2_up_early0_SrcPlugin_SRC2_lane0;
  reg        [31:0]   toplevel_execute_ctrl2_up_early0_SrcPlugin_SRC1_lane0;
  reg        [1:0]    toplevel_execute_ctrl2_up_AguPlugin_SIZE_lane0;
  reg        [0:0]    toplevel_execute_ctrl2_up_LANE_AGE_lane1;
  reg        [4:0]    toplevel_execute_ctrl2_up_RS2_PHYS_lane1;
  reg        [4:0]    toplevel_execute_ctrl2_up_RS1_PHYS_lane1;
  reg        [15:0]   toplevel_execute_ctrl2_up_Decode_UOP_ID_lane1;
  reg        [31:0]   toplevel_execute_ctrl2_up_PC_lane1;
  reg        [0:0]    toplevel_execute_ctrl2_up_Decode_INSTRUCTION_SLICE_COUNT_lane1;
  reg        [11:0]   toplevel_execute_ctrl2_up_Prediction_BRANCH_HISTORY_lane1;
  reg        [1:0]    toplevel_execute_ctrl2_up_GSharePlugin_GSHARE_COUNTER_lane1_0;
  reg        [1:0]    toplevel_execute_ctrl2_up_GSharePlugin_GSHARE_COUNTER_lane1_1;
  reg        [1:0]    toplevel_execute_ctrl2_up_GSharePlugin_GSHARE_COUNTER_lane1_2;
  reg        [1:0]    toplevel_execute_ctrl2_up_GSharePlugin_GSHARE_COUNTER_lane1_3;
  reg        [3:0]    toplevel_execute_ctrl2_up_Prediction_ALIGNED_SLICES_BRANCH_lane1;
  reg        [3:0]    toplevel_execute_ctrl2_up_Prediction_ALIGNED_SLICES_TAKEN_lane1;
  reg        [31:0]   toplevel_execute_ctrl2_up_Prediction_ALIGNED_JUMPED_PC_lane1;
  reg                 toplevel_execute_ctrl2_up_Prediction_ALIGNED_JUMPED_lane1;
  reg        [31:0]   toplevel_execute_ctrl2_up_Decode_UOP_lane1;
  reg        [0:0]    toplevel_execute_ctrl2_up_LANE_AGE_lane0;
  reg        [4:0]    toplevel_execute_ctrl2_up_RS2_PHYS_lane0;
  reg        [4:0]    toplevel_execute_ctrl2_up_RS1_PHYS_lane0;
  reg        [15:0]   toplevel_execute_ctrl2_up_Decode_UOP_ID_lane0;
  reg        [31:0]   toplevel_execute_ctrl2_up_PC_lane0;
  reg        [0:0]    toplevel_execute_ctrl2_up_Decode_INSTRUCTION_SLICE_COUNT_lane0;
  reg        [11:0]   toplevel_execute_ctrl2_up_Prediction_BRANCH_HISTORY_lane0;
  reg        [1:0]    toplevel_execute_ctrl2_up_GSharePlugin_GSHARE_COUNTER_lane0_0;
  reg        [1:0]    toplevel_execute_ctrl2_up_GSharePlugin_GSHARE_COUNTER_lane0_1;
  reg        [1:0]    toplevel_execute_ctrl2_up_GSharePlugin_GSHARE_COUNTER_lane0_2;
  reg        [1:0]    toplevel_execute_ctrl2_up_GSharePlugin_GSHARE_COUNTER_lane0_3;
  reg        [3:0]    toplevel_execute_ctrl2_up_Prediction_ALIGNED_SLICES_BRANCH_lane0;
  reg        [3:0]    toplevel_execute_ctrl2_up_Prediction_ALIGNED_SLICES_TAKEN_lane0;
  reg        [31:0]   toplevel_execute_ctrl2_up_Prediction_ALIGNED_JUMPED_PC_lane0;
  reg                 toplevel_execute_ctrl2_up_Prediction_ALIGNED_JUMPED_lane0;
  reg        [31:0]   toplevel_execute_ctrl2_up_Decode_UOP_lane0;
  wire       [0:0]    toplevel_execute_ctrl0_down_execute_lane1_LAYER_SEL_lane1;
  wire                toplevel_execute_ctrl0_down_COMPLETED_lane1;
  wire       [4:0]    toplevel_execute_ctrl0_down_RD_PHYS_lane1;
  wire                toplevel_execute_ctrl0_down_TRAP_lane1;
  wire       [31:0]   toplevel_execute_ctrl0_down_PC_lane1;
  wire       [0:0]    toplevel_execute_ctrl0_down_Decode_INSTRUCTION_SLICE_COUNT_lane1;
  wire       [11:0]   toplevel_execute_ctrl0_down_Prediction_BRANCH_HISTORY_lane1;
  wire       [1:0]    toplevel_execute_ctrl0_down_GSharePlugin_GSHARE_COUNTER_lane1_0;
  wire       [1:0]    toplevel_execute_ctrl0_down_GSharePlugin_GSHARE_COUNTER_lane1_1;
  wire       [1:0]    toplevel_execute_ctrl0_down_GSharePlugin_GSHARE_COUNTER_lane1_2;
  wire       [1:0]    toplevel_execute_ctrl0_down_GSharePlugin_GSHARE_COUNTER_lane1_3;
  wire       [3:0]    toplevel_execute_ctrl0_down_Prediction_ALIGNED_SLICES_BRANCH_lane1;
  wire       [3:0]    toplevel_execute_ctrl0_down_Prediction_ALIGNED_SLICES_TAKEN_lane1;
  wire       [31:0]   toplevel_execute_ctrl0_down_Prediction_ALIGNED_JUMPED_PC_lane1;
  wire                toplevel_execute_ctrl0_down_Prediction_ALIGNED_JUMPED_lane1;
  wire       [31:0]   toplevel_execute_ctrl0_down_Decode_UOP_lane1;
  wire       [0:0]    toplevel_execute_ctrl0_down_execute_lane0_LAYER_SEL_lane0;
  wire                toplevel_execute_ctrl0_down_COMPLETED_lane0;
  wire       [4:0]    toplevel_execute_ctrl0_down_RD_PHYS_lane0;
  wire                toplevel_execute_ctrl0_down_TRAP_lane0;
  wire       [31:0]   toplevel_execute_ctrl0_down_PC_lane0;
  wire       [0:0]    toplevel_execute_ctrl0_down_Decode_INSTRUCTION_SLICE_COUNT_lane0;
  wire       [11:0]   toplevel_execute_ctrl0_down_Prediction_BRANCH_HISTORY_lane0;
  wire       [1:0]    toplevel_execute_ctrl0_down_GSharePlugin_GSHARE_COUNTER_lane0_0;
  wire       [1:0]    toplevel_execute_ctrl0_down_GSharePlugin_GSHARE_COUNTER_lane0_1;
  wire       [1:0]    toplevel_execute_ctrl0_down_GSharePlugin_GSHARE_COUNTER_lane0_2;
  wire       [1:0]    toplevel_execute_ctrl0_down_GSharePlugin_GSHARE_COUNTER_lane0_3;
  wire       [3:0]    toplevel_execute_ctrl0_down_Prediction_ALIGNED_SLICES_BRANCH_lane0;
  wire       [3:0]    toplevel_execute_ctrl0_down_Prediction_ALIGNED_SLICES_TAKEN_lane0;
  wire       [31:0]   toplevel_execute_ctrl0_down_Prediction_ALIGNED_JUMPED_PC_lane0;
  wire                toplevel_execute_ctrl0_down_Prediction_ALIGNED_JUMPED_lane0;
  reg        [1:0]    toplevel_execute_ctrl1_up_AguPlugin_SIZE_lane0;
  reg        [0:0]    toplevel_execute_ctrl1_up_execute_lane1_LAYER_SEL_lane1;
  reg                 toplevel_execute_ctrl1_up_COMPLETED_lane1;
  reg        [0:0]    toplevel_execute_ctrl1_up_LANE_AGE_lane1;
  reg        [4:0]    toplevel_execute_ctrl1_up_RS2_PHYS_lane1;
  reg        [4:0]    toplevel_execute_ctrl1_up_RS1_PHYS_lane1;
  reg        [15:0]   toplevel_execute_ctrl1_up_Decode_UOP_ID_lane1;
  reg                 toplevel_execute_ctrl1_up_TRAP_lane1;
  reg        [31:0]   toplevel_execute_ctrl1_up_PC_lane1;
  reg        [0:0]    toplevel_execute_ctrl1_up_Decode_INSTRUCTION_SLICE_COUNT_lane1;
  reg        [11:0]   toplevel_execute_ctrl1_up_Prediction_BRANCH_HISTORY_lane1;
  reg        [1:0]    toplevel_execute_ctrl1_up_GSharePlugin_GSHARE_COUNTER_lane1_0;
  reg        [1:0]    toplevel_execute_ctrl1_up_GSharePlugin_GSHARE_COUNTER_lane1_1;
  reg        [1:0]    toplevel_execute_ctrl1_up_GSharePlugin_GSHARE_COUNTER_lane1_2;
  reg        [1:0]    toplevel_execute_ctrl1_up_GSharePlugin_GSHARE_COUNTER_lane1_3;
  reg        [3:0]    toplevel_execute_ctrl1_up_Prediction_ALIGNED_SLICES_BRANCH_lane1;
  reg        [3:0]    toplevel_execute_ctrl1_up_Prediction_ALIGNED_SLICES_TAKEN_lane1;
  reg        [31:0]   toplevel_execute_ctrl1_up_Prediction_ALIGNED_JUMPED_PC_lane1;
  reg                 toplevel_execute_ctrl1_up_Prediction_ALIGNED_JUMPED_lane1;
  reg        [31:0]   toplevel_execute_ctrl1_up_Decode_UOP_lane1;
  reg        [0:0]    toplevel_execute_ctrl1_up_execute_lane0_LAYER_SEL_lane0;
  reg                 toplevel_execute_ctrl1_up_COMPLETED_lane0;
  reg        [0:0]    toplevel_execute_ctrl1_up_LANE_AGE_lane0;
  reg        [4:0]    toplevel_execute_ctrl1_up_RS2_PHYS_lane0;
  reg        [4:0]    toplevel_execute_ctrl1_up_RS1_PHYS_lane0;
  reg        [15:0]   toplevel_execute_ctrl1_up_Decode_UOP_ID_lane0;
  reg                 toplevel_execute_ctrl1_up_TRAP_lane0;
  reg        [31:0]   toplevel_execute_ctrl1_up_PC_lane0;
  reg        [0:0]    toplevel_execute_ctrl1_up_Decode_INSTRUCTION_SLICE_COUNT_lane0;
  reg        [11:0]   toplevel_execute_ctrl1_up_Prediction_BRANCH_HISTORY_lane0;
  reg        [1:0]    toplevel_execute_ctrl1_up_GSharePlugin_GSHARE_COUNTER_lane0_0;
  reg        [1:0]    toplevel_execute_ctrl1_up_GSharePlugin_GSHARE_COUNTER_lane0_1;
  reg        [1:0]    toplevel_execute_ctrl1_up_GSharePlugin_GSHARE_COUNTER_lane0_2;
  reg        [1:0]    toplevel_execute_ctrl1_up_GSharePlugin_GSHARE_COUNTER_lane0_3;
  reg        [3:0]    toplevel_execute_ctrl1_up_Prediction_ALIGNED_SLICES_BRANCH_lane0;
  reg        [3:0]    toplevel_execute_ctrl1_up_Prediction_ALIGNED_SLICES_TAKEN_lane0;
  reg        [31:0]   toplevel_execute_ctrl1_up_Prediction_ALIGNED_JUMPED_PC_lane0;
  reg                 toplevel_execute_ctrl1_up_Prediction_ALIGNED_JUMPED_lane0;
  reg        [31:0]   toplevel_execute_ctrl1_up_Decode_UOP_lane0;
  wire                toplevel_decode_ctrls_1_down_isReady;
  wire                toplevel_decode_ctrls_0_down_Prediction_ALIGN_REDO_1;
  wire       [3:0]    toplevel_decode_ctrls_0_down_Prediction_ALIGNED_SLICES_TAKEN_1;
  wire       [3:0]    toplevel_decode_ctrls_0_down_Prediction_ALIGNED_SLICES_BRANCH_1;
  wire       [31:0]   toplevel_decode_ctrls_0_down_Prediction_ALIGNED_JUMPED_PC_1;
  wire                toplevel_decode_ctrls_0_down_Prediction_ALIGNED_JUMPED_1;
  wire       [11:0]   toplevel_decode_ctrls_0_down_Prediction_BRANCH_HISTORY_1;
  wire       [1:0]    toplevel_decode_ctrls_0_down_GSharePlugin_GSHARE_COUNTER_1_0;
  wire       [1:0]    toplevel_decode_ctrls_0_down_GSharePlugin_GSHARE_COUNTER_1_1;
  wire       [1:0]    toplevel_decode_ctrls_0_down_GSharePlugin_GSHARE_COUNTER_1_2;
  wire       [1:0]    toplevel_decode_ctrls_0_down_GSharePlugin_GSHARE_COUNTER_1_3;
  wire       [0:0]    toplevel_decode_ctrls_0_down_Decode_INSTRUCTION_SLICE_COUNT_1;
  wire       [31:0]   toplevel_decode_ctrls_0_down_Decode_INSTRUCTION_RAW_1;
  wire                toplevel_decode_ctrls_0_down_Decode_DECOMPRESSION_FAULT_1;
  wire       [31:0]   toplevel_decode_ctrls_0_down_Decode_INSTRUCTION_1;
  wire                toplevel_decode_ctrls_0_down_Prediction_ALIGN_REDO_0;
  wire       [3:0]    toplevel_decode_ctrls_0_down_Prediction_ALIGNED_SLICES_TAKEN_0;
  wire       [3:0]    toplevel_decode_ctrls_0_down_Prediction_ALIGNED_SLICES_BRANCH_0;
  wire       [31:0]   toplevel_decode_ctrls_0_down_Prediction_ALIGNED_JUMPED_PC_0;
  wire                toplevel_decode_ctrls_0_down_Prediction_ALIGNED_JUMPED_0;
  wire       [11:0]   toplevel_decode_ctrls_0_down_Prediction_BRANCH_HISTORY_0;
  wire       [1:0]    toplevel_decode_ctrls_0_down_GSharePlugin_GSHARE_COUNTER_0_0;
  wire       [1:0]    toplevel_decode_ctrls_0_down_GSharePlugin_GSHARE_COUNTER_0_1;
  wire       [1:0]    toplevel_decode_ctrls_0_down_GSharePlugin_GSHARE_COUNTER_0_2;
  wire       [1:0]    toplevel_decode_ctrls_0_down_GSharePlugin_GSHARE_COUNTER_0_3;
  wire       [0:0]    toplevel_decode_ctrls_0_down_Decode_INSTRUCTION_SLICE_COUNT_0;
  wire       [31:0]   toplevel_decode_ctrls_0_down_Decode_INSTRUCTION_RAW_0;
  wire                toplevel_decode_ctrls_0_down_Decode_DECOMPRESSION_FAULT_0;
  wire       [31:0]   toplevel_decode_ctrls_0_down_Decode_INSTRUCTION_0;
  wire                toplevel_decode_ctrls_0_down_isValid;
  wire                toplevel_decode_ctrls_0_down_isReady;
  reg                 toplevel_decode_ctrls_1_up_Prediction_ALIGN_REDO_1;
  reg        [3:0]    toplevel_decode_ctrls_1_up_Prediction_ALIGNED_SLICES_TAKEN_1;
  reg        [3:0]    toplevel_decode_ctrls_1_up_Prediction_ALIGNED_SLICES_BRANCH_1;
  reg        [31:0]   toplevel_decode_ctrls_1_up_Prediction_ALIGNED_JUMPED_PC_1;
  reg                 toplevel_decode_ctrls_1_up_Prediction_ALIGNED_JUMPED_1;
  reg        [11:0]   toplevel_decode_ctrls_1_up_Prediction_BRANCH_HISTORY_1;
  reg        [1:0]    toplevel_decode_ctrls_1_up_GSharePlugin_GSHARE_COUNTER_1_0;
  reg        [1:0]    toplevel_decode_ctrls_1_up_GSharePlugin_GSHARE_COUNTER_1_1;
  reg        [1:0]    toplevel_decode_ctrls_1_up_GSharePlugin_GSHARE_COUNTER_1_2;
  reg        [1:0]    toplevel_decode_ctrls_1_up_GSharePlugin_GSHARE_COUNTER_1_3;
  reg        [9:0]    toplevel_decode_ctrls_1_up_Decode_DOP_ID_1;
  reg        [31:0]   toplevel_decode_ctrls_1_up_PC_1;
  reg        [0:0]    toplevel_decode_ctrls_1_up_Decode_INSTRUCTION_SLICE_COUNT_1;
  reg        [31:0]   toplevel_decode_ctrls_1_up_Decode_INSTRUCTION_RAW_1;
  reg                 toplevel_decode_ctrls_1_up_Decode_DECOMPRESSION_FAULT_1;
  reg        [31:0]   toplevel_decode_ctrls_1_up_Decode_INSTRUCTION_1;
  reg                 toplevel_decode_ctrls_1_up_Prediction_ALIGN_REDO_0;
  reg        [3:0]    toplevel_decode_ctrls_1_up_Prediction_ALIGNED_SLICES_TAKEN_0;
  reg        [3:0]    toplevel_decode_ctrls_1_up_Prediction_ALIGNED_SLICES_BRANCH_0;
  reg        [31:0]   toplevel_decode_ctrls_1_up_Prediction_ALIGNED_JUMPED_PC_0;
  reg                 toplevel_decode_ctrls_1_up_Prediction_ALIGNED_JUMPED_0;
  reg        [11:0]   toplevel_decode_ctrls_1_up_Prediction_BRANCH_HISTORY_0;
  reg        [1:0]    toplevel_decode_ctrls_1_up_GSharePlugin_GSHARE_COUNTER_0_0;
  reg        [1:0]    toplevel_decode_ctrls_1_up_GSharePlugin_GSHARE_COUNTER_0_1;
  reg        [1:0]    toplevel_decode_ctrls_1_up_GSharePlugin_GSHARE_COUNTER_0_2;
  reg        [1:0]    toplevel_decode_ctrls_1_up_GSharePlugin_GSHARE_COUNTER_0_3;
  reg        [9:0]    toplevel_decode_ctrls_1_up_Decode_DOP_ID_0;
  reg        [31:0]   toplevel_decode_ctrls_1_up_PC_0;
  reg        [0:0]    toplevel_decode_ctrls_1_up_Decode_INSTRUCTION_SLICE_COUNT_0;
  reg        [31:0]   toplevel_decode_ctrls_1_up_Decode_INSTRUCTION_RAW_0;
  reg                 toplevel_decode_ctrls_1_up_Decode_DECOMPRESSION_FAULT_0;
  reg        [31:0]   toplevel_decode_ctrls_1_up_Decode_INSTRUCTION_0;
  wire       [11:0]   fetch_logic_ctrls_1_down_Prediction_BRANCH_HISTORY;
  wire       [9:0]    fetch_logic_ctrls_1_down_Fetch_ID;
  wire                fetch_logic_ctrls_1_down_Fetch_PC_FAULT;
  wire                fetch_logic_ctrls_1_down_isValid;
  reg                 fetch_logic_ctrls_2_up_MMU_ACCESS_FAULT;
  reg                 fetch_logic_ctrls_2_up_MMU_PAGE_FAULT;
  reg                 fetch_logic_ctrls_2_up_MMU_ALLOW_EXECUTE;
  reg        [31:0]   fetch_logic_ctrls_2_up_MMU_TRANSLATED;
  reg                 fetch_logic_ctrls_2_up_MMU_REFILL;
  reg                 fetch_logic_ctrls_2_up_MMU_HAZARD;
  reg                 fetch_logic_ctrls_2_up_BtbPlugin_logic_chunksLogic_1_hitCalc_HIT;
  reg        [15:0]   fetch_logic_ctrls_2_up_BtbPlugin_logic_chunksLogic_1_readRsp_ENTRY_hash;
  reg        [0:0]    fetch_logic_ctrls_2_up_BtbPlugin_logic_chunksLogic_1_readRsp_ENTRY_sliceLow;
  reg        [30:0]   fetch_logic_ctrls_2_up_BtbPlugin_logic_chunksLogic_1_readRsp_ENTRY_pcTarget;
  reg                 fetch_logic_ctrls_2_up_BtbPlugin_logic_chunksLogic_1_readRsp_ENTRY_isBranch;
  reg                 fetch_logic_ctrls_2_up_BtbPlugin_logic_chunksLogic_1_readRsp_ENTRY_isPush;
  reg                 fetch_logic_ctrls_2_up_BtbPlugin_logic_chunksLogic_1_readRsp_ENTRY_isPop;
  reg                 fetch_logic_ctrls_2_up_BtbPlugin_logic_chunksLogic_0_hitCalc_HIT;
  reg        [15:0]   fetch_logic_ctrls_2_up_BtbPlugin_logic_chunksLogic_0_readRsp_ENTRY_hash;
  reg        [0:0]    fetch_logic_ctrls_2_up_BtbPlugin_logic_chunksLogic_0_readRsp_ENTRY_sliceLow;
  reg        [30:0]   fetch_logic_ctrls_2_up_BtbPlugin_logic_chunksLogic_0_readRsp_ENTRY_pcTarget;
  reg                 fetch_logic_ctrls_2_up_BtbPlugin_logic_chunksLogic_0_readRsp_ENTRY_isBranch;
  reg                 fetch_logic_ctrls_2_up_BtbPlugin_logic_chunksLogic_0_readRsp_ENTRY_isPush;
  reg                 fetch_logic_ctrls_2_up_BtbPlugin_logic_chunksLogic_0_readRsp_ENTRY_isPop;
  reg        [1:0]    fetch_logic_ctrls_2_up_GSharePlugin_GSHARE_COUNTER_0;
  reg        [1:0]    fetch_logic_ctrls_2_up_GSharePlugin_GSHARE_COUNTER_1;
  reg        [1:0]    fetch_logic_ctrls_2_up_GSharePlugin_GSHARE_COUNTER_2;
  reg        [1:0]    fetch_logic_ctrls_2_up_GSharePlugin_GSHARE_COUNTER_3;
  reg                 fetch_logic_ctrls_2_up_FetchL1Plugin_logic_WAYS_HIT;
  reg                 fetch_logic_ctrls_2_up_MMU_BYPASS_TRANSLATION;
  reg                 fetch_logic_ctrls_2_up_FetchL1Plugin_logic_WAYS_HITS_0;
  reg                 fetch_logic_ctrls_2_up_FetchL1Plugin_logic_WAYS_HITS_1;
  reg                 fetch_logic_ctrls_2_up_FetchL1Plugin_logic_HAZARD;
  reg        [63:0]   fetch_logic_ctrls_2_up_FetchL1Plugin_logic_BANKS_MUXES_0;
  reg        [63:0]   fetch_logic_ctrls_2_up_FetchL1Plugin_logic_BANKS_MUXES_1;
  reg        [0:0]    fetch_logic_ctrls_2_up_FetchL1Plugin_logic_PLRU_BYPASSED_0;
  reg                 fetch_logic_ctrls_2_up_FetchL1Plugin_logic_WAYS_TAGS_0_loaded;
  reg                 fetch_logic_ctrls_2_up_FetchL1Plugin_logic_WAYS_TAGS_0_error;
  reg        [19:0]   fetch_logic_ctrls_2_up_FetchL1Plugin_logic_WAYS_TAGS_0_address;
  reg                 fetch_logic_ctrls_2_up_FetchL1Plugin_logic_WAYS_TAGS_1_loaded;
  reg                 fetch_logic_ctrls_2_up_FetchL1Plugin_logic_WAYS_TAGS_1_error;
  reg        [19:0]   fetch_logic_ctrls_2_up_FetchL1Plugin_logic_WAYS_TAGS_1_address;
  reg        [11:0]   fetch_logic_ctrls_2_up_Prediction_BRANCH_HISTORY;
  reg        [9:0]    fetch_logic_ctrls_2_up_Fetch_ID;
  reg                 fetch_logic_ctrls_2_up_Fetch_PC_FAULT;
  reg        [31:0]   fetch_logic_ctrls_2_up_Fetch_WORD_PC;
  wire                fetch_logic_ctrls_0_down_Fetch_PC_FAULT;
  wire                fetch_logic_ctrls_0_down_isValid;
  reg        [1:0]    fetch_logic_ctrls_1_up_BtbPlugin_logic_readCmd_HAZARDS;
  reg                 fetch_logic_ctrls_1_up_GSharePlugin_logic_BYPASS_valid;
  reg        [11:0]   fetch_logic_ctrls_1_up_GSharePlugin_logic_BYPASS_payload_address;
  reg        [1:0]    fetch_logic_ctrls_1_up_GSharePlugin_logic_BYPASS_payload_data_0;
  reg        [1:0]    fetch_logic_ctrls_1_up_GSharePlugin_logic_BYPASS_payload_data_1;
  reg        [1:0]    fetch_logic_ctrls_1_up_GSharePlugin_logic_BYPASS_payload_data_2;
  reg        [1:0]    fetch_logic_ctrls_1_up_GSharePlugin_logic_BYPASS_payload_data_3;
  reg        [11:0]   fetch_logic_ctrls_1_up_Prediction_BRANCH_HISTORY;
  reg        [11:0]   fetch_logic_ctrls_1_up_GSharePlugin_logic_HASH;
  reg        [5:0]    fetch_logic_ctrls_1_up_FetchL1Plugin_logic_cmd_TAGS_UPDATE_ADDRESS;
  reg                 fetch_logic_ctrls_1_up_FetchL1Plugin_logic_cmd_TAGS_UPDATE;
  reg        [0:0]    fetch_logic_ctrls_1_up_FetchL1Plugin_logic_cmd_PLRU_BYPASS_DATA_0;
  reg                 fetch_logic_ctrls_1_up_FetchL1Plugin_logic_cmd_PLRU_BYPASS_VALID;
  reg                 _zz_1;
  reg        [9:0]    fetch_logic_ctrls_1_up_Fetch_ID;
  reg                 fetch_logic_ctrls_1_up_Fetch_PC_FAULT;
  reg        [31:0]   fetch_logic_ctrls_1_up_Fetch_WORD_PC;
  reg                 fetch_logic_ctrls_2_up_valid;
  wire                toplevel_decode_ctrls_1_down_valid;
  reg                 fetch_logic_ctrls_1_down_valid;
  wire                toplevel_decode_ctrls_0_down_valid;
  reg                 fetch_logic_ctrls_0_down_valid;
  wire                toplevel_execute_ctrl0_up_ready;
  wire                toplevel_execute_ctrl0_down_ready;
  wire                toplevel_execute_ctrl1_up_ready;
  wire                toplevel_execute_ctrl1_down_ready;
  wire                toplevel_execute_ctrl2_up_ready;
  wire                toplevel_execute_ctrl2_down_ready;
  wire                toplevel_execute_ctrl3_up_ready;
  wire                toplevel_execute_ctrl3_down_ready;
  wire                fetch_logic_ctrls_0_down_ready;
  wire                toplevel_execute_ctrl4_up_ready;
  wire                toplevel_decode_ctrls_0_up_ready;
  wire                fetch_logic_ctrls_1_up_cancel;
  wire                toplevel_execute_ctrl4_down_ready;
  reg                 toplevel_decode_ctrls_0_down_ready;
  wire                fetch_logic_ctrls_1_down_ready;
  wire                toplevel_execute_ctrl5_up_ready;
  wire                fetch_logic_ctrls_2_up_ready;
  wire                fetch_logic_ctrls_2_up_cancel;
  wire                toplevel_execute_ctrl4_down_AguPlugin_ATOMIC_lane0;
  wire       [11:0]   toplevel_execute_ctrl4_down_Decode_STORE_ID_lane0;
  wire       [31:0]   toplevel_execute_ctrl4_down_MMU_TRANSLATED_lane0;
  wire       [1:0]    toplevel_execute_ctrl4_down_AguPlugin_SIZE_lane0;
  wire                toplevel_execute_ctrl4_down_LsuPlugin_logic_LSU_PREFETCH_lane0;
  wire                toplevel_execute_ctrl4_down_AguPlugin_LOAD_lane0;
  wire                toplevel_execute_ctrl5_down_ready;
  reg                 toplevel_execute_ctrl2_up_TRAP_lane1;
  wire                toplevel_execute_ctrl2_up_COMMIT_lane1;
  wire       [0:0]    toplevel_execute_ctrl5_down_LANE_AGE_lane1;
  wire                toplevel_execute_ctrl4_down_RD_ENABLE_lane1;
  reg                 toplevel_execute_ctrl4_RD_ENABLE_lane1_bypass;
  reg                 toplevel_execute_ctrl4_LANE_SEL_lane1_bypass;
  wire                toplevel_execute_ctrl3_down_RD_ENABLE_lane1;
  reg                 toplevel_execute_ctrl3_RD_ENABLE_lane1_bypass;
  reg                 toplevel_execute_ctrl3_LANE_SEL_lane1_bypass;
  wire                toplevel_execute_ctrl2_down_RD_ENABLE_lane1;
  reg                 toplevel_execute_ctrl2_RD_ENABLE_lane1_bypass;
  reg                 toplevel_execute_ctrl2_LANE_SEL_lane1_bypass;
  wire       [0:0]    toplevel_execute_ctrl2_down_LANE_AGE_lane1;
  wire                toplevel_execute_ctrl1_down_RD_ENABLE_lane1;
  reg                 toplevel_execute_ctrl1_RD_ENABLE_lane1_bypass;
  wire                toplevel_execute_ctrl1_down_LANE_SEL_lane1;
  reg                 toplevel_execute_ctrl1_LANE_SEL_lane1_bypass;
  wire       [0:0]    toplevel_execute_ctrl1_down_LANE_AGE_lane1;
  wire                toplevel_execute_ctrl0_down_RD_ENABLE_lane1;
  reg                 toplevel_execute_ctrl0_RD_ENABLE_lane1_bypass;
  reg                 toplevel_execute_ctrl0_LANE_SEL_lane1_bypass;
  wire       [0:0]    toplevel_execute_ctrl0_down_LANE_AGE_lane1;
  wire                toplevel_execute_ctrl1_down_TRAP_lane1;
  wire       [1:0]    toplevel_execute_ctrl1_down_late1_SrcPlugin_logic_SRC2_CTRL_lane1;
  wire       [0:0]    toplevel_execute_ctrl1_down_late1_SrcPlugin_logic_SRC1_CTRL_lane1;
  wire       [1:0]    toplevel_execute_ctrl1_down_late1_IntAluPlugin_ALU_BITWISE_CTRL_lane1;
  wire                toplevel_execute_ctrl1_down_late1_IntAluPlugin_ALU_SLTX_lane1;
  wire                toplevel_execute_ctrl1_down_late1_IntAluPlugin_ALU_ADD_SUB_lane1;
  wire       [1:0]    toplevel_execute_ctrl1_down_BranchPlugin_BRANCH_CTRL_lane1;
  wire                toplevel_execute_ctrl1_down_BarrelShifterPlugin_SIGNED_lane1;
  wire                toplevel_execute_ctrl1_down_BarrelShifterPlugin_LEFT_lane1;
  wire                toplevel_execute_ctrl1_down_SrcStageables_UNSIGNED_lane1;
  wire                toplevel_execute_ctrl1_down_BYPASSED_AT_3_lane1;
  wire                toplevel_execute_ctrl1_down_lane1_IntFormatPlugin_logic_SIGNED_lane1;
  wire                toplevel_execute_ctrl1_down_SrcStageables_ZERO_lane1;
  wire                toplevel_execute_ctrl1_down_SrcStageables_REVERT_lane1;
  wire       [1:0]    toplevel_execute_ctrl1_down_early1_IntAluPlugin_ALU_BITWISE_CTRL_lane1;
  wire                toplevel_execute_ctrl1_down_early1_IntAluPlugin_ALU_SLTX_lane1;
  wire                toplevel_execute_ctrl1_down_early1_IntAluPlugin_ALU_ADD_SUB_lane1;
  reg                 toplevel_execute_ctrl1_down_execute_lane1_logic_completions_onCtrl_2_ENABLE_lane1;
  reg                 toplevel_execute_ctrl1_down_execute_lane1_logic_completions_onCtrl_1_ENABLE_lane1;
  reg                 toplevel_execute_ctrl1_down_execute_lane1_logic_completions_onCtrl_0_ENABLE_lane1;
  reg                 toplevel_execute_ctrl1_down_COMPLETION_AT_4_lane1;
  reg                 toplevel_execute_ctrl1_down_COMPLETION_AT_3_lane1;
  reg                 toplevel_execute_ctrl1_down_COMPLETION_AT_2_lane1;
  reg                 toplevel_execute_ctrl1_down_lane1_integer_WriteBackPlugin_SEL_lane1;
  reg                 toplevel_execute_ctrl1_down_late1_BranchPlugin_SEL_lane1;
  reg                 toplevel_execute_ctrl1_down_late1_BarrelShifterPlugin_SEL_lane1;
  reg                 toplevel_execute_ctrl1_down_late1_IntAluPlugin_SEL_lane1;
  reg                 toplevel_execute_ctrl1_down_early1_BranchPlugin_SEL_lane1;
  reg                 toplevel_execute_ctrl1_down_early1_BarrelShifterPlugin_SEL_lane1;
  reg                 toplevel_execute_ctrl1_down_early1_IntAluPlugin_SEL_lane1;
  wire       [0:0]    toplevel_execute_ctrl1_down_execute_lane1_LAYER_SEL_lane1;
  wire                toplevel_execute_ctrl4_down_execute_lane1_logic_completions_onCtrl_2_ENABLE_lane1;
  wire                toplevel_execute_ctrl3_down_TRAP_lane1;
  wire                toplevel_execute_ctrl3_down_execute_lane1_logic_completions_onCtrl_1_ENABLE_lane1;
  wire                toplevel_execute_ctrl2_down_TRAP_lane1;
  wire                toplevel_execute_ctrl2_down_execute_lane1_logic_completions_onCtrl_0_ENABLE_lane1;
  reg        [31:0]   toplevel_execute_ctrl3_up_integer_RS2_lane1;
  wire       [31:0]   toplevel_execute_ctrl3_integer_RS2_lane1_bypass;
  wire       [4:0]    toplevel_execute_ctrl3_down_RS2_PHYS_lane1;
  reg        [31:0]   toplevel_execute_ctrl2_up_integer_RS2_lane1;
  wire       [31:0]   toplevel_execute_ctrl2_down_integer_RS2_lane1;
  wire       [31:0]   toplevel_execute_ctrl2_integer_RS2_lane1_bypass;
  wire       [4:0]    toplevel_execute_ctrl2_down_RS2_PHYS_lane1;
  wire       [4:0]    toplevel_execute_ctrl1_down_RS2_PHYS_lane1;
  wire       [4:0]    toplevel_execute_ctrl0_down_RS2_PHYS_lane1;
  reg        [31:0]   toplevel_execute_ctrl3_up_integer_RS1_lane1;
  wire       [31:0]   toplevel_execute_ctrl3_integer_RS1_lane1_bypass;
  wire       [4:0]    toplevel_execute_ctrl3_down_RS1_PHYS_lane1;
  reg        [31:0]   toplevel_execute_ctrl2_up_integer_RS1_lane1;
  wire       [31:0]   toplevel_execute_ctrl2_down_integer_RS1_lane1;
  wire       [31:0]   toplevel_execute_ctrl2_integer_RS1_lane1_bypass;
  wire       [4:0]    toplevel_execute_ctrl2_down_RS1_PHYS_lane1;
  wire       [4:0]    toplevel_execute_ctrl1_down_RS1_PHYS_lane1;
  wire       [0:0]    toplevel_execute_ctrl5_down_LANE_AGE_lane0;
  wire                toplevel_execute_ctrl4_down_RD_ENABLE_lane0;
  reg                 toplevel_execute_ctrl4_RD_ENABLE_lane0_bypass;
  reg                 toplevel_execute_ctrl4_LANE_SEL_lane0_bypass;
  wire                toplevel_execute_ctrl3_down_RD_ENABLE_lane0;
  reg                 toplevel_execute_ctrl3_RD_ENABLE_lane0_bypass;
  reg                 toplevel_execute_ctrl3_LANE_SEL_lane0_bypass;
  wire                toplevel_execute_ctrl2_down_RD_ENABLE_lane0;
  reg                 toplevel_execute_ctrl2_RD_ENABLE_lane0_bypass;
  reg                 toplevel_execute_ctrl2_LANE_SEL_lane0_bypass;
  wire                toplevel_execute_ctrl1_down_RD_ENABLE_lane0;
  reg                 toplevel_execute_ctrl1_RD_ENABLE_lane0_bypass;
  wire                toplevel_execute_ctrl1_down_LANE_SEL_lane0;
  reg                 toplevel_execute_ctrl1_LANE_SEL_lane0_bypass;
  wire       [0:0]    toplevel_execute_ctrl1_down_LANE_AGE_lane0;
  wire                toplevel_execute_ctrl0_down_RD_ENABLE_lane0;
  reg                 toplevel_execute_ctrl0_RD_ENABLE_lane0_bypass;
  reg                 toplevel_execute_ctrl0_LANE_SEL_lane0_bypass;
  wire       [0:0]    toplevel_execute_ctrl0_down_LANE_AGE_lane0;
  wire                toplevel_execute_ctrl1_down_TRAP_lane0;
  wire       [1:0]    toplevel_execute_ctrl1_down_late0_SrcPlugin_logic_SRC2_CTRL_lane0;
  wire       [0:0]    toplevel_execute_ctrl1_down_late0_SrcPlugin_logic_SRC1_CTRL_lane0;
  wire       [1:0]    toplevel_execute_ctrl1_down_late0_IntAluPlugin_ALU_BITWISE_CTRL_lane0;
  wire                toplevel_execute_ctrl1_down_late0_IntAluPlugin_ALU_SLTX_lane0;
  wire                toplevel_execute_ctrl1_down_late0_IntAluPlugin_ALU_ADD_SUB_lane0;
  wire       [2:0]    toplevel_execute_ctrl1_down_early0_EnvPlugin_OP_lane0;
  wire                toplevel_execute_ctrl1_down_LsuPlugin_logic_LSU_PREFETCH_lane0;
  wire                toplevel_execute_ctrl1_down_AguPlugin_FLOAT_lane0;
  wire                toplevel_execute_ctrl1_down_AguPlugin_ATOMIC_lane0;
  wire                toplevel_execute_ctrl1_down_AguPlugin_STORE_lane0;
  wire                toplevel_execute_ctrl1_down_AguPlugin_LOAD_lane0;
  wire                toplevel_execute_ctrl1_down_CsrAccessPlugin_CSR_CLEAR_lane0;
  wire                toplevel_execute_ctrl1_down_CsrAccessPlugin_CSR_MASK_lane0;
  wire                toplevel_execute_ctrl1_down_CsrAccessPlugin_CSR_IMM_lane0;
  wire                toplevel_execute_ctrl1_down_DivPlugin_REM_lane0;
  wire                toplevel_execute_ctrl1_down_RsUnsignedPlugin_RS2_SIGNED_lane0;
  wire                toplevel_execute_ctrl1_down_RsUnsignedPlugin_RS1_SIGNED_lane0;
  wire       [1:0]    toplevel_execute_ctrl1_down_BranchPlugin_BRANCH_CTRL_lane0;
  wire                toplevel_execute_ctrl1_down_BarrelShifterPlugin_SIGNED_lane0;
  wire                toplevel_execute_ctrl1_down_BarrelShifterPlugin_LEFT_lane0;
  wire                toplevel_execute_ctrl1_down_SrcStageables_UNSIGNED_lane0;
  wire                toplevel_execute_ctrl1_down_BYPASSED_AT_3_lane0;
  wire       [1:0]    toplevel_execute_ctrl1_down_lane0_IntFormatPlugin_logic_WIDTH_ID_lane0;
  wire                toplevel_execute_ctrl1_down_lane0_IntFormatPlugin_logic_SIGNED_lane0;
  wire                toplevel_execute_ctrl1_down_SrcStageables_ZERO_lane0;
  wire                toplevel_execute_ctrl1_down_SrcStageables_REVERT_lane0;
  wire       [1:0]    toplevel_execute_ctrl1_down_early0_IntAluPlugin_ALU_BITWISE_CTRL_lane0;
  wire                toplevel_execute_ctrl1_down_early0_IntAluPlugin_ALU_SLTX_lane0;
  wire                toplevel_execute_ctrl1_down_early0_IntAluPlugin_ALU_ADD_SUB_lane0;
  reg                 toplevel_execute_ctrl1_down_execute_lane0_logic_completions_onCtrl_2_ENABLE_lane0;
  reg                 toplevel_execute_ctrl1_down_execute_lane0_logic_completions_onCtrl_1_ENABLE_lane0;
  reg                 toplevel_execute_ctrl1_down_execute_lane0_logic_completions_onCtrl_0_ENABLE_lane0;
  reg                 toplevel_execute_ctrl1_down_COMPLETION_AT_4_lane0;
  reg                 toplevel_execute_ctrl1_down_COMPLETION_AT_3_lane0;
  reg                 toplevel_execute_ctrl1_down_COMPLETION_AT_2_lane0;
  reg                 toplevel_execute_ctrl1_down_lane0_integer_WriteBackPlugin_SEL_lane0;
  reg                 toplevel_execute_ctrl1_down_LsuPlugin_logic_FENCE_lane0;
  reg                 toplevel_execute_ctrl1_down_AguPlugin_SEL_lane0;
  reg                 toplevel_execute_ctrl1_down_CsrAccessPlugin_SEL_lane0;
  reg                 toplevel_execute_ctrl1_down_MulPlugin_HIGH_lane0;
  reg                 toplevel_execute_ctrl1_down_late0_BranchPlugin_SEL_lane0;
  reg                 toplevel_execute_ctrl1_down_late0_BarrelShifterPlugin_SEL_lane0;
  reg                 toplevel_execute_ctrl1_down_late0_IntAluPlugin_SEL_lane0;
  reg                 toplevel_execute_ctrl1_down_early0_EnvPlugin_SEL_lane0;
  reg                 toplevel_execute_ctrl1_down_early0_DivPlugin_SEL_lane0;
  reg                 toplevel_execute_ctrl1_down_early0_MulPlugin_SEL_lane0;
  reg                 toplevel_execute_ctrl1_down_early0_BranchPlugin_SEL_lane0;
  reg                 toplevel_execute_ctrl1_down_early0_BarrelShifterPlugin_SEL_lane0;
  reg                 toplevel_execute_ctrl1_down_early0_IntAluPlugin_SEL_lane0;
  wire       [0:0]    toplevel_execute_ctrl1_down_execute_lane0_LAYER_SEL_lane0;
  wire                toplevel_execute_ctrl4_down_execute_lane0_logic_completions_onCtrl_2_ENABLE_lane0;
  wire                toplevel_execute_ctrl3_down_TRAP_lane0;
  wire                toplevel_execute_ctrl3_down_execute_lane0_logic_completions_onCtrl_1_ENABLE_lane0;
  wire                toplevel_execute_ctrl2_down_execute_lane0_logic_completions_onCtrl_0_ENABLE_lane0;
  reg        [31:0]   toplevel_execute_ctrl3_up_integer_RS2_lane0;
  wire       [31:0]   toplevel_execute_ctrl3_integer_RS2_lane0_bypass;
  wire       [4:0]    toplevel_execute_ctrl3_down_RS2_PHYS_lane0;
  wire       [31:0]   toplevel_execute_ctrl2_down_integer_RS2_lane0;
  wire       [31:0]   toplevel_execute_ctrl2_integer_RS2_lane0_bypass;
  wire       [4:0]    toplevel_execute_ctrl2_down_RS2_PHYS_lane0;
  wire       [4:0]    toplevel_execute_ctrl1_down_RS2_PHYS_lane0;
  wire       [4:0]    toplevel_execute_ctrl0_down_RS2_PHYS_lane0;
  reg        [31:0]   toplevel_execute_ctrl3_up_integer_RS1_lane0;
  wire       [31:0]   toplevel_execute_ctrl3_integer_RS1_lane0_bypass;
  wire       [4:0]    toplevel_execute_ctrl3_down_RS1_PHYS_lane0;
  wire       [31:0]   toplevel_execute_ctrl2_down_integer_RS1_lane0;
  wire       [31:0]   toplevel_execute_ctrl2_integer_RS1_lane0_bypass;
  wire       [4:0]    toplevel_execute_ctrl2_down_RS1_PHYS_lane0;
  wire       [31:0]   toplevel_execute_ctrl5_down_lane1_integer_WriteBackPlugin_logic_DATA_lane1;
  wire       [31:0]   toplevel_execute_ctrl5_down_lane0_integer_WriteBackPlugin_logic_DATA_lane0;
  wire       [4:0]    toplevel_execute_ctrl5_down_RD_PHYS_lane1;
  reg                 toplevel_execute_ctrl5_up_RD_ENABLE_lane1;
  reg                 toplevel_execute_ctrl5_up_LANE_SEL_lane1;
  wire       [4:0]    toplevel_execute_ctrl5_down_RD_PHYS_lane0;
  reg                 toplevel_execute_ctrl5_up_RD_ENABLE_lane0;
  reg                 toplevel_execute_ctrl5_up_LANE_SEL_lane0;
  wire       [4:0]    toplevel_execute_ctrl3_down_RD_PHYS_lane1;
  wire       [4:0]    toplevel_execute_ctrl3_down_RD_PHYS_lane0;
  wire       [4:0]    toplevel_execute_ctrl2_down_RD_PHYS_lane1;
  wire       [4:0]    toplevel_execute_ctrl1_down_RS1_PHYS_lane0;
  wire       [4:0]    toplevel_execute_ctrl0_down_RS1_PHYS_lane0;
  reg                 _zz_2;
  wire                toplevel_execute_ctrl3_down_CsrAccessPlugin_SEL_lane0;
  wire       [4:0]    toplevel_execute_ctrl2_down_RD_PHYS_lane0;
  wire                toplevel_execute_ctrl2_down_CsrAccessPlugin_CSR_CLEAR_lane0;
  wire                toplevel_execute_ctrl2_down_CsrAccessPlugin_CSR_MASK_lane0;
  wire                toplevel_execute_ctrl2_down_CsrAccessPlugin_CSR_IMM_lane0;
  wire                toplevel_execute_ctrl2_down_CsrAccessPlugin_SEL_lane0;
  wire                fetch_logic_ctrls_0_up_isFiring;
  reg        [9:0]    fetch_logic_ctrls_0_up_Fetch_ID;
  wire                fetch_logic_ctrls_0_up_Fetch_PC_FAULT;
  wire       [31:0]   fetch_logic_ctrls_0_up_Fetch_WORD_PC;
  reg                 fetch_logic_ctrls_0_up_ready;
  wire                fetch_logic_ctrls_0_up_valid;
  reg                 fetch_logic_ctrls_1_down_MMU_ACCESS_FAULT;
  reg                 fetch_logic_ctrls_1_down_MMU_PAGE_FAULT;
  reg                 fetch_logic_ctrls_1_down_MMU_ALLOW_WRITE;
  reg                 fetch_logic_ctrls_1_down_MMU_ALLOW_READ;
  reg                 fetch_logic_ctrls_1_down_MMU_ALLOW_EXECUTE;
  reg        [31:0]   fetch_logic_ctrls_1_down_MMU_TRANSLATED;
  reg                 fetch_logic_ctrls_1_down_MMU_REFILL;
  reg                 fetch_logic_ctrls_1_down_MMU_HAZARD;
  wire       [0:0]    fetch_logic_ctrls_1_down_MMU_L1_HITS;
  wire       [0:0]    fetch_logic_ctrls_1_down_MMU_L1_HITS_PRE_VALID;
  wire                fetch_logic_ctrls_1_down_MMU_L1_ENTRIES_0_valid;
  wire       [3:0]    fetch_logic_ctrls_1_down_MMU_L1_ENTRIES_0_virtualAddress;
  wire       [9:0]    fetch_logic_ctrls_1_down_MMU_L1_ENTRIES_0_physicalAddress;
  wire                fetch_logic_ctrls_1_down_MMU_L1_ENTRIES_0_allowRead;
  wire                fetch_logic_ctrls_1_down_MMU_L1_ENTRIES_0_allowWrite;
  wire                fetch_logic_ctrls_1_down_MMU_L1_ENTRIES_0_allowExecute;
  wire                fetch_logic_ctrls_1_down_MMU_L1_ENTRIES_0_allowUser;
  reg        [1:0]    fetch_logic_ctrls_1_down_MMU_L0_HITS;
  reg        [1:0]    fetch_logic_ctrls_1_down_MMU_L0_HITS_PRE_VALID;
  wire                fetch_logic_ctrls_1_down_MMU_L0_ENTRIES_0_valid;
  wire       [13:0]   fetch_logic_ctrls_1_down_MMU_L0_ENTRIES_0_virtualAddress;
  wire       [19:0]   fetch_logic_ctrls_1_down_MMU_L0_ENTRIES_0_physicalAddress;
  wire                fetch_logic_ctrls_1_down_MMU_L0_ENTRIES_0_allowRead;
  wire                fetch_logic_ctrls_1_down_MMU_L0_ENTRIES_0_allowWrite;
  wire                fetch_logic_ctrls_1_down_MMU_L0_ENTRIES_0_allowExecute;
  wire                fetch_logic_ctrls_1_down_MMU_L0_ENTRIES_0_allowUser;
  wire                fetch_logic_ctrls_1_down_MMU_L0_ENTRIES_1_valid;
  wire       [13:0]   fetch_logic_ctrls_1_down_MMU_L0_ENTRIES_1_virtualAddress;
  wire       [19:0]   fetch_logic_ctrls_1_down_MMU_L0_ENTRIES_1_physicalAddress;
  wire                fetch_logic_ctrls_1_down_MMU_L0_ENTRIES_1_allowRead;
  wire                fetch_logic_ctrls_1_down_MMU_L0_ENTRIES_1_allowWrite;
  wire                fetch_logic_ctrls_1_down_MMU_L0_ENTRIES_1_allowExecute;
  wire                fetch_logic_ctrls_1_down_MMU_L0_ENTRIES_1_allowUser;
  wire       [31:0]   toplevel_execute_ctrl3_down_MMU_WAYS_PHYSICAL_lane0_0;
  wire       [31:0]   toplevel_execute_ctrl3_down_MMU_WAYS_PHYSICAL_lane0_1;
  wire       [31:0]   toplevel_execute_ctrl3_down_MMU_WAYS_PHYSICAL_lane0_2;
  wire       [2:0]    toplevel_execute_ctrl3_down_MMU_WAYS_OH_lane0;
  wire                toplevel_execute_ctrl3_down_MMU_BYPASS_TRANSLATION_lane0;
  reg                 toplevel_execute_ctrl3_down_MMU_ALLOW_EXECUTE_lane0;
  wire                toplevel_execute_ctrl3_down_LsuPlugin_logic_FORCE_PHYSICAL_lane0;
  wire       [0:0]    toplevel_execute_ctrl3_down_MMU_L1_HITS_lane0;
  wire       [0:0]    toplevel_execute_ctrl3_down_MMU_L1_HITS_PRE_VALID_lane0;
  wire                toplevel_execute_ctrl3_down_MMU_L1_ENTRIES_lane0_0_valid;
  wire       [3:0]    toplevel_execute_ctrl3_down_MMU_L1_ENTRIES_lane0_0_virtualAddress;
  wire       [9:0]    toplevel_execute_ctrl3_down_MMU_L1_ENTRIES_lane0_0_physicalAddress;
  wire                toplevel_execute_ctrl3_down_MMU_L1_ENTRIES_lane0_0_allowRead;
  wire                toplevel_execute_ctrl3_down_MMU_L1_ENTRIES_lane0_0_allowWrite;
  wire                toplevel_execute_ctrl3_down_MMU_L1_ENTRIES_lane0_0_allowExecute;
  wire                toplevel_execute_ctrl3_down_MMU_L1_ENTRIES_lane0_0_allowUser;
  reg        [1:0]    toplevel_execute_ctrl3_down_MMU_L0_HITS_lane0;
  reg        [1:0]    toplevel_execute_ctrl3_down_MMU_L0_HITS_PRE_VALID_lane0;
  wire                toplevel_execute_ctrl3_down_MMU_L0_ENTRIES_lane0_0_valid;
  wire       [13:0]   toplevel_execute_ctrl3_down_MMU_L0_ENTRIES_lane0_0_virtualAddress;
  wire       [19:0]   toplevel_execute_ctrl3_down_MMU_L0_ENTRIES_lane0_0_physicalAddress;
  wire                toplevel_execute_ctrl3_down_MMU_L0_ENTRIES_lane0_0_allowRead;
  wire                toplevel_execute_ctrl3_down_MMU_L0_ENTRIES_lane0_0_allowWrite;
  wire                toplevel_execute_ctrl3_down_MMU_L0_ENTRIES_lane0_0_allowExecute;
  wire                toplevel_execute_ctrl3_down_MMU_L0_ENTRIES_lane0_0_allowUser;
  wire                toplevel_execute_ctrl3_down_MMU_L0_ENTRIES_lane0_1_valid;
  wire       [13:0]   toplevel_execute_ctrl3_down_MMU_L0_ENTRIES_lane0_1_virtualAddress;
  wire       [19:0]   toplevel_execute_ctrl3_down_MMU_L0_ENTRIES_lane0_1_physicalAddress;
  wire                toplevel_execute_ctrl3_down_MMU_L0_ENTRIES_lane0_1_allowRead;
  wire                toplevel_execute_ctrl3_down_MMU_L0_ENTRIES_lane0_1_allowWrite;
  wire                toplevel_execute_ctrl3_down_MMU_L0_ENTRIES_lane0_1_allowExecute;
  wire                toplevel_execute_ctrl3_down_MMU_L0_ENTRIES_lane0_1_allowUser;
  wire       [0:0]    toplevel_execute_ctrl4_down_Decode_INSTRUCTION_SLICE_COUNT_lane1;
  wire       [0:0]    toplevel_execute_ctrl4_down_Decode_INSTRUCTION_SLICE_COUNT_lane0;
  wire                toplevel_execute_ctrl4_down_TRAP_lane1;
  wire                toplevel_execute_ctrl5_down_COMMIT_lane1;
  wire                toplevel_execute_ctrl5_down_LANE_SEL_lane1;
  wire                toplevel_execute_ctrl5_down_COMMIT_lane0;
  wire                toplevel_execute_ctrl5_down_isReady;
  wire                toplevel_execute_ctrl5_down_LANE_SEL_lane0;
  wire                toplevel_execute_ctrl4_down_AguPlugin_FLOAT_lane0;
  wire                toplevel_execute_ctrl4_down_LsuPlugin_logic_FROM_ACCESS_lane0;
  wire                toplevel_execute_ctrl4_down_LsuPlugin_logic_MMU_FAILURE_lane0;
  reg                 toplevel_execute_ctrl4_up_COMMIT_lane0;
  reg                 toplevel_execute_ctrl4_COMMIT_lane0_bypass;
  reg                 toplevel_execute_ctrl4_up_TRAP_lane0;
  wire                toplevel_execute_ctrl4_down_TRAP_lane0;
  reg                 toplevel_execute_ctrl4_TRAP_lane0_bypass;
  wire                toplevel_execute_ctrl4_down_AguPlugin_SEL_lane0;
  wire                toplevel_execute_ctrl4_down_LsuPlugin_logic_FROM_PREFETCH_lane0;
  wire                toplevel_execute_ctrl4_down_LsuPlugin_logic_FENCE_lane0;
  wire                toplevel_execute_ctrl4_down_LsuPlugin_logic_onTrigger_HIT_lane0;
  wire                toplevel_execute_ctrl4_down_LsuPlugin_logic_preCtrl_MISS_ALIGNED_lane0;
  wire                toplevel_execute_ctrl4_down_MMU_BYPASS_TRANSLATION_lane0;
  wire                toplevel_execute_ctrl4_down_LsuPlugin_logic_onPma_FROM_LSU_MSB_FAILED_lane0;
  wire                toplevel_execute_ctrl4_down_MMU_HAZARD_lane0;
  wire                toplevel_execute_ctrl4_down_MMU_REFILL_lane0;
  wire                toplevel_execute_ctrl4_down_MMU_ACCESS_FAULT_lane0;
  wire                toplevel_execute_ctrl4_down_LsuPlugin_logic_MMU_PAGE_FAULT_lane0;
  wire                toplevel_execute_ctrl4_down_LsuPlugin_logic_onPma_IO_RSP_lane0_fault;
  wire                toplevel_execute_ctrl4_down_LsuPlugin_logic_onPma_IO_RSP_lane0_io;
  wire                toplevel_execute_ctrl4_down_AguPlugin_STORE_lane0;
  wire                toplevel_execute_ctrl4_down_LsuPlugin_logic_onPma_CACHED_RSP_lane0_fault;
  wire                toplevel_execute_ctrl4_down_LsuPlugin_logic_onPma_CACHED_RSP_lane0_io;
  wire                toplevel_execute_ctrl4_down_LsuPlugin_logic_preCtrl_IS_AMO_lane0;
  wire       [31:0]   toplevel_execute_ctrl4_down_integer_RS2_lane0;
  wire                toplevel_execute_ctrl4_down_LsuPlugin_logic_onCtrl_SC_MISS_lane0;
  wire       [31:0]   toplevel_execute_ctrl4_down_LsuPlugin_logic_onCtrl_loadData_RESULT_lane0;
  wire       [1:0]    toplevel_execute_ctrl4_down_LsuL1_SIZE_lane0;
  wire                toplevel_execute_ctrl4_down_LsuPlugin_logic_onPma_IO_lane0;
  reg        [31:0]   toplevel_execute_ctrl4_up_integer_RS2_lane0;
  reg                 toplevel_execute_ctrl3_down_MMU_HAZARD_lane0;
  reg                 toplevel_execute_ctrl3_down_MMU_REFILL_lane0;
  reg                 toplevel_execute_ctrl3_down_MMU_ACCESS_FAULT_lane0;
  wire                toplevel_execute_ctrl3_down_LsuPlugin_logic_MMU_FAILURE_lane0;
  reg                 toplevel_execute_ctrl3_down_MMU_ALLOW_READ_lane0;
  reg                 toplevel_execute_ctrl3_down_MMU_ALLOW_WRITE_lane0;
  wire                toplevel_execute_ctrl3_down_AguPlugin_STORE_lane0;
  reg                 toplevel_execute_ctrl3_down_MMU_PAGE_FAULT_lane0;
  wire                toplevel_execute_ctrl3_down_LsuPlugin_logic_MMU_PAGE_FAULT_lane0;
  wire                toplevel_execute_ctrl3_down_LsuPlugin_logic_onPma_FROM_LSU_MSB_FAILED_lane0;
  wire       [31:0]   toplevel_execute_ctrl3_down_early0_SrcPlugin_ADD_SUB_lane0;
  wire                toplevel_execute_ctrl3_down_LsuPlugin_logic_onPma_IO_lane0;
  wire                toplevel_execute_ctrl3_down_LsuPlugin_logic_FROM_PREFETCH_lane0;
  wire                toplevel_execute_ctrl3_down_LsuPlugin_logic_FENCE_lane0;
  wire                toplevel_execute_ctrl3_down_LsuPlugin_logic_onPma_IO_RSP_lane0_fault;
  wire                toplevel_execute_ctrl3_down_LsuPlugin_logic_onPma_IO_RSP_lane0_io;
  wire                toplevel_execute_ctrl3_down_LsuPlugin_logic_onPma_CACHED_RSP_lane0_fault;
  wire                toplevel_execute_ctrl3_down_LsuPlugin_logic_onPma_CACHED_RSP_lane0_io;
  wire                toplevel_execute_ctrl3_down_LsuPlugin_logic_preCtrl_IS_AMO_lane0;
  wire                toplevel_execute_ctrl3_down_LsuL1_ATOMIC_lane0;
  wire                toplevel_execute_ctrl3_down_AguPlugin_SEL_lane0;
  wire                toplevel_execute_ctrl3_down_LsuPlugin_logic_preCtrl_MISS_ALIGNED_lane0;
  reg                 toplevel_execute_ctrl4_LsuL1_SEL_lane0_bypass;
  wire                toplevel_execute_ctrl4_down_LsuPlugin_logic_FROM_LSU_lane0;
  reg                 toplevel_execute_ctrl4_up_LsuL1_SEL_lane0;
  reg                 toplevel_execute_ctrl3_LsuL1_SEL_lane0_bypass;
  wire                toplevel_execute_ctrl3_down_LsuPlugin_logic_FROM_LSU_lane0;
  reg                 toplevel_execute_ctrl3_up_LsuL1_SEL_lane0;
  reg        [31:0]   toplevel_execute_ctrl3_down_MMU_TRANSLATED_lane0;
  wire                toplevel_execute_ctrl2_down_LsuPlugin_logic_FROM_PREFETCH_lane0;
  wire                toplevel_execute_ctrl2_down_LsuPlugin_logic_FROM_LSU_lane0;
  wire       [11:0]   toplevel_execute_ctrl2_down_Decode_STORE_ID_lane0;
  wire                toplevel_execute_ctrl2_down_LsuL1_FLUSH_lane0;
  wire                toplevel_execute_ctrl2_down_LsuL1_PREFETCH_lane0;
  wire                toplevel_execute_ctrl2_down_LsuL1_STORE_lane0;
  wire                toplevel_execute_ctrl2_down_LsuL1_ATOMIC_lane0;
  wire                toplevel_execute_ctrl2_down_LsuL1_LOAD_lane0;
  wire       [1:0]    toplevel_execute_ctrl2_down_LsuL1_SIZE_lane0;
  wire       [3:0]    toplevel_execute_ctrl2_down_LsuL1_MASK_lane0;
  wire                toplevel_execute_ctrl2_down_LsuL1_SEL_lane0;
  wire                toplevel_execute_ctrl2_down_AguPlugin_ATOMIC_lane0;
  wire                toplevel_execute_ctrl2_down_AguPlugin_STORE_lane0;
  wire                toplevel_execute_ctrl2_down_AguPlugin_LOAD_lane0;
  wire       [1:0]    toplevel_execute_ctrl2_down_AguPlugin_SIZE_lane0;
  wire                toplevel_execute_ctrl2_down_AguPlugin_SEL_lane0;
  wire                toplevel_execute_ctrl2_down_LsuPlugin_logic_FROM_WB_lane0;
  wire                toplevel_execute_ctrl2_down_LsuPlugin_logic_FROM_ACCESS_lane0;
  wire                toplevel_execute_ctrl2_down_LsuPlugin_logic_FORCE_PHYSICAL_lane0;
  wire                toplevel_execute_ctrl3_down_LsuPlugin_logic_onTrigger_HIT_lane0;
  wire       [1:0]    toplevel_execute_ctrl3_down_LsuL1_SIZE_lane0;
  wire                toplevel_execute_ctrl3_down_LsuL1_STORE_lane0;
  wire                toplevel_execute_ctrl3_down_LsuL1_LOAD_lane0;
  wire       [31:0]   toplevel_execute_ctrl4_down_LsuL1_READ_DATA_lane0;
  wire       [31:0]   toplevel_execute_ctrl3_down_LsuL1Plugin_logic_EVENT_WRITE_DATA_lane0;
  wire       [3:0]    toplevel_execute_ctrl3_down_LsuL1Plugin_logic_EVENT_WRITE_MASK_lane0;
  wire       [31:0]   toplevel_execute_ctrl4_down_LsuL1Plugin_logic_EVENT_WRITE_DATA_lane0;
  wire       [3:0]    toplevel_execute_ctrl4_down_LsuL1Plugin_logic_EVENT_WRITE_MASK_lane0;
  wire       [1:0]    toplevel_execute_ctrl4_down_LsuL1Plugin_logic_WRITE_TO_READ_HAZARDS_lane0;
  reg        [31:0]   toplevel_execute_ctrl4_down_LsuL1Plugin_logic_BYPASSED_DATA_lane0;
  wire       [3:0]    toplevel_execute_ctrl2_down_LsuL1Plugin_logic_EVENT_WRITE_MASK_lane0;
  wire       [31:0]   toplevel_execute_ctrl2_down_LsuL1Plugin_logic_EVENT_WRITE_DATA_lane0;
  wire                toplevel_execute_ctrl4_down_LsuL1_FLUSH_HIT_lane0;
  wire       [3:0]    toplevel_execute_ctrl4_down_LsuL1_MASK_lane0;
  wire       [31:0]   toplevel_execute_ctrl4_down_LsuL1_WRITE_DATA_lane0;
  wire       [31:0]   toplevel_execute_ctrl4_down_LsuL1_MIXED_ADDRESS_lane0;
  wire                toplevel_execute_ctrl4_down_LsuL1_ABORD_lane0;
  wire       [0:0]    toplevel_execute_ctrl4_down_LsuL1_WAIT_WRITEBACK_lane0;
  wire       [0:0]    toplevel_execute_ctrl4_down_LsuL1_WAIT_REFILL_lane0;
  wire                toplevel_execute_ctrl4_down_LsuL1_SKIP_WRITE_lane0;
  wire                toplevel_execute_ctrl4_down_LsuL1_REFILL_HIT_lane0;
  wire                toplevel_execute_ctrl4_down_LsuL1_MISS_UNIQUE_lane0;
  wire                toplevel_execute_ctrl4_down_LsuL1_FAULT_lane0;
  wire                toplevel_execute_ctrl4_down_LsuL1_MISS_lane0;
  wire                toplevel_execute_ctrl4_down_LsuL1_FLUSH_HAZARD_lane0;
  wire                toplevel_execute_ctrl4_down_LsuL1_HAZARD_lane0;
  wire                toplevel_execute_ctrl4_down_LsuL1Plugin_logic_HAZARD_FORCED_lane0;
  wire                toplevel_execute_ctrl4_down_LsuL1_PREFETCH_lane0;
  wire                toplevel_execute_ctrl4_down_LsuL1_LOAD_lane0;
  wire       [1:0]    toplevel_execute_ctrl4_down_LsuL1Plugin_logic_BANK_BUSY_REMAPPED_lane0;
  wire       [31:0]   toplevel_execute_ctrl4_down_LsuL1_PHYSICAL_ADDRESS_lane0;
  wire                toplevel_execute_ctrl4_down_LsuL1Plugin_logic_WAYS_TAGS_lane0_0_loaded;
  wire       [19:0]   toplevel_execute_ctrl4_down_LsuL1Plugin_logic_WAYS_TAGS_lane0_0_address;
  wire                toplevel_execute_ctrl4_down_LsuL1Plugin_logic_WAYS_TAGS_lane0_0_fault;
  wire                toplevel_execute_ctrl4_down_LsuL1Plugin_logic_WAYS_TAGS_lane0_1_loaded;
  wire       [19:0]   toplevel_execute_ctrl4_down_LsuL1Plugin_logic_WAYS_TAGS_lane0_1_address;
  wire                toplevel_execute_ctrl4_down_LsuL1Plugin_logic_WAYS_TAGS_lane0_1_fault;
  wire       [0:0]    toplevel_execute_ctrl4_down_LsuL1Plugin_logic_SHARED_lane0_plru_0;
  wire       [1:0]    toplevel_execute_ctrl4_down_LsuL1Plugin_logic_SHARED_lane0_dirty;
  wire                toplevel_execute_ctrl4_down_LsuL1_ATOMIC_lane0;
  wire                toplevel_execute_ctrl4_down_LsuL1_STORE_lane0;
  wire                toplevel_execute_ctrl4_down_LsuL1Plugin_logic_NEED_UNIQUE_lane0;
  wire                toplevel_execute_ctrl4_down_LsuL1Plugin_logic_WAYS_HIT_lane0;
  reg        [1:0]    toplevel_execute_ctrl3_down_LsuL1Plugin_logic_WAYS_HITS_lane0;
  wire       [0:0]    toplevel_execute_ctrl3_down_LsuL1Plugin_logic_SHARED_lane0_plru_0;
  wire       [1:0]    toplevel_execute_ctrl3_down_LsuL1Plugin_logic_SHARED_lane0_dirty;
  wire       [0:0]    toplevel_execute_ctrl3_LsuL1Plugin_logic_SHARED_lane0_bypass_plru_0;
  wire       [1:0]    toplevel_execute_ctrl3_LsuL1Plugin_logic_SHARED_lane0_bypass_dirty;
  wire       [0:0]    toplevel_execute_ctrl3_down_LsuL1Plugin_logic_ls_rt0_SHARED_BYPASS_VALUE_lane0_plru_0;
  wire       [1:0]    toplevel_execute_ctrl3_down_LsuL1Plugin_logic_ls_rt0_SHARED_BYPASS_VALUE_lane0_dirty;
  wire                toplevel_execute_ctrl3_down_LsuL1Plugin_logic_ls_rt0_SHARED_BYPASS_VALID_lane0;
  wire                toplevel_execute_ctrl3_down_LsuL1Plugin_logic_WAYS_TAGS_lane0_0_loaded;
  wire       [19:0]   toplevel_execute_ctrl3_down_LsuL1Plugin_logic_WAYS_TAGS_lane0_0_address;
  wire                toplevel_execute_ctrl3_down_LsuL1Plugin_logic_WAYS_TAGS_lane0_0_fault;
  wire                toplevel_execute_ctrl3_down_LsuL1Plugin_logic_WAYS_TAGS_lane0_1_loaded;
  wire       [19:0]   toplevel_execute_ctrl3_down_LsuL1Plugin_logic_WAYS_TAGS_lane0_1_address;
  wire                toplevel_execute_ctrl3_down_LsuL1Plugin_logic_WAYS_TAGS_lane0_1_fault;
  reg        [0:0]    toplevel_execute_ctrl3_up_LsuL1Plugin_logic_SHARED_lane0_plru_0;
  reg        [1:0]    toplevel_execute_ctrl3_up_LsuL1Plugin_logic_SHARED_lane0_dirty;
  wire       [0:0]    toplevel_execute_ctrl2_down_LsuL1Plugin_logic_ls_rt0_SHARED_BYPASS_VALUE_lane0_plru_0;
  wire       [1:0]    toplevel_execute_ctrl2_down_LsuL1Plugin_logic_ls_rt0_SHARED_BYPASS_VALUE_lane0_dirty;
  wire                toplevel_execute_ctrl2_down_LsuL1Plugin_logic_ls_rt0_SHARED_BYPASS_VALID_lane0;
  wire       [31:0]   toplevel_execute_ctrl3_down_LsuL1Plugin_logic_EVENT_WRITE_ADDRESS_lane0;
  wire                toplevel_execute_ctrl3_down_LsuL1Plugin_logic_EVENT_WRITE_VALID_lane0;
  wire       [31:0]   toplevel_execute_ctrl3_down_LsuL1_PHYSICAL_ADDRESS_lane0;
  wire       [31:0]   toplevel_execute_ctrl2_down_LsuL1Plugin_logic_EVENT_WRITE_ADDRESS_lane0;
  wire                toplevel_execute_ctrl2_down_LsuL1Plugin_logic_EVENT_WRITE_VALID_lane0;
  reg        [1:0]    toplevel_execute_ctrl3_down_LsuL1Plugin_logic_WRITE_TO_READ_HAZARDS_lane0;
  wire       [31:0]   toplevel_execute_ctrl4_down_LsuL1Plugin_logic_BANKS_MUXES_lane0_0;
  wire       [31:0]   toplevel_execute_ctrl4_down_LsuL1Plugin_logic_BANKS_MUXES_lane0_1;
  wire       [1:0]    toplevel_execute_ctrl4_down_LsuL1Plugin_logic_WAYS_HITS_lane0;
  wire       [31:0]   toplevel_execute_ctrl4_down_LsuL1Plugin_logic_MUXED_DATA_lane0;
  wire       [31:0]   toplevel_execute_ctrl3_down_LsuL1_MIXED_ADDRESS_lane0;
  wire       [31:0]   toplevel_execute_ctrl3_down_LsuL1Plugin_logic_BANKS_MUXES_lane0_0;
  wire       [31:0]   toplevel_execute_ctrl3_down_LsuL1Plugin_logic_BANKS_MUXES_lane0_1;
  wire       [1:0]    toplevel_execute_ctrl3_down_LsuL1Plugin_logic_BANK_BUSY_lane0;
  reg        [1:0]    toplevel_execute_ctrl3_down_LsuL1Plugin_logic_BANK_BUSY_REMAPPED_lane0;
  wire       [63:0]   toplevel_execute_ctrl3_down_LsuL1Plugin_logic_BANKS_WORDS_lane0_0;
  wire       [63:0]   toplevel_execute_ctrl3_down_LsuL1Plugin_logic_BANKS_WORDS_lane0_1;
  reg        [1:0]    toplevel_execute_ctrl2_down_LsuL1Plugin_logic_BANK_BUSY_lane0;
  wire       [31:0]   toplevel_execute_ctrl2_down_LsuL1_MIXED_ADDRESS_lane0;
  reg                 _zz_3;
  reg                 _zz_4;
  wire       [4:0]    toplevel_execute_ctrl0_down_RS1_PHYS_lane1;
  wire                toplevel_decode_ctrls_0_down_TRAP_1;
  wire                toplevel_decode_ctrls_0_down_TRAP_0;
  wire                toplevel_decode_ctrls_1_down_LANE_SEL_1;
  reg                 toplevel_decode_ctrls_1_LANE_SEL_1_bypass;
  wire                toplevel_decode_ctrls_1_down_LANE_SEL_0;
  reg                 toplevel_decode_ctrls_1_LANE_SEL_0_bypass;
  wire                toplevel_decode_ctrls_0_down_LANE_SEL_1;
  reg                 toplevel_decode_ctrls_0_LANE_SEL_1_bypass;
  wire                toplevel_decode_ctrls_0_down_LANE_SEL_0;
  reg                 toplevel_decode_ctrls_0_LANE_SEL_0_bypass;
  wire       [0:0]    toplevel_execute_ctrl0_up_execute_lane1_LAYER_SEL_lane1;
  wire                toplevel_execute_ctrl0_up_COMPLETED_lane1;
  wire       [0:0]    toplevel_execute_ctrl0_up_LANE_AGE_lane1;
  wire                toplevel_execute_ctrl0_up_DispatchPlugin_logic_hcs_3_onRs_1_ENABLES_0_lane1;
  wire                toplevel_execute_ctrl0_up_DispatchPlugin_logic_hcs_3_onRs_0_ENABLES_0_lane1;
  wire                toplevel_execute_ctrl0_up_DispatchPlugin_logic_hcs_2_onRs_1_ENABLES_0_lane1;
  wire                toplevel_execute_ctrl0_up_DispatchPlugin_logic_hcs_2_onRs_0_ENABLES_0_lane1;
  wire                toplevel_execute_ctrl0_up_DispatchPlugin_logic_hcs_1_onRs_1_ENABLES_1_lane1;
  wire                toplevel_execute_ctrl0_up_DispatchPlugin_logic_hcs_1_onRs_1_ENABLES_0_lane1;
  wire                toplevel_execute_ctrl0_up_DispatchPlugin_logic_hcs_1_onRs_0_ENABLES_0_lane1;
  wire                toplevel_execute_ctrl0_up_DispatchPlugin_logic_hcs_0_onRs_1_ENABLES_0_lane1;
  wire                toplevel_execute_ctrl0_up_DispatchPlugin_logic_hcs_0_onRs_0_ENABLES_0_lane1;
  wire       [4:0]    toplevel_execute_ctrl0_up_RD_PHYS_lane1;
  reg                 toplevel_execute_ctrl0_up_RD_ENABLE_lane1;
  wire       [4:0]    toplevel_execute_ctrl0_up_RS2_PHYS_lane1;
  wire                toplevel_execute_ctrl0_up_RS2_ENABLE_lane1;
  wire       [4:0]    toplevel_execute_ctrl0_up_RS1_PHYS_lane1;
  wire                toplevel_execute_ctrl0_up_RS1_ENABLE_lane1;
  wire       [15:0]   toplevel_execute_ctrl0_up_Decode_UOP_ID_lane1;
  wire                toplevel_execute_ctrl0_up_TRAP_lane1;
  wire       [31:0]   toplevel_execute_ctrl0_up_PC_lane1;
  wire                toplevel_execute_ctrl0_up_DONT_FLUSH_PRECISE_4_lane1;
  wire                toplevel_execute_ctrl0_up_DONT_FLUSH_PRECISE_3_lane1;
  wire       [0:0]    toplevel_execute_ctrl0_up_Decode_INSTRUCTION_SLICE_COUNT_lane1;
  wire                toplevel_execute_ctrl0_up_DispatchPlugin_DONT_FLUSH_FROM_LANES_lane1;
  wire                toplevel_execute_ctrl0_up_DispatchPlugin_DONT_FLUSH_lane1;
  reg                 toplevel_execute_ctrl0_up_DispatchPlugin_MAY_FLUSH_lane1;
  wire                toplevel_execute_ctrl0_up_DispatchPlugin_FENCE_OLDER_lane1;
  wire       [11:0]   toplevel_execute_ctrl0_up_Prediction_BRANCH_HISTORY_lane1;
  wire       [1:0]    toplevel_execute_ctrl0_up_GSharePlugin_GSHARE_COUNTER_lane1_0;
  wire       [1:0]    toplevel_execute_ctrl0_up_GSharePlugin_GSHARE_COUNTER_lane1_1;
  wire       [1:0]    toplevel_execute_ctrl0_up_GSharePlugin_GSHARE_COUNTER_lane1_2;
  wire       [1:0]    toplevel_execute_ctrl0_up_GSharePlugin_GSHARE_COUNTER_lane1_3;
  wire       [3:0]    toplevel_execute_ctrl0_up_Prediction_ALIGNED_SLICES_BRANCH_lane1;
  wire       [3:0]    toplevel_execute_ctrl0_up_Prediction_ALIGNED_SLICES_TAKEN_lane1;
  wire       [31:0]   toplevel_execute_ctrl0_up_Prediction_ALIGNED_JUMPED_PC_lane1;
  wire                toplevel_execute_ctrl0_up_Prediction_ALIGNED_JUMPED_lane1;
  wire       [31:0]   toplevel_execute_ctrl0_up_Decode_UOP_lane1;
  wire                toplevel_execute_ctrl0_up_LANE_SEL_lane1;
  wire       [0:0]    toplevel_execute_ctrl0_up_execute_lane0_LAYER_SEL_lane0;
  wire                toplevel_execute_ctrl0_up_COMPLETED_lane0;
  wire       [0:0]    toplevel_execute_ctrl0_up_LANE_AGE_lane0;
  wire                toplevel_execute_ctrl0_up_DispatchPlugin_logic_hcs_3_onRs_1_ENABLES_0_lane0;
  wire                toplevel_execute_ctrl0_up_DispatchPlugin_logic_hcs_3_onRs_0_ENABLES_0_lane0;
  wire                toplevel_execute_ctrl0_up_DispatchPlugin_logic_hcs_2_onRs_1_ENABLES_0_lane0;
  wire                toplevel_execute_ctrl0_up_DispatchPlugin_logic_hcs_2_onRs_0_ENABLES_0_lane0;
  wire                toplevel_execute_ctrl0_up_DispatchPlugin_logic_hcs_1_onRs_1_ENABLES_1_lane0;
  wire                toplevel_execute_ctrl0_up_DispatchPlugin_logic_hcs_1_onRs_1_ENABLES_0_lane0;
  wire                toplevel_execute_ctrl0_up_DispatchPlugin_logic_hcs_1_onRs_0_ENABLES_0_lane0;
  wire                toplevel_execute_ctrl0_up_DispatchPlugin_logic_hcs_0_onRs_1_ENABLES_0_lane0;
  wire                toplevel_execute_ctrl0_up_DispatchPlugin_logic_hcs_0_onRs_0_ENABLES_0_lane0;
  wire       [4:0]    toplevel_execute_ctrl0_up_RD_PHYS_lane0;
  reg                 toplevel_execute_ctrl0_up_RD_ENABLE_lane0;
  wire       [4:0]    toplevel_execute_ctrl0_up_RS2_PHYS_lane0;
  wire                toplevel_execute_ctrl0_up_RS2_ENABLE_lane0;
  wire       [4:0]    toplevel_execute_ctrl0_up_RS1_PHYS_lane0;
  wire                toplevel_execute_ctrl0_up_RS1_ENABLE_lane0;
  wire       [15:0]   toplevel_execute_ctrl0_up_Decode_UOP_ID_lane0;
  wire                toplevel_execute_ctrl0_up_TRAP_lane0;
  wire       [31:0]   toplevel_execute_ctrl0_up_PC_lane0;
  wire                toplevel_execute_ctrl0_up_DONT_FLUSH_PRECISE_4_lane0;
  wire                toplevel_execute_ctrl0_up_DONT_FLUSH_PRECISE_3_lane0;
  wire       [0:0]    toplevel_execute_ctrl0_up_Decode_INSTRUCTION_SLICE_COUNT_lane0;
  wire                toplevel_execute_ctrl0_up_DispatchPlugin_DONT_FLUSH_FROM_LANES_lane0;
  wire                toplevel_execute_ctrl0_up_DispatchPlugin_DONT_FLUSH_lane0;
  reg                 toplevel_execute_ctrl0_up_DispatchPlugin_MAY_FLUSH_lane0;
  wire                toplevel_execute_ctrl0_up_DispatchPlugin_FENCE_OLDER_lane0;
  wire       [11:0]   toplevel_execute_ctrl0_up_Prediction_BRANCH_HISTORY_lane0;
  wire       [1:0]    toplevel_execute_ctrl0_up_GSharePlugin_GSHARE_COUNTER_lane0_0;
  wire       [1:0]    toplevel_execute_ctrl0_up_GSharePlugin_GSHARE_COUNTER_lane0_1;
  wire       [1:0]    toplevel_execute_ctrl0_up_GSharePlugin_GSHARE_COUNTER_lane0_2;
  wire       [1:0]    toplevel_execute_ctrl0_up_GSharePlugin_GSHARE_COUNTER_lane0_3;
  wire       [3:0]    toplevel_execute_ctrl0_up_Prediction_ALIGNED_SLICES_BRANCH_lane0;
  wire       [3:0]    toplevel_execute_ctrl0_up_Prediction_ALIGNED_SLICES_TAKEN_lane0;
  wire       [31:0]   toplevel_execute_ctrl0_up_Prediction_ALIGNED_JUMPED_PC_lane0;
  wire                toplevel_execute_ctrl0_up_Prediction_ALIGNED_JUMPED_lane0;
  wire       [31:0]   toplevel_execute_ctrl0_up_Decode_UOP_lane0;
  wire                toplevel_execute_ctrl0_up_LANE_SEL_lane0;
  wire                toplevel_decode_ctrls_0_up_isMoving;
  wire                fetch_logic_ctrls_2_down_BtbPlugin_logic_chunksLogic_1_hitCalc_HIT;
  wire                fetch_logic_ctrls_2_down_BtbPlugin_logic_chunksLogic_0_hitCalc_HIT;
  wire                fetch_logic_ctrls_1_down_isReady;
  wire                fetch_logic_ctrls_2_down_BtbPlugin_logic_chunksLogic_1_predict_TAKEN;
  wire       [15:0]   fetch_logic_ctrls_2_down_BtbPlugin_logic_chunksLogic_1_readRsp_ENTRY_hash;
  wire       [0:0]    fetch_logic_ctrls_2_down_BtbPlugin_logic_chunksLogic_1_readRsp_ENTRY_sliceLow;
  wire       [30:0]   fetch_logic_ctrls_2_down_BtbPlugin_logic_chunksLogic_1_readRsp_ENTRY_pcTarget;
  wire                fetch_logic_ctrls_2_down_BtbPlugin_logic_chunksLogic_1_readRsp_ENTRY_isBranch;
  wire                fetch_logic_ctrls_2_down_BtbPlugin_logic_chunksLogic_1_readRsp_ENTRY_isPush;
  wire                fetch_logic_ctrls_2_down_BtbPlugin_logic_chunksLogic_1_readRsp_ENTRY_isPop;
  wire                fetch_logic_ctrls_1_down_BtbPlugin_logic_chunksLogic_1_hitCalc_HIT;
  (* keep , syn_keep *) wire       [15:0]   fetch_logic_ctrls_1_down_BtbPlugin_logic_chunksLogic_1_readRsp_ENTRY_hash /* synthesis syn_keep = 1 */ ;
  (* keep , syn_keep *) wire       [0:0]    fetch_logic_ctrls_1_down_BtbPlugin_logic_chunksLogic_1_readRsp_ENTRY_sliceLow /* synthesis syn_keep = 1 */ ;
  (* keep , syn_keep *) wire       [30:0]   fetch_logic_ctrls_1_down_BtbPlugin_logic_chunksLogic_1_readRsp_ENTRY_pcTarget /* synthesis syn_keep = 1 */ ;
  (* keep , syn_keep *) wire                fetch_logic_ctrls_1_down_BtbPlugin_logic_chunksLogic_1_readRsp_ENTRY_isBranch /* synthesis syn_keep = 1 */ ;
  (* keep , syn_keep *) wire                fetch_logic_ctrls_1_down_BtbPlugin_logic_chunksLogic_1_readRsp_ENTRY_isPush /* synthesis syn_keep = 1 */ ;
  (* keep , syn_keep *) wire                fetch_logic_ctrls_1_down_BtbPlugin_logic_chunksLogic_1_readRsp_ENTRY_isPop /* synthesis syn_keep = 1 */ ;
  wire                fetch_logic_ctrls_2_down_BtbPlugin_logic_chunksLogic_0_predict_TAKEN;
  wire       [15:0]   fetch_logic_ctrls_2_down_BtbPlugin_logic_chunksLogic_0_readRsp_ENTRY_hash;
  wire       [0:0]    fetch_logic_ctrls_2_down_BtbPlugin_logic_chunksLogic_0_readRsp_ENTRY_sliceLow;
  wire       [30:0]   fetch_logic_ctrls_2_down_BtbPlugin_logic_chunksLogic_0_readRsp_ENTRY_pcTarget;
  wire                fetch_logic_ctrls_2_down_BtbPlugin_logic_chunksLogic_0_readRsp_ENTRY_isBranch;
  wire                fetch_logic_ctrls_2_down_BtbPlugin_logic_chunksLogic_0_readRsp_ENTRY_isPush;
  wire                fetch_logic_ctrls_2_down_BtbPlugin_logic_chunksLogic_0_readRsp_ENTRY_isPop;
  wire       [1:0]    fetch_logic_ctrls_1_down_BtbPlugin_logic_readCmd_HAZARDS;
  wire                fetch_logic_ctrls_1_up_isValid;
  wire                fetch_logic_ctrls_1_down_BtbPlugin_logic_chunksLogic_0_hitCalc_HIT;
  (* keep , syn_keep *) wire       [15:0]   fetch_logic_ctrls_1_down_BtbPlugin_logic_chunksLogic_0_readRsp_ENTRY_hash /* synthesis syn_keep = 1 */ ;
  (* keep , syn_keep *) wire       [0:0]    fetch_logic_ctrls_1_down_BtbPlugin_logic_chunksLogic_0_readRsp_ENTRY_sliceLow /* synthesis syn_keep = 1 */ ;
  (* keep , syn_keep *) wire       [30:0]   fetch_logic_ctrls_1_down_BtbPlugin_logic_chunksLogic_0_readRsp_ENTRY_pcTarget /* synthesis syn_keep = 1 */ ;
  (* keep , syn_keep *) wire                fetch_logic_ctrls_1_down_BtbPlugin_logic_chunksLogic_0_readRsp_ENTRY_isBranch /* synthesis syn_keep = 1 */ ;
  (* keep , syn_keep *) wire                fetch_logic_ctrls_1_down_BtbPlugin_logic_chunksLogic_0_readRsp_ENTRY_isPush /* synthesis syn_keep = 1 */ ;
  (* keep , syn_keep *) wire                fetch_logic_ctrls_1_down_BtbPlugin_logic_chunksLogic_0_readRsp_ENTRY_isPop /* synthesis syn_keep = 1 */ ;
  wire       [1:0]    fetch_logic_ctrls_0_down_BtbPlugin_logic_readCmd_HAZARDS;
  wire       [15:0]   toplevel_execute_ctrl0_down_Decode_UOP_ID_lane1;
  wire                toplevel_execute_ctrl0_down_LANE_SEL_lane1;
  wire       [15:0]   toplevel_execute_ctrl0_down_Decode_UOP_ID_lane0;
  wire                toplevel_execute_ctrl0_down_isReady;
  wire                toplevel_execute_ctrl0_down_LANE_SEL_lane0;
  wire       [9:0]    toplevel_decode_ctrls_1_down_Decode_DOP_ID_1;
  wire       [9:0]    toplevel_decode_ctrls_1_down_Decode_DOP_ID_0;
  wire                toplevel_decode_ctrls_1_down_DecoderPlugin_logic_NEED_RM_1;
  wire                toplevel_decode_ctrls_1_down_DecoderPlugin_logic_NEED_FPU_1;
  wire                toplevel_decode_ctrls_1_down_DecoderPlugin_logic_NEED_RM_0;
  wire                toplevel_decode_ctrls_1_down_DecoderPlugin_logic_NEED_FPU_0;
  wire                toplevel_decode_ctrls_1_down_DispatchPlugin_logic_hcs_3_onRs_1_ENABLES_0_1;
  wire                toplevel_decode_ctrls_1_down_DispatchPlugin_logic_hcs_3_onRs_0_ENABLES_0_1;
  wire                toplevel_decode_ctrls_1_down_DispatchPlugin_logic_hcs_2_onRs_1_ENABLES_0_1;
  wire                toplevel_decode_ctrls_1_down_DispatchPlugin_logic_hcs_2_onRs_0_ENABLES_0_1;
  wire                toplevel_decode_ctrls_1_down_DispatchPlugin_logic_hcs_1_onRs_1_ENABLES_1_1;
  wire                toplevel_decode_ctrls_1_down_DispatchPlugin_logic_hcs_1_onRs_1_ENABLES_0_1;
  wire                toplevel_decode_ctrls_1_down_DispatchPlugin_logic_hcs_1_onRs_0_ENABLES_0_1;
  wire                toplevel_decode_ctrls_1_down_DispatchPlugin_logic_hcs_0_onRs_1_ENABLES_0_1;
  wire                toplevel_decode_ctrls_1_down_DispatchPlugin_logic_hcs_0_onRs_0_ENABLES_0_1;
  wire                toplevel_decode_ctrls_1_down_DONT_FLUSH_PRECISE_4_1;
  wire                toplevel_decode_ctrls_1_down_DONT_FLUSH_PRECISE_3_1;
  wire                toplevel_decode_ctrls_1_down_DispatchPlugin_DONT_FLUSH_FROM_LANES_1;
  wire                toplevel_decode_ctrls_1_down_DispatchPlugin_DONT_FLUSH_1;
  wire                toplevel_decode_ctrls_1_down_DispatchPlugin_MAY_FLUSH_1;
  wire                toplevel_decode_ctrls_1_down_DispatchPlugin_FENCE_OLDER_1;
  wire       [11:0]   toplevel_decode_ctrls_1_down_Prediction_BRANCH_HISTORY_1;
  wire       [1:0]    toplevel_decode_ctrls_1_down_GSharePlugin_GSHARE_COUNTER_1_0;
  wire       [1:0]    toplevel_decode_ctrls_1_down_GSharePlugin_GSHARE_COUNTER_1_1;
  wire       [1:0]    toplevel_decode_ctrls_1_down_GSharePlugin_GSHARE_COUNTER_1_2;
  wire       [1:0]    toplevel_decode_ctrls_1_down_GSharePlugin_GSHARE_COUNTER_1_3;
  wire       [3:0]    toplevel_decode_ctrls_1_down_Prediction_ALIGNED_SLICES_BRANCH_1;
  wire       [3:0]    toplevel_decode_ctrls_1_down_Prediction_ALIGNED_SLICES_TAKEN_1;
  wire       [31:0]   toplevel_decode_ctrls_1_down_Prediction_ALIGNED_JUMPED_PC_1;
  wire                toplevel_decode_ctrls_1_down_DispatchPlugin_logic_LANES_LAYER_HIT_3_1;
  wire                toplevel_decode_ctrls_1_down_DispatchPlugin_logic_LANES_LAYER_HIT_2_1;
  wire                toplevel_decode_ctrls_1_down_DispatchPlugin_logic_LANES_LAYER_HIT_1_1;
  wire                toplevel_decode_ctrls_1_down_DispatchPlugin_logic_LANES_LAYER_HIT_0_1;
  wire                toplevel_decode_ctrls_1_down_DispatchPlugin_logic_hcs_3_onRs_1_ENABLES_0_0;
  wire                toplevel_decode_ctrls_1_down_DispatchPlugin_logic_hcs_3_onRs_0_ENABLES_0_0;
  wire                toplevel_decode_ctrls_1_down_DispatchPlugin_logic_hcs_2_onRs_1_ENABLES_0_0;
  wire                toplevel_decode_ctrls_1_down_DispatchPlugin_logic_hcs_2_onRs_0_ENABLES_0_0;
  wire                toplevel_decode_ctrls_1_down_DispatchPlugin_logic_hcs_1_onRs_1_ENABLES_1_0;
  wire                toplevel_decode_ctrls_1_down_DispatchPlugin_logic_hcs_1_onRs_1_ENABLES_0_0;
  wire                toplevel_decode_ctrls_1_down_DispatchPlugin_logic_hcs_1_onRs_0_ENABLES_0_0;
  wire                toplevel_decode_ctrls_1_down_DispatchPlugin_logic_hcs_0_onRs_1_ENABLES_0_0;
  wire                toplevel_decode_ctrls_1_down_DispatchPlugin_logic_hcs_0_onRs_0_ENABLES_0_0;
  wire                toplevel_decode_ctrls_1_down_DONT_FLUSH_PRECISE_4_0;
  wire                toplevel_decode_ctrls_1_down_DONT_FLUSH_PRECISE_3_0;
  wire                toplevel_decode_ctrls_1_down_DispatchPlugin_DONT_FLUSH_FROM_LANES_0;
  wire                toplevel_decode_ctrls_1_down_DispatchPlugin_DONT_FLUSH_0;
  wire                toplevel_decode_ctrls_1_down_DispatchPlugin_MAY_FLUSH_0;
  wire                toplevel_decode_ctrls_1_down_DispatchPlugin_FENCE_OLDER_0;
  wire       [11:0]   toplevel_decode_ctrls_1_down_Prediction_BRANCH_HISTORY_0;
  wire       [1:0]    toplevel_decode_ctrls_1_down_GSharePlugin_GSHARE_COUNTER_0_0;
  wire       [1:0]    toplevel_decode_ctrls_1_down_GSharePlugin_GSHARE_COUNTER_0_1;
  wire       [1:0]    toplevel_decode_ctrls_1_down_GSharePlugin_GSHARE_COUNTER_0_2;
  wire       [1:0]    toplevel_decode_ctrls_1_down_GSharePlugin_GSHARE_COUNTER_0_3;
  wire       [3:0]    toplevel_decode_ctrls_1_down_Prediction_ALIGNED_SLICES_BRANCH_0;
  wire       [3:0]    toplevel_decode_ctrls_1_down_Prediction_ALIGNED_SLICES_TAKEN_0;
  wire       [31:0]   toplevel_decode_ctrls_1_down_Prediction_ALIGNED_JUMPED_PC_0;
  wire                toplevel_decode_ctrls_1_down_DispatchPlugin_logic_LANES_LAYER_HIT_3_0;
  wire                toplevel_decode_ctrls_1_down_DispatchPlugin_logic_LANES_LAYER_HIT_2_0;
  wire                toplevel_decode_ctrls_1_down_DispatchPlugin_logic_LANES_LAYER_HIT_1_0;
  wire                toplevel_decode_ctrls_1_down_DispatchPlugin_logic_LANES_LAYER_HIT_0_0;
  wire                toplevel_decode_ctrls_1_up_isValid;
  reg                 toplevel_decode_ctrls_1_down_ready;
  wire                toplevel_execute_ctrl2_down_MAY_FLUSH_PRECISE_3_lane1;
  wire                toplevel_execute_ctrl1_down_MAY_FLUSH_PRECISE_4_lane1;
  wire                toplevel_execute_ctrl1_down_MAY_FLUSH_PRECISE_3_lane1;
  wire                toplevel_execute_ctrl2_down_MAY_FLUSH_PRECISE_3_lane0;
  wire                toplevel_execute_ctrl1_down_MAY_FLUSH_PRECISE_4_lane0;
  wire                toplevel_execute_ctrl1_down_MAY_FLUSH_PRECISE_3_lane0;
  wire                toplevel_execute_ctrl2_down_BYPASSED_AT_3_lane1;
  reg        [4:0]    toplevel_execute_ctrl2_up_RD_PHYS_lane1;
  wire                toplevel_execute_ctrl1_down_BYPASSED_AT_2_lane1;
  reg        [4:0]    toplevel_execute_ctrl1_up_RD_PHYS_lane1;
  reg                 toplevel_execute_ctrl1_up_RD_ENABLE_lane1;
  wire                toplevel_execute_ctrl2_down_BYPASSED_AT_3_lane0;
  reg        [4:0]    toplevel_execute_ctrl2_up_RD_PHYS_lane0;
  wire                toplevel_execute_ctrl1_down_BYPASSED_AT_2_lane0;
  reg        [4:0]    toplevel_execute_ctrl1_up_RD_PHYS_lane0;
  reg                 toplevel_execute_ctrl1_up_RD_ENABLE_lane0;
  wire       [4:0]    toplevel_execute_ctrl4_down_RD_PHYS_lane1;
  wire                toplevel_execute_ctrl4_down_lane1_integer_WriteBackPlugin_SEL_lane1;
  wire                toplevel_execute_ctrl4_down_COMMIT_lane1;
  reg                 toplevel_execute_ctrl4_up_RD_ENABLE_lane1;
  wire                toplevel_execute_ctrl4_down_LANE_SEL_lane1;
  wire       [31:0]   toplevel_execute_ctrl4_down_lane1_integer_WriteBackPlugin_logic_DATA_lane1;
  wire       [31:0]   toplevel_execute_ctrl4_lane1_integer_WriteBackPlugin_logic_DATA_lane1_bypass;
  reg        [31:0]   toplevel_execute_ctrl4_up_lane1_integer_WriteBackPlugin_logic_DATA_lane1;
  wire                toplevel_execute_ctrl3_down_COMMIT_lane1;
  reg                 toplevel_execute_ctrl3_up_RD_ENABLE_lane1;
  wire                toplevel_execute_ctrl3_down_LANE_SEL_lane1;
  wire       [31:0]   toplevel_execute_ctrl3_down_lane1_integer_WriteBackPlugin_logic_DATA_lane1;
  wire       [31:0]   toplevel_execute_ctrl3_lane1_integer_WriteBackPlugin_logic_DATA_lane1_bypass;
  reg        [31:0]   toplevel_execute_ctrl3_up_lane1_integer_WriteBackPlugin_logic_DATA_lane1;
  wire       [15:0]   toplevel_execute_ctrl2_down_Decode_UOP_ID_lane1;
  wire                toplevel_execute_ctrl2_down_COMMIT_lane1;
  reg                 toplevel_execute_ctrl2_up_RD_ENABLE_lane1;
  wire                toplevel_execute_ctrl2_down_LANE_SEL_lane1;
  wire       [31:0]   toplevel_execute_ctrl2_down_lane1_integer_WriteBackPlugin_logic_DATA_lane1;
  wire       [31:0]   toplevel_execute_ctrl2_lane1_integer_WriteBackPlugin_logic_DATA_lane1_bypass;
  wire       [4:0]    toplevel_execute_ctrl4_down_RD_PHYS_lane0;
  wire                toplevel_execute_ctrl4_down_lane0_integer_WriteBackPlugin_SEL_lane0;
  wire                toplevel_execute_ctrl4_down_COMMIT_lane0;
  reg                 toplevel_execute_ctrl4_up_RD_ENABLE_lane0;
  wire                toplevel_execute_ctrl4_down_LANE_SEL_lane0;
  wire       [31:0]   toplevel_execute_ctrl4_down_lane0_integer_WriteBackPlugin_logic_DATA_lane0;
  wire       [31:0]   toplevel_execute_ctrl4_lane0_integer_WriteBackPlugin_logic_DATA_lane0_bypass;
  reg        [31:0]   toplevel_execute_ctrl4_up_lane0_integer_WriteBackPlugin_logic_DATA_lane0;
  wire                toplevel_execute_ctrl3_down_COMMIT_lane0;
  reg                 toplevel_execute_ctrl3_up_RD_ENABLE_lane0;
  wire                toplevel_execute_ctrl3_down_isReady;
  wire                toplevel_execute_ctrl3_down_LANE_SEL_lane0;
  wire       [31:0]   toplevel_execute_ctrl3_down_lane0_integer_WriteBackPlugin_logic_DATA_lane0;
  wire       [31:0]   toplevel_execute_ctrl3_lane0_integer_WriteBackPlugin_logic_DATA_lane0_bypass;
  reg        [31:0]   toplevel_execute_ctrl3_up_lane0_integer_WriteBackPlugin_logic_DATA_lane0;
  reg                 toplevel_execute_ctrl2_up_RD_ENABLE_lane0;
  wire                toplevel_execute_ctrl2_down_LANE_SEL_lane0;
  wire       [31:0]   toplevel_execute_ctrl2_down_lane0_integer_WriteBackPlugin_logic_DATA_lane0;
  wire       [31:0]   toplevel_execute_ctrl2_lane0_integer_WriteBackPlugin_logic_DATA_lane0_bypass;
  wire       [31:0]   toplevel_decode_ctrls_1_down_Decode_UOP_1;
  reg                 toplevel_decode_ctrls_1_up_TRAP_1;
  reg                 toplevel_decode_ctrls_1_TRAP_1_bypass;
  wire       [15:0]   toplevel_decode_ctrls_1_down_Decode_UOP_ID_1;
  wire                toplevel_decode_ctrls_1_down_TRAP_1;
  wire       [0:0]    toplevel_decode_ctrls_1_down_Decode_INSTRUCTION_SLICE_COUNT_1;
  wire       [31:0]   toplevel_decode_ctrls_1_down_PC_1;
  wire                toplevel_decode_ctrls_1_down_Prediction_ALIGN_REDO_1;
  wire                toplevel_decode_ctrls_1_down_Prediction_ALIGNED_JUMPED_1;
  reg                 toplevel_decode_ctrls_1_up_LANE_SEL_1;
  wire       [31:0]   toplevel_decode_ctrls_1_down_Decode_INSTRUCTION_RAW_1;
  wire                toplevel_decode_ctrls_1_down_Decode_DECOMPRESSION_FAULT_1;
  wire                toplevel_decode_ctrls_1_down_Decode_LEGAL_1;
  wire       [4:0]    toplevel_decode_ctrls_1_down_RD_PHYS_1;
  reg                 toplevel_decode_ctrls_1_down_RD_ENABLE_1;
  wire       [4:0]    toplevel_decode_ctrls_1_down_RS2_PHYS_1;
  wire                toplevel_decode_ctrls_1_down_RS2_ENABLE_1;
  wire       [4:0]    toplevel_decode_ctrls_1_down_RS1_PHYS_1;
  wire       [31:0]   toplevel_decode_ctrls_1_down_Decode_INSTRUCTION_1;
  wire                toplevel_decode_ctrls_1_down_RS1_ENABLE_1;
  wire                toplevel_decode_ctrls_1_lane1_upIsCancel;
  wire                toplevel_decode_ctrls_1_lane1_downIsCancel;
  wire       [31:0]   toplevel_decode_ctrls_1_down_Decode_UOP_0;
  reg                 toplevel_decode_ctrls_1_up_TRAP_0;
  reg                 toplevel_decode_ctrls_1_TRAP_0_bypass;
  wire       [15:0]   toplevel_decode_ctrls_1_down_Decode_UOP_ID_0;
  wire                toplevel_decode_ctrls_1_up_isReady;
  wire                toplevel_decode_ctrls_1_down_TRAP_0;
  wire       [0:0]    toplevel_decode_ctrls_1_down_Decode_INSTRUCTION_SLICE_COUNT_0;
  wire       [31:0]   toplevel_decode_ctrls_1_down_PC_0;
  wire                toplevel_decode_ctrls_1_down_Prediction_ALIGN_REDO_0;
  wire                toplevel_decode_ctrls_1_down_Prediction_ALIGNED_JUMPED_0;
  reg                 toplevel_decode_ctrls_1_up_LANE_SEL_0;
  wire       [31:0]   toplevel_decode_ctrls_1_down_Decode_INSTRUCTION_RAW_0;
  wire                toplevel_decode_ctrls_1_down_Decode_DECOMPRESSION_FAULT_0;
  wire                toplevel_decode_ctrls_1_down_Decode_LEGAL_0;
  wire       [4:0]    toplevel_decode_ctrls_1_down_RD_PHYS_0;
  reg                 toplevel_decode_ctrls_1_down_RD_ENABLE_0;
  wire       [4:0]    toplevel_decode_ctrls_1_down_RS2_PHYS_0;
  wire                toplevel_decode_ctrls_1_down_RS2_ENABLE_0;
  wire       [4:0]    toplevel_decode_ctrls_1_down_RS1_PHYS_0;
  wire       [31:0]   toplevel_decode_ctrls_1_down_Decode_INSTRUCTION_0;
  wire                toplevel_decode_ctrls_1_down_RS1_ENABLE_0;
  wire                toplevel_decode_ctrls_1_up_isCanceling;
  wire                toplevel_decode_ctrls_1_up_ready;
  reg                 toplevel_decode_ctrls_1_up_valid;
  wire                toplevel_decode_ctrls_1_up_isMoving;
  wire                toplevel_execute_ctrl4_down_COMPLETION_AT_4_lane0;
  reg                 toplevel_execute_ctrl4_up_COMPLETED_lane0;
  wire                toplevel_execute_ctrl4_down_COMPLETED_lane0;
  wire                toplevel_execute_ctrl4_COMPLETED_lane0_bypass;
  wire                toplevel_execute_ctrl3_down_COMPLETION_AT_3_lane0;
  reg                 toplevel_execute_ctrl3_up_COMPLETED_lane0;
  wire                toplevel_execute_ctrl3_down_COMPLETED_lane0;
  wire                toplevel_execute_ctrl3_COMPLETED_lane0_bypass;
  wire                toplevel_execute_ctrl2_down_COMPLETION_AT_2_lane0;
  reg                 toplevel_execute_ctrl2_up_COMPLETED_lane0;
  wire                toplevel_execute_ctrl2_down_COMPLETED_lane0;
  wire                toplevel_execute_ctrl2_COMPLETED_lane0_bypass;
  reg                 toplevel_execute_ctrl1_up_LANE_SEL_lane0;
  wire                toplevel_execute_ctrl4_down_COMPLETION_AT_4_lane1;
  reg                 toplevel_execute_ctrl4_up_COMPLETED_lane1;
  wire                toplevel_execute_ctrl4_down_COMPLETED_lane1;
  wire                toplevel_execute_ctrl4_COMPLETED_lane1_bypass;
  wire                toplevel_execute_ctrl3_down_COMPLETION_AT_3_lane1;
  reg                 toplevel_execute_ctrl3_up_COMPLETED_lane1;
  wire                toplevel_execute_ctrl3_down_COMPLETED_lane1;
  wire                toplevel_execute_ctrl3_COMPLETED_lane1_bypass;
  wire                toplevel_execute_ctrl2_down_COMPLETION_AT_2_lane1;
  reg                 toplevel_execute_ctrl2_up_COMPLETED_lane1;
  wire                toplevel_execute_ctrl2_down_COMPLETED_lane1;
  wire                toplevel_execute_ctrl2_COMPLETED_lane1_bypass;
  reg                 toplevel_execute_ctrl1_up_LANE_SEL_lane1;
  wire       [1:0]    toplevel_execute_ctrl4_down_GSharePlugin_GSHARE_COUNTER_lane1_0;
  wire       [1:0]    toplevel_execute_ctrl4_down_GSharePlugin_GSHARE_COUNTER_lane1_1;
  wire       [1:0]    toplevel_execute_ctrl4_down_GSharePlugin_GSHARE_COUNTER_lane1_2;
  wire       [1:0]    toplevel_execute_ctrl4_down_GSharePlugin_GSHARE_COUNTER_lane1_3;
  wire       [31:0]   toplevel_execute_ctrl4_down_early1_BranchPlugin_pcCalc_PC_LAST_SLICE_lane1;
  wire                toplevel_execute_ctrl4_down_early1_BranchPlugin_SEL_lane1;
  wire                toplevel_execute_ctrl4_down_late1_BranchPlugin_logic_jumpLogic_IS_JALR_lane1;
  wire                toplevel_execute_ctrl4_down_late1_BranchPlugin_logic_jumpLogic_IS_JAL_lane1;
  wire                toplevel_execute_ctrl4_down_late1_BranchPlugin_logic_jumpLogic_MISSALIGNED_lane1;
  wire       [15:0]   toplevel_execute_ctrl4_down_Decode_UOP_ID_lane1;
  wire       [0:0]    toplevel_execute_ctrl4_down_LANE_AGE_lane1;
  reg        [11:0]   late1_BranchPlugin_logic_jumpLogic_history_fromFetch_shifter_4;
  reg        [11:0]   late1_BranchPlugin_logic_jumpLogic_history_fromFetch_shifter_3;
  reg        [11:0]   late1_BranchPlugin_logic_jumpLogic_history_fromFetch_shifter_2;
  reg        [11:0]   late1_BranchPlugin_logic_jumpLogic_history_fromFetch_shifter_1;
  wire       [3:0]    toplevel_execute_ctrl4_down_Prediction_ALIGNED_SLICES_TAKEN_lane1;
  wire       [3:0]    toplevel_execute_ctrl4_down_Prediction_ALIGNED_SLICES_BRANCH_lane1;
  wire       [11:0]   toplevel_execute_ctrl4_down_Prediction_BRANCH_HISTORY_lane1;
  wire       [31:0]   toplevel_execute_ctrl4_down_PC_lane1;
  wire                toplevel_execute_ctrl4_down_late1_BranchPlugin_SEL_lane1;
  wire                toplevel_execute_ctrl4_down_Prediction_ALIGNED_JUMPED_lane1;
  wire       [31:0]   toplevel_execute_ctrl4_down_late1_BranchPlugin_logic_jumpLogic_btb_REAL_TARGET_lane1;
  wire       [31:0]   toplevel_execute_ctrl4_down_early1_BranchPlugin_pcCalc_PC_FALSE_lane1;
  wire                toplevel_execute_ctrl4_down_late1_BranchPlugin_logic_jumpLogic_COND_lane1;
  wire       [31:0]   toplevel_execute_ctrl4_down_Decode_UOP_lane1;
  wire                toplevel_execute_ctrl4_down_late1_BranchPlugin_logic_alu_MSB_FAILED_lane1;
  wire       [1:0]    toplevel_execute_ctrl4_down_BranchPlugin_BRANCH_CTRL_lane1;
  wire                toplevel_execute_ctrl4_down_late1_BranchPlugin_logic_alu_btb_BAD_TARGET_lane1;
  wire       [31:0]   toplevel_execute_ctrl4_down_early1_BranchPlugin_pcCalc_PC_TRUE_lane1;
  wire       [31:0]   toplevel_execute_ctrl4_down_Prediction_ALIGNED_JUMPED_PC_lane1;
  wire                toplevel_execute_ctrl4_down_late1_BranchPlugin_logic_alu_EQ_lane1;
  wire       [1:0]    toplevel_execute_ctrl4_down_GSharePlugin_GSHARE_COUNTER_lane0_0;
  wire       [1:0]    toplevel_execute_ctrl4_down_GSharePlugin_GSHARE_COUNTER_lane0_1;
  wire       [1:0]    toplevel_execute_ctrl4_down_GSharePlugin_GSHARE_COUNTER_lane0_2;
  wire       [1:0]    toplevel_execute_ctrl4_down_GSharePlugin_GSHARE_COUNTER_lane0_3;
  wire       [31:0]   toplevel_execute_ctrl4_down_early0_BranchPlugin_pcCalc_PC_LAST_SLICE_lane0;
  wire                toplevel_execute_ctrl4_down_early0_BranchPlugin_SEL_lane0;
  wire                toplevel_execute_ctrl4_down_late0_BranchPlugin_logic_jumpLogic_IS_JALR_lane0;
  wire                toplevel_execute_ctrl4_down_late0_BranchPlugin_logic_jumpLogic_IS_JAL_lane0;
  wire                toplevel_execute_ctrl4_down_late0_BranchPlugin_logic_jumpLogic_MISSALIGNED_lane0;
  wire       [15:0]   toplevel_execute_ctrl4_down_Decode_UOP_ID_lane0;
  wire       [0:0]    toplevel_execute_ctrl4_down_LANE_AGE_lane0;
  reg        [11:0]   late0_BranchPlugin_logic_jumpLogic_history_fromFetch_shifter_4;
  reg        [11:0]   late0_BranchPlugin_logic_jumpLogic_history_fromFetch_shifter_3;
  reg        [11:0]   late0_BranchPlugin_logic_jumpLogic_history_fromFetch_shifter_2;
  reg        [11:0]   late0_BranchPlugin_logic_jumpLogic_history_fromFetch_shifter_1;
  wire       [3:0]    toplevel_execute_ctrl4_down_Prediction_ALIGNED_SLICES_TAKEN_lane0;
  wire       [3:0]    toplevel_execute_ctrl4_down_Prediction_ALIGNED_SLICES_BRANCH_lane0;
  wire       [11:0]   toplevel_execute_ctrl4_down_Prediction_BRANCH_HISTORY_lane0;
  wire       [31:0]   toplevel_execute_ctrl4_down_PC_lane0;
  wire                toplevel_execute_ctrl4_down_late0_BranchPlugin_SEL_lane0;
  wire                toplevel_execute_ctrl4_down_Prediction_ALIGNED_JUMPED_lane0;
  wire       [31:0]   toplevel_execute_ctrl4_down_late0_BranchPlugin_logic_jumpLogic_btb_REAL_TARGET_lane0;
  wire       [31:0]   toplevel_execute_ctrl4_down_early0_BranchPlugin_pcCalc_PC_FALSE_lane0;
  wire                toplevel_execute_ctrl4_down_late0_BranchPlugin_logic_jumpLogic_COND_lane0;
  wire       [31:0]   toplevel_execute_ctrl4_down_Decode_UOP_lane0;
  wire                toplevel_execute_ctrl4_down_late0_BranchPlugin_logic_alu_MSB_FAILED_lane0;
  wire       [1:0]    toplevel_execute_ctrl4_down_BranchPlugin_BRANCH_CTRL_lane0;
  wire                toplevel_execute_ctrl4_down_late0_BranchPlugin_logic_alu_btb_BAD_TARGET_lane0;
  wire       [31:0]   toplevel_execute_ctrl4_down_early0_BranchPlugin_pcCalc_PC_TRUE_lane0;
  wire       [31:0]   toplevel_execute_ctrl4_down_Prediction_ALIGNED_JUMPED_PC_lane0;
  wire                toplevel_execute_ctrl4_down_late0_BranchPlugin_logic_alu_EQ_lane0;
  wire                toplevel_execute_ctrl4_down_SrcStageables_UNSIGNED_lane1;
  wire                toplevel_execute_ctrl4_down_SrcStageables_ZERO_lane1;
  wire                toplevel_execute_ctrl4_down_SrcStageables_REVERT_lane1;
  wire       [31:0]   toplevel_execute_ctrl3_down_integer_RS2_lane1;
  wire       [1:0]    toplevel_execute_ctrl3_down_late1_SrcPlugin_logic_SRC2_CTRL_lane1;
  wire       [31:0]   toplevel_execute_ctrl3_down_late1_SrcPlugin_SRC2_lane1;
  wire       [31:0]   toplevel_execute_ctrl3_down_integer_RS1_lane1;
  wire       [0:0]    toplevel_execute_ctrl3_down_late1_SrcPlugin_logic_SRC1_CTRL_lane1;
  wire       [31:0]   toplevel_execute_ctrl3_down_late1_SrcPlugin_SRC1_lane1;
  reg                 toplevel_execute_ctrl4_up_LANE_SEL_lane1;
  reg                 toplevel_execute_ctrl2_up_LANE_SEL_lane1;
  wire                toplevel_execute_ctrl2_down_SrcStageables_UNSIGNED_lane1;
  wire                toplevel_execute_ctrl2_down_SrcStageables_ZERO_lane1;
  wire                toplevel_execute_ctrl2_down_SrcStageables_REVERT_lane1;
  wire       [31:0]   toplevel_execute_ctrl1_down_PC_lane1;
  wire       [31:0]   toplevel_execute_ctrl1_down_integer_RS2_lane1;
  wire       [1:0]    toplevel_execute_ctrl1_down_early1_SrcPlugin_logic_SRC2_CTRL_lane1;
  wire       [31:0]   toplevel_execute_ctrl1_down_early1_SrcPlugin_SRC2_lane1;
  wire       [31:0]   toplevel_execute_ctrl1_down_integer_RS1_lane1;
  wire       [0:0]    toplevel_execute_ctrl1_down_early1_SrcPlugin_logic_SRC1_CTRL_lane1;
  wire       [31:0]   toplevel_execute_ctrl1_down_early1_SrcPlugin_SRC1_lane1;
  wire       [31:0]   toplevel_execute_ctrl1_down_Decode_UOP_lane1;
  wire                toplevel_execute_ctrl4_down_SrcStageables_UNSIGNED_lane0;
  wire                toplevel_execute_ctrl4_down_SrcStageables_ZERO_lane0;
  wire                toplevel_execute_ctrl4_down_SrcStageables_REVERT_lane0;
  wire       [31:0]   toplevel_execute_ctrl3_down_integer_RS2_lane0;
  wire       [1:0]    toplevel_execute_ctrl3_down_late0_SrcPlugin_logic_SRC2_CTRL_lane0;
  wire       [31:0]   toplevel_execute_ctrl3_down_late0_SrcPlugin_SRC2_lane0;
  wire       [31:0]   toplevel_execute_ctrl3_down_integer_RS1_lane0;
  wire       [0:0]    toplevel_execute_ctrl3_down_late0_SrcPlugin_logic_SRC1_CTRL_lane0;
  wire       [31:0]   toplevel_execute_ctrl3_down_late0_SrcPlugin_SRC1_lane0;
  wire       [1:0]    toplevel_execute_ctrl4_down_lane0_IntFormatPlugin_logic_WIDTH_ID_lane0;
  wire                toplevel_execute_ctrl4_down_lane0_IntFormatPlugin_logic_SIGNED_lane0;
  wire                toplevel_execute_ctrl2_down_SrcStageables_UNSIGNED_lane0;
  wire                toplevel_execute_ctrl2_down_SrcStageables_ZERO_lane0;
  wire                toplevel_execute_ctrl2_down_SrcStageables_REVERT_lane0;
  wire       [31:0]   toplevel_execute_ctrl1_down_PC_lane0;
  wire       [31:0]   toplevel_execute_ctrl1_down_integer_RS2_lane0;
  wire       [1:0]    toplevel_execute_ctrl1_down_early0_SrcPlugin_logic_SRC2_CTRL_lane0;
  wire       [31:0]   toplevel_execute_ctrl1_down_early0_SrcPlugin_SRC2_lane0;
  wire       [31:0]   toplevel_execute_ctrl1_down_integer_RS1_lane0;
  wire       [0:0]    toplevel_execute_ctrl1_down_early0_SrcPlugin_logic_SRC1_CTRL_lane0;
  wire       [31:0]   toplevel_execute_ctrl1_down_early0_SrcPlugin_SRC1_lane0;
  wire       [31:0]   toplevel_execute_ctrl1_down_Decode_UOP_lane0;
  wire                toplevel_execute_ctrl2_down_early1_BranchPlugin_SEL_lane1;
  wire                toplevel_execute_ctrl3_down_early1_BranchPlugin_logic_jumpLogic_IS_JALR_lane1;
  wire                toplevel_execute_ctrl3_down_early1_BranchPlugin_logic_jumpLogic_IS_JAL_lane1;
  wire                toplevel_execute_ctrl3_down_early1_BranchPlugin_logic_jumpLogic_MISSALIGNED_lane1;
  wire       [15:0]   toplevel_execute_ctrl3_down_Decode_UOP_ID_lane1;
  wire       [0:0]    toplevel_execute_ctrl3_down_LANE_AGE_lane1;
  reg        [11:0]   early1_BranchPlugin_logic_jumpLogic_history_fromFetch_shifter_4;
  reg        [11:0]   early1_BranchPlugin_logic_jumpLogic_history_fromFetch_shifter_3;
  reg        [11:0]   early1_BranchPlugin_logic_jumpLogic_history_fromFetch_shifter_2;
  reg        [11:0]   early1_BranchPlugin_logic_jumpLogic_history_fromFetch_shifter_1;
  wire       [3:0]    toplevel_execute_ctrl3_down_Prediction_ALIGNED_SLICES_TAKEN_lane1;
  wire       [3:0]    toplevel_execute_ctrl3_down_Prediction_ALIGNED_SLICES_BRANCH_lane1;
  wire       [11:0]   toplevel_execute_ctrl3_down_Prediction_BRANCH_HISTORY_lane1;
  wire       [31:0]   toplevel_execute_ctrl3_down_PC_lane1;
  wire                toplevel_execute_ctrl3_down_early1_BranchPlugin_SEL_lane1;
  reg                 toplevel_execute_ctrl3_up_LANE_SEL_lane1;
  wire                toplevel_execute_ctrl3_down_early1_BranchPlugin_logic_alu_MSB_FAILED_lane1;
  wire                toplevel_execute_ctrl3_down_early1_BranchPlugin_logic_alu_btb_BAD_TARGET_lane1;
  wire                toplevel_execute_ctrl3_down_Prediction_ALIGNED_JUMPED_lane1;
  wire       [31:0]   toplevel_execute_ctrl3_down_early1_BranchPlugin_logic_jumpLogic_btb_REAL_TARGET_lane1;
  wire       [31:0]   toplevel_execute_ctrl3_down_early1_BranchPlugin_pcCalc_PC_FALSE_lane1;
  wire       [31:0]   toplevel_execute_ctrl3_down_early1_BranchPlugin_pcCalc_PC_TRUE_lane1;
  wire                toplevel_execute_ctrl3_down_early1_BranchPlugin_logic_jumpLogic_COND_lane1;
  wire                toplevel_execute_ctrl3_down_early1_SrcPlugin_LESS_lane1;
  wire                toplevel_execute_ctrl3_down_early1_BranchPlugin_logic_alu_EQ_lane1;
  wire       [31:0]   toplevel_execute_ctrl3_down_Decode_UOP_lane1;
  wire       [1:0]    toplevel_execute_ctrl3_down_BranchPlugin_BRANCH_CTRL_lane1;
  wire                toplevel_execute_ctrl2_down_early1_BranchPlugin_logic_alu_MSB_FAILED_lane1;
  wire                toplevel_execute_ctrl2_down_early1_BranchPlugin_logic_alu_btb_BAD_TARGET_lane1;
  wire       [31:0]   toplevel_execute_ctrl2_down_Prediction_ALIGNED_JUMPED_PC_lane1;
  wire                toplevel_execute_ctrl2_down_early1_BranchPlugin_logic_alu_EQ_lane1;
  wire                toplevel_execute_ctrl2_up_COMMIT_lane0;
  wire                toplevel_execute_ctrl2_down_COMMIT_lane0;
  reg                 toplevel_execute_ctrl2_COMMIT_lane0_bypass;
  reg                 toplevel_execute_ctrl2_up_TRAP_lane0;
  wire                toplevel_execute_ctrl2_down_TRAP_lane0;
  reg                 toplevel_execute_ctrl2_TRAP_lane0_bypass;
  wire                toplevel_execute_ctrl2_down_early0_EnvPlugin_SEL_lane0;
  wire       [2:0]    toplevel_execute_ctrl2_down_early0_EnvPlugin_OP_lane0;
  wire       [0:0]    toplevel_execute_ctrl2_down_LANE_AGE_lane0;
  wire       [15:0]   toplevel_execute_ctrl2_down_Decode_UOP_ID_lane0;
  wire                toplevel_execute_ctrl2_down_early0_BranchPlugin_SEL_lane0;
  wire                toplevel_execute_ctrl3_down_early0_BranchPlugin_logic_jumpLogic_IS_JALR_lane0;
  wire                toplevel_execute_ctrl3_down_early0_BranchPlugin_logic_jumpLogic_IS_JAL_lane0;
  wire                toplevel_execute_ctrl3_down_early0_BranchPlugin_logic_jumpLogic_MISSALIGNED_lane0;
  wire       [15:0]   toplevel_execute_ctrl3_down_Decode_UOP_ID_lane0;
  wire       [0:0]    toplevel_execute_ctrl3_down_LANE_AGE_lane0;
  reg        [11:0]   early0_BranchPlugin_logic_jumpLogic_history_fromFetch_shifter_4;
  reg        [11:0]   early0_BranchPlugin_logic_jumpLogic_history_fromFetch_shifter_3;
  reg        [11:0]   early0_BranchPlugin_logic_jumpLogic_history_fromFetch_shifter_2;
  reg        [11:0]   early0_BranchPlugin_logic_jumpLogic_history_fromFetch_shifter_1;
  wire       [3:0]    toplevel_execute_ctrl3_down_Prediction_ALIGNED_SLICES_TAKEN_lane0;
  wire       [3:0]    toplevel_execute_ctrl3_down_Prediction_ALIGNED_SLICES_BRANCH_lane0;
  wire       [11:0]   toplevel_execute_ctrl3_down_Prediction_BRANCH_HISTORY_lane0;
  wire       [31:0]   toplevel_execute_ctrl3_down_PC_lane0;
  wire                toplevel_execute_ctrl3_down_early0_BranchPlugin_SEL_lane0;
  reg                 toplevel_execute_ctrl3_up_LANE_SEL_lane0;
  wire                toplevel_execute_ctrl3_down_early0_BranchPlugin_logic_alu_MSB_FAILED_lane0;
  wire                toplevel_execute_ctrl3_down_early0_BranchPlugin_logic_alu_btb_BAD_TARGET_lane0;
  wire                toplevel_execute_ctrl3_down_Prediction_ALIGNED_JUMPED_lane0;
  wire       [31:0]   toplevel_execute_ctrl3_down_early0_BranchPlugin_logic_jumpLogic_btb_REAL_TARGET_lane0;
  wire       [31:0]   toplevel_execute_ctrl3_down_early0_BranchPlugin_pcCalc_PC_FALSE_lane0;
  wire       [31:0]   toplevel_execute_ctrl3_down_early0_BranchPlugin_pcCalc_PC_TRUE_lane0;
  wire                toplevel_execute_ctrl3_down_early0_BranchPlugin_logic_jumpLogic_COND_lane0;
  wire                toplevel_execute_ctrl3_down_early0_SrcPlugin_LESS_lane0;
  wire                toplevel_execute_ctrl3_down_early0_BranchPlugin_logic_alu_EQ_lane0;
  wire       [31:0]   toplevel_execute_ctrl3_down_Decode_UOP_lane0;
  wire       [1:0]    toplevel_execute_ctrl3_down_BranchPlugin_BRANCH_CTRL_lane0;
  wire                toplevel_execute_ctrl2_down_early0_BranchPlugin_logic_alu_MSB_FAILED_lane0;
  wire                toplevel_execute_ctrl2_down_early0_BranchPlugin_logic_alu_btb_BAD_TARGET_lane0;
  wire       [31:0]   toplevel_execute_ctrl2_down_Prediction_ALIGNED_JUMPED_PC_lane0;
  wire                toplevel_execute_ctrl2_down_early0_BranchPlugin_logic_alu_EQ_lane0;
  wire                toplevel_decode_ctrls_1_lane0_upIsCancel;
  wire                toplevel_decode_ctrls_1_lane0_downIsCancel;
  wire       [9:0]    toplevel_decode_ctrls_0_down_Fetch_ID_1;
  wire       [31:0]   toplevel_decode_ctrls_0_down_PC_1;
  wire       [9:0]    toplevel_decode_ctrls_0_down_Fetch_ID_0;
  wire       [31:0]   toplevel_decode_ctrls_0_down_PC_0;
  wire       [9:0]    fetch_logic_ctrls_0_down_Fetch_ID;
  reg                 _zz_5;
  reg        [1:0]    BtbPlugin_logic_ras_ptr_pop_aheadValue;
  wire       [11:0]   fetch_logic_ctrls_1_down_GSharePlugin_logic_HASH;
  wire                fetch_logic_ctrls_1_down_GSharePlugin_logic_BYPASS_valid;
  wire       [11:0]   fetch_logic_ctrls_1_down_GSharePlugin_logic_BYPASS_payload_address;
  wire       [1:0]    fetch_logic_ctrls_1_down_GSharePlugin_logic_BYPASS_payload_data_0;
  wire       [1:0]    fetch_logic_ctrls_1_down_GSharePlugin_logic_BYPASS_payload_data_1;
  wire       [1:0]    fetch_logic_ctrls_1_down_GSharePlugin_logic_BYPASS_payload_data_2;
  wire       [1:0]    fetch_logic_ctrls_1_down_GSharePlugin_logic_BYPASS_payload_data_3;
  wire                fetch_logic_ctrls_0_down_isReady;
  (* keep , syn_keep *) reg        [1:0]    fetch_logic_ctrls_1_down_GSharePlugin_GSHARE_COUNTER_0 /* synthesis syn_keep = 1 */ ;
  (* keep , syn_keep *) reg        [1:0]    fetch_logic_ctrls_1_down_GSharePlugin_GSHARE_COUNTER_1 /* synthesis syn_keep = 1 */ ;
  (* keep , syn_keep *) reg        [1:0]    fetch_logic_ctrls_1_down_GSharePlugin_GSHARE_COUNTER_2 /* synthesis syn_keep = 1 */ ;
  (* keep , syn_keep *) reg        [1:0]    fetch_logic_ctrls_1_down_GSharePlugin_GSHARE_COUNTER_3 /* synthesis syn_keep = 1 */ ;
  wire                fetch_logic_ctrls_0_down_GSharePlugin_logic_BYPASS_valid;
  wire       [11:0]   fetch_logic_ctrls_0_down_GSharePlugin_logic_BYPASS_payload_address;
  wire       [1:0]    fetch_logic_ctrls_0_down_GSharePlugin_logic_BYPASS_payload_data_0;
  wire       [1:0]    fetch_logic_ctrls_0_down_GSharePlugin_logic_BYPASS_payload_data_1;
  wire       [1:0]    fetch_logic_ctrls_0_down_GSharePlugin_logic_BYPASS_payload_data_2;
  wire       [1:0]    fetch_logic_ctrls_0_down_GSharePlugin_logic_BYPASS_payload_data_3;
  wire       [11:0]   fetch_logic_ctrls_0_down_Prediction_BRANCH_HISTORY;
  wire       [11:0]   fetch_logic_ctrls_0_down_GSharePlugin_logic_HASH;
  reg                 _zz_6;
  wire                toplevel_execute_ctrl4_down_LsuL1_FLUSH_lane0;
  wire                toplevel_execute_ctrl4_down_LsuL1_SEL_lane0;
  wire                toplevel_execute_ctrl3_down_LsuL1_FLUSH_lane0;
  wire                toplevel_execute_ctrl3_down_LsuL1_SEL_lane0;
  wire       [31:0]   toplevel_execute_ctrl0_down_Decode_UOP_lane0;
  wire       [1:0]    toplevel_execute_ctrl0_down_AguPlugin_SIZE_lane0;
  wire                fetch_logic_ctrls_2_up_isCanceling;
  wire                fetch_logic_ctrls_2_down_MMU_BYPASS_TRANSLATION;
  wire                fetch_logic_ctrls_2_down_Fetch_PC_FAULT;
  wire                fetch_logic_ctrls_2_down_MMU_HAZARD;
  wire                fetch_logic_ctrls_2_down_MMU_REFILL;
  wire                fetch_logic_ctrls_2_down_MMU_ACCESS_FAULT;
  wire                fetch_logic_ctrls_2_down_MMU_ALLOW_EXECUTE;
  wire                fetch_logic_ctrls_2_down_MMU_PAGE_FAULT;
  wire                fetch_logic_ctrls_2_down_FetchL1Plugin_logic_WAYS_HIT;
  wire                fetch_logic_ctrls_2_up_isCancel;
  wire                fetch_logic_ctrls_2_down_FetchL1Plugin_logic_HAZARD;
  wire                fetch_logic_ctrls_2_down_FetchL1Plugin_logic_WAYS_TAGS_0_loaded;
  wire                fetch_logic_ctrls_2_down_FetchL1Plugin_logic_WAYS_TAGS_0_error;
  wire       [19:0]   fetch_logic_ctrls_2_down_FetchL1Plugin_logic_WAYS_TAGS_0_address;
  wire                fetch_logic_ctrls_2_down_FetchL1Plugin_logic_WAYS_TAGS_1_loaded;
  wire                fetch_logic_ctrls_2_down_FetchL1Plugin_logic_WAYS_TAGS_1_error;
  wire       [19:0]   fetch_logic_ctrls_2_down_FetchL1Plugin_logic_WAYS_TAGS_1_address;
  wire                fetch_logic_ctrls_2_up_isReady;
  wire       [0:0]    fetch_logic_ctrls_2_down_FetchL1Plugin_logic_PLRU_BYPASSED_0;
  wire       [31:0]   fetch_logic_ctrls_2_down_MMU_TRANSLATED;
  wire                fetch_logic_ctrls_1_down_FetchL1Plugin_logic_WAYS_HIT;
  wire                fetch_logic_ctrls_1_down_MMU_BYPASS_TRANSLATION;
  wire                fetch_logic_ctrls_1_down_FetchL1Plugin_logic_WAYS_HITS_0;
  wire                fetch_logic_ctrls_1_down_FetchL1Plugin_logic_WAYS_HITS_1;
  wire       [2:0]    fetch_logic_ctrls_1_down_MMU_WAYS_OH;
  wire       [31:0]   fetch_logic_ctrls_1_down_MMU_WAYS_PHYSICAL_0;
  wire       [31:0]   fetch_logic_ctrls_1_down_MMU_WAYS_PHYSICAL_1;
  wire       [31:0]   fetch_logic_ctrls_1_down_MMU_WAYS_PHYSICAL_2;
  wire       [5:0]    fetch_logic_ctrls_1_down_FetchL1Plugin_logic_cmd_TAGS_UPDATE_ADDRESS;
  wire                fetch_logic_ctrls_1_down_FetchL1Plugin_logic_cmd_TAGS_UPDATE;
  wire                fetch_logic_ctrls_1_down_FetchL1Plugin_logic_HAZARD;
  wire       [63:0]   fetch_logic_ctrls_2_down_FetchL1Plugin_logic_BANKS_MUXES_0;
  wire       [63:0]   fetch_logic_ctrls_2_down_FetchL1Plugin_logic_BANKS_MUXES_1;
  wire                fetch_logic_ctrls_2_down_FetchL1Plugin_logic_WAYS_HITS_0;
  wire                fetch_logic_ctrls_2_down_FetchL1Plugin_logic_WAYS_HITS_1;
  wire       [31:0]   fetch_logic_ctrls_1_down_Fetch_WORD_PC;
  wire       [63:0]   fetch_logic_ctrls_1_down_FetchL1Plugin_logic_BANKS_MUXES_0;
  wire       [63:0]   fetch_logic_ctrls_1_down_FetchL1Plugin_logic_BANKS_MUXES_1;
  wire       [0:0]    fetch_logic_ctrls_1_down_FetchL1Plugin_logic_cmd_PLRU_BYPASS_DATA_0;
  wire                fetch_logic_ctrls_1_down_FetchL1Plugin_logic_cmd_PLRU_BYPASS_VALID;
  reg        [0:0]    fetch_logic_ctrls_1_down_FetchL1Plugin_logic_PLRU_BYPASSED_0;
  wire       [5:0]    fetch_logic_ctrls_0_down_FetchL1Plugin_logic_cmd_TAGS_UPDATE_ADDRESS;
  wire                fetch_logic_ctrls_0_down_FetchL1Plugin_logic_cmd_TAGS_UPDATE;
  wire       [0:0]    fetch_logic_ctrls_0_down_FetchL1Plugin_logic_cmd_PLRU_BYPASS_DATA_0;
  wire                fetch_logic_ctrls_0_down_FetchL1Plugin_logic_cmd_PLRU_BYPASS_VALID;
  reg                 fetch_logic_ctrls_1_up_valid;
  wire                fetch_logic_ctrls_1_up_ready;
  wire       [31:0]   fetch_logic_ctrls_0_down_Fetch_WORD_PC;
  reg                 _zz_fetch_logic_ctrls_0_haltRequest_FetchL1Plugin_l233;
  wire       [0:0]    fetch_logic_ctrls_1_down_FetchL1Plugin_logic_PLRU_READ_0;
  reg                 _zz_7;
  wire                fetch_logic_ctrls_1_down_FetchL1Plugin_logic_WAYS_TAGS_0_loaded;
  wire                fetch_logic_ctrls_1_down_FetchL1Plugin_logic_WAYS_TAGS_0_error;
  wire       [19:0]   fetch_logic_ctrls_1_down_FetchL1Plugin_logic_WAYS_TAGS_0_address;
  wire                fetch_logic_ctrls_1_down_FetchL1Plugin_logic_WAYS_TAGS_1_loaded;
  wire                fetch_logic_ctrls_1_down_FetchL1Plugin_logic_WAYS_TAGS_1_error;
  wire       [19:0]   fetch_logic_ctrls_1_down_FetchL1Plugin_logic_WAYS_TAGS_1_address;
  reg                 _zz_8;
  wire       [63:0]   fetch_logic_ctrls_1_down_FetchL1Plugin_logic_BANKS_WORDS_0;
  wire       [63:0]   fetch_logic_ctrls_1_down_FetchL1Plugin_logic_BANKS_WORDS_1;
  reg                 _zz_9;
  wire       [31:0]   fetch_logic_ctrls_2_down_Prediction_WORD_JUMP_PC;
  reg        [3:0]    fetch_logic_ctrls_2_down_Prediction_WORD_SLICES_TAKEN;
  reg        [3:0]    fetch_logic_ctrls_2_down_Prediction_WORD_SLICES_BRANCH;
  wire       [11:0]   fetch_logic_ctrls_2_down_Prediction_BRANCH_HISTORY;
  wire       [1:0]    fetch_logic_ctrls_2_down_GSharePlugin_GSHARE_COUNTER_0;
  wire       [1:0]    fetch_logic_ctrls_2_down_GSharePlugin_GSHARE_COUNTER_1;
  wire       [1:0]    fetch_logic_ctrls_2_down_GSharePlugin_GSHARE_COUNTER_2;
  wire       [1:0]    fetch_logic_ctrls_2_down_GSharePlugin_GSHARE_COUNTER_3;
  wire       [9:0]    fetch_logic_ctrls_2_down_Fetch_ID;
  wire                fetch_logic_ctrls_2_down_TRAP;
  wire                fetch_logic_ctrls_2_down_isCancel;
  wire                fetch_logic_ctrls_2_down_isReady;
  wire                fetch_logic_ctrls_2_down_isValid;
  wire                fetch_logic_ctrls_2_down_ready;
  wire                toplevel_decode_ctrls_0_up_isCancel;
  wire                toplevel_decode_ctrls_0_up_isReady;
  wire                fetch_logic_ctrls_2_down_valid;
  wire       [63:0]   fetch_logic_ctrls_2_down_Fetch_WORD;
  wire                toplevel_decode_ctrls_0_up_valid;
  wire                toplevel_decode_ctrls_0_up_Prediction_ALIGN_REDO_1;
  wire       [3:0]    toplevel_decode_ctrls_0_up_Prediction_ALIGNED_SLICES_TAKEN_1;
  wire       [3:0]    toplevel_decode_ctrls_0_up_Prediction_ALIGNED_SLICES_BRANCH_1;
  wire       [31:0]   toplevel_decode_ctrls_0_up_Prediction_ALIGNED_JUMPED_PC_1;
  wire                toplevel_decode_ctrls_0_up_Prediction_ALIGNED_JUMPED_1;
  wire                toplevel_decode_ctrls_0_up_TRAP_1;
  wire       [1:0]    toplevel_decode_ctrls_0_up_Prediction_WORD_JUMP_SLICE_1;
  wire                toplevel_decode_ctrls_0_up_Prediction_WORD_JUMPED_1;
  wire       [31:0]   toplevel_decode_ctrls_0_up_Prediction_WORD_JUMP_PC_1;
  wire       [3:0]    toplevel_decode_ctrls_0_up_Prediction_WORD_SLICES_TAKEN_1;
  wire       [3:0]    toplevel_decode_ctrls_0_up_Prediction_WORD_SLICES_BRANCH_1;
  wire       [11:0]   toplevel_decode_ctrls_0_up_Prediction_BRANCH_HISTORY_1;
  wire       [1:0]    toplevel_decode_ctrls_0_up_GSharePlugin_GSHARE_COUNTER_1_0;
  wire       [1:0]    toplevel_decode_ctrls_0_up_GSharePlugin_GSHARE_COUNTER_1_1;
  wire       [1:0]    toplevel_decode_ctrls_0_up_GSharePlugin_GSHARE_COUNTER_1_2;
  wire       [1:0]    toplevel_decode_ctrls_0_up_GSharePlugin_GSHARE_COUNTER_1_3;
  wire       [9:0]    toplevel_decode_ctrls_0_up_Fetch_ID_1;
  wire       [9:0]    toplevel_decode_ctrls_0_down_Decode_DOP_ID_0;
  wire       [9:0]    toplevel_decode_ctrls_0_up_Decode_DOP_ID_1;
  wire       [31:0]   toplevel_decode_ctrls_0_up_PC_1;
  wire       [0:0]    toplevel_decode_ctrls_0_up_Decode_INSTRUCTION_SLICE_COUNT_1;
  reg        [31:0]   toplevel_decode_ctrls_0_up_Decode_INSTRUCTION_RAW_1;
  reg                 toplevel_decode_ctrls_0_up_Decode_DECOMPRESSION_FAULT_1;
  reg        [31:0]   toplevel_decode_ctrls_0_up_Decode_INSTRUCTION_1;
  wire                toplevel_decode_ctrls_0_up_LANE_SEL_1;
  wire                toplevel_decode_ctrls_0_up_Prediction_ALIGN_REDO_0;
  wire       [3:0]    toplevel_decode_ctrls_0_up_Prediction_ALIGNED_SLICES_TAKEN_0;
  wire       [3:0]    toplevel_decode_ctrls_0_up_Prediction_ALIGNED_SLICES_BRANCH_0;
  wire       [31:0]   toplevel_decode_ctrls_0_up_Prediction_ALIGNED_JUMPED_PC_0;
  wire                toplevel_decode_ctrls_0_up_Prediction_ALIGNED_JUMPED_0;
  wire                toplevel_decode_ctrls_0_up_TRAP_0;
  wire       [1:0]    toplevel_decode_ctrls_0_up_Prediction_WORD_JUMP_SLICE_0;
  wire                toplevel_decode_ctrls_0_up_Prediction_WORD_JUMPED_0;
  wire       [31:0]   toplevel_decode_ctrls_0_up_Prediction_WORD_JUMP_PC_0;
  wire       [3:0]    toplevel_decode_ctrls_0_up_Prediction_WORD_SLICES_TAKEN_0;
  wire       [3:0]    toplevel_decode_ctrls_0_up_Prediction_WORD_SLICES_BRANCH_0;
  wire       [11:0]   toplevel_decode_ctrls_0_up_Prediction_BRANCH_HISTORY_0;
  wire       [1:0]    toplevel_decode_ctrls_0_up_GSharePlugin_GSHARE_COUNTER_0_0;
  wire       [1:0]    toplevel_decode_ctrls_0_up_GSharePlugin_GSHARE_COUNTER_0_1;
  wire       [1:0]    toplevel_decode_ctrls_0_up_GSharePlugin_GSHARE_COUNTER_0_2;
  wire       [1:0]    toplevel_decode_ctrls_0_up_GSharePlugin_GSHARE_COUNTER_0_3;
  wire       [9:0]    toplevel_decode_ctrls_0_up_Fetch_ID_0;
  wire       [9:0]    toplevel_decode_ctrls_0_up_Decode_DOP_ID_0;
  wire       [31:0]   toplevel_decode_ctrls_0_up_PC_0;
  wire       [0:0]    toplevel_decode_ctrls_0_up_Decode_INSTRUCTION_SLICE_COUNT_0;
  reg        [31:0]   toplevel_decode_ctrls_0_up_Decode_INSTRUCTION_RAW_0;
  reg                 toplevel_decode_ctrls_0_up_Decode_DECOMPRESSION_FAULT_0;
  reg        [31:0]   toplevel_decode_ctrls_0_up_Decode_INSTRUCTION_0;
  wire                toplevel_decode_ctrls_0_up_LANE_SEL_0;
  wire                toplevel_decode_ctrls_0_lane0_upIsCancel;
  wire                toplevel_decode_ctrls_0_lane0_downIsCancel;
  wire       [9:0]    toplevel_decode_ctrls_0_down_Decode_DOP_ID_1;
  wire                toplevel_decode_ctrls_0_lane1_upIsCancel;
  wire                toplevel_decode_ctrls_0_lane1_downIsCancel;
  wire                toplevel_decode_ctrls_0_up_isFiring;
  wire                fetch_logic_ctrls_2_up_isValid;
  wire       [3:0]    fetch_logic_ctrls_2_down_AlignerPlugin_logic_FETCH_LAST;
  wire                fetch_logic_ctrls_2_down_Prediction_WORD_JUMPED;
  wire       [1:0]    fetch_logic_ctrls_2_down_Prediction_WORD_JUMP_SLICE;
  wire       [31:0]   fetch_logic_ctrls_2_down_Fetch_WORD_PC;
  wire       [3:0]    fetch_logic_ctrls_2_down_AlignerPlugin_logic_FETCH_MASK;
  (* keep , syn_keep *) wire       [31:0]   toplevel_execute_ctrl2_down_early1_BranchPlugin_pcCalc_PC_LAST_SLICE_lane1 /* synthesis syn_keep = 1 */ ;
  (* keep , syn_keep *) wire       [31:0]   toplevel_execute_ctrl2_down_early1_BranchPlugin_pcCalc_PC_FALSE_lane1 /* synthesis syn_keep = 1 */ ;
  (* keep , syn_keep *) reg        [31:0]   toplevel_execute_ctrl2_down_early1_BranchPlugin_pcCalc_PC_TRUE_lane1 /* synthesis syn_keep = 1 */ ;
  wire       [0:0]    toplevel_execute_ctrl2_down_Decode_INSTRUCTION_SLICE_COUNT_lane1;
  wire       [31:0]   toplevel_execute_ctrl2_down_PC_lane1;
  wire       [1:0]    toplevel_execute_ctrl2_down_BranchPlugin_BRANCH_CTRL_lane1;
  wire       [31:0]   toplevel_execute_ctrl2_down_Decode_UOP_lane1;
  (* keep , syn_keep *) wire       [31:0]   toplevel_execute_ctrl2_down_early0_BranchPlugin_pcCalc_PC_LAST_SLICE_lane0 /* synthesis syn_keep = 1 */ ;
  (* keep , syn_keep *) wire       [31:0]   toplevel_execute_ctrl2_down_early0_BranchPlugin_pcCalc_PC_FALSE_lane0 /* synthesis syn_keep = 1 */ ;
  (* keep , syn_keep *) reg        [31:0]   toplevel_execute_ctrl2_down_early0_BranchPlugin_pcCalc_PC_TRUE_lane0 /* synthesis syn_keep = 1 */ ;
  wire       [0:0]    toplevel_execute_ctrl2_down_Decode_INSTRUCTION_SLICE_COUNT_lane0;
  wire       [31:0]   toplevel_execute_ctrl2_down_PC_lane0;
  wire       [1:0]    toplevel_execute_ctrl2_down_BranchPlugin_BRANCH_CTRL_lane0;
  wire       [31:0]   toplevel_execute_ctrl2_down_Decode_UOP_lane0;
  wire                fetch_logic_ctrls_0_down_isFiring;
  wire                toplevel_execute_ctrl4_down_late1_BarrelShifterPlugin_SEL_lane1;
  wire       [31:0]   toplevel_execute_ctrl4_down_late1_BarrelShifterPlugin_SHIFT_RESULT_lane1;
  wire                toplevel_execute_ctrl4_down_BarrelShifterPlugin_SIGNED_lane1;
  wire                toplevel_execute_ctrl4_down_BarrelShifterPlugin_LEFT_lane1;
  wire                toplevel_execute_ctrl4_down_late1_IntAluPlugin_SEL_lane1;
  wire       [31:0]   toplevel_execute_ctrl4_down_late1_IntAluPlugin_ALU_RESULT_lane1;
  wire                toplevel_execute_ctrl4_down_late1_IntAluPlugin_ALU_SLTX_lane1;
  wire                toplevel_execute_ctrl4_down_late1_SrcPlugin_LESS_lane1;
  wire                toplevel_execute_ctrl4_down_late1_IntAluPlugin_ALU_ADD_SUB_lane1;
  wire       [31:0]   toplevel_execute_ctrl4_down_late1_SrcPlugin_ADD_SUB_lane1;
  wire       [31:0]   toplevel_execute_ctrl4_down_late1_SrcPlugin_SRC2_lane1;
  wire       [31:0]   toplevel_execute_ctrl4_down_late1_SrcPlugin_SRC1_lane1;
  wire       [1:0]    toplevel_execute_ctrl4_down_late1_IntAluPlugin_ALU_BITWISE_CTRL_lane1;
  wire       [31:0]   toplevel_execute_ctrl3_down_early1_BarrelShifterPlugin_SHIFT_RESULT_lane1;
  wire                toplevel_execute_ctrl3_down_early1_BarrelShifterPlugin_SEL_lane1;
  wire       [31:0]   toplevel_execute_ctrl2_down_early1_BarrelShifterPlugin_SHIFT_RESULT_lane1;
  wire                toplevel_execute_ctrl2_down_BarrelShifterPlugin_SIGNED_lane1;
  wire                toplevel_execute_ctrl2_down_BarrelShifterPlugin_LEFT_lane1;
  wire                toplevel_execute_ctrl2_down_early1_IntAluPlugin_SEL_lane1;
  wire       [31:0]   toplevel_execute_ctrl2_down_early1_IntAluPlugin_ALU_RESULT_lane1;
  wire                toplevel_execute_ctrl2_down_early1_IntAluPlugin_ALU_SLTX_lane1;
  wire                toplevel_execute_ctrl2_down_early1_SrcPlugin_LESS_lane1;
  wire                toplevel_execute_ctrl2_down_early1_IntAluPlugin_ALU_ADD_SUB_lane1;
  wire       [31:0]   toplevel_execute_ctrl2_down_early1_SrcPlugin_ADD_SUB_lane1;
  wire       [31:0]   toplevel_execute_ctrl2_down_early1_SrcPlugin_SRC2_lane1;
  wire       [31:0]   toplevel_execute_ctrl2_down_early1_SrcPlugin_SRC1_lane1;
  wire       [1:0]    toplevel_execute_ctrl2_down_early1_IntAluPlugin_ALU_BITWISE_CTRL_lane1;
  wire                toplevel_execute_ctrl4_down_late0_BarrelShifterPlugin_SEL_lane0;
  wire       [31:0]   toplevel_execute_ctrl4_down_late0_BarrelShifterPlugin_SHIFT_RESULT_lane0;
  wire                toplevel_execute_ctrl4_down_BarrelShifterPlugin_SIGNED_lane0;
  wire                toplevel_execute_ctrl4_down_BarrelShifterPlugin_LEFT_lane0;
  wire                toplevel_execute_ctrl4_down_late0_IntAluPlugin_SEL_lane0;
  wire       [31:0]   toplevel_execute_ctrl4_down_late0_IntAluPlugin_ALU_RESULT_lane0;
  wire                toplevel_execute_ctrl4_down_late0_IntAluPlugin_ALU_SLTX_lane0;
  wire                toplevel_execute_ctrl4_down_late0_SrcPlugin_LESS_lane0;
  wire                toplevel_execute_ctrl4_down_late0_IntAluPlugin_ALU_ADD_SUB_lane0;
  wire       [31:0]   toplevel_execute_ctrl4_down_late0_SrcPlugin_ADD_SUB_lane0;
  wire       [31:0]   toplevel_execute_ctrl4_down_late0_SrcPlugin_SRC2_lane0;
  wire       [31:0]   toplevel_execute_ctrl4_down_late0_SrcPlugin_SRC1_lane0;
  wire       [1:0]    toplevel_execute_ctrl4_down_late0_IntAluPlugin_ALU_BITWISE_CTRL_lane0;
  wire       [31:0]   toplevel_execute_ctrl3_down_DivPlugin_DIV_RESULT_lane0;
  wire                toplevel_execute_ctrl3_down_early0_DivPlugin_SEL_lane0;
  wire       [31:0]   toplevel_execute_ctrl2_down_DivPlugin_DIV_RESULT_lane0;
  wire                toplevel_execute_ctrl2_down_early0_DivPlugin_SEL_lane0;
  reg                 toplevel_execute_ctrl2_up_LANE_SEL_lane0;
  wire                toplevel_execute_ctrl2_down_isReady;
  wire                toplevel_execute_ctrl2_down_DivPlugin_REM_lane0;
  wire       [31:0]   toplevel_execute_ctrl2_down_RsUnsignedPlugin_RS2_UNSIGNED_lane0;
  wire       [31:0]   toplevel_execute_ctrl2_down_RsUnsignedPlugin_RS1_UNSIGNED_lane0;
  wire                toplevel_execute_ctrl2_down_RsUnsignedPlugin_RS2_REVERT_lane0;
  wire                toplevel_execute_ctrl2_down_RsUnsignedPlugin_RS1_REVERT_lane0;
  wire       [31:0]   toplevel_execute_ctrl2_down_RsUnsignedPlugin_RS2_FORMATED_lane0;
  wire       [31:0]   toplevel_execute_ctrl2_down_RsUnsignedPlugin_RS1_FORMATED_lane0;
  wire                toplevel_execute_ctrl4_down_early0_MulPlugin_SEL_lane0;
  wire                toplevel_execute_ctrl4_down_MulPlugin_HIGH_lane0;
  wire                toplevel_execute_ctrl4_down_isReady;
  reg                 toplevel_execute_ctrl4_up_LANE_SEL_lane0;
  wire       [65:0]   toplevel_execute_ctrl4_down_early0_MulPlugin_logic_steps_1_adders_0_lane0;
  wire       [4:0]    toplevel_execute_ctrl4_down_early0_MulPlugin_logic_steps_0_adders_1_lane0;
  wire       [62:0]   toplevel_execute_ctrl4_down_early0_MulPlugin_logic_steps_0_adders_0_lane0;
  wire       [4:0]    toplevel_execute_ctrl3_down_early0_MulPlugin_logic_steps_0_adders_1_lane0;
  wire       [62:0]   toplevel_execute_ctrl3_down_early0_MulPlugin_logic_steps_0_adders_0_lane0;
  wire       [29:0]   toplevel_execute_ctrl3_down_early0_MulPlugin_logic_mul_VALUES_3_lane0;
  wire       [46:0]   toplevel_execute_ctrl3_down_early0_MulPlugin_logic_mul_VALUES_2_lane0;
  wire       [46:0]   toplevel_execute_ctrl3_down_early0_MulPlugin_logic_mul_VALUES_1_lane0;
  wire       [33:0]   toplevel_execute_ctrl3_down_early0_MulPlugin_logic_mul_VALUES_0_lane0;
  wire       [32:0]   toplevel_execute_ctrl3_down_MUL_SRC2_lane0;
  wire       [32:0]   toplevel_execute_ctrl3_down_MUL_SRC1_lane0;
  wire                toplevel_execute_ctrl2_down_RsUnsignedPlugin_RS2_SIGNED_lane0;
  wire       [32:0]   toplevel_execute_ctrl2_down_MUL_SRC2_lane0;
  wire                toplevel_execute_ctrl2_down_RsUnsignedPlugin_RS1_SIGNED_lane0;
  wire       [32:0]   toplevel_execute_ctrl2_down_MUL_SRC1_lane0;
  reg        [31:0]   toplevel_execute_ctrl2_up_integer_RS2_lane0;
  reg        [31:0]   toplevel_execute_ctrl2_up_integer_RS1_lane0;
  wire       [31:0]   toplevel_execute_ctrl3_down_early0_BarrelShifterPlugin_SHIFT_RESULT_lane0;
  wire                toplevel_execute_ctrl3_down_early0_BarrelShifterPlugin_SEL_lane0;
  wire       [31:0]   toplevel_execute_ctrl2_down_early0_BarrelShifterPlugin_SHIFT_RESULT_lane0;
  wire                toplevel_execute_ctrl2_down_BarrelShifterPlugin_SIGNED_lane0;
  wire                toplevel_execute_ctrl2_down_BarrelShifterPlugin_LEFT_lane0;
  wire                toplevel_execute_ctrl2_down_early0_IntAluPlugin_SEL_lane0;
  wire       [31:0]   toplevel_execute_ctrl2_down_early0_IntAluPlugin_ALU_RESULT_lane0;
  wire                toplevel_execute_ctrl2_down_early0_IntAluPlugin_ALU_SLTX_lane0;
  wire                toplevel_execute_ctrl2_down_early0_SrcPlugin_LESS_lane0;
  wire                toplevel_execute_ctrl2_down_early0_IntAluPlugin_ALU_ADD_SUB_lane0;
  wire       [31:0]   toplevel_execute_ctrl2_down_early0_SrcPlugin_ADD_SUB_lane0;
  wire       [31:0]   toplevel_execute_ctrl2_down_early0_SrcPlugin_SRC2_lane0;
  wire       [31:0]   toplevel_execute_ctrl2_down_early0_SrcPlugin_SRC1_lane0;
  wire       [1:0]    toplevel_execute_ctrl2_down_early0_IntAluPlugin_ALU_BITWISE_CTRL_lane0;
  reg                 MmuPlugin_api_fetchTranslationEnable;
  reg                 MmuPlugin_api_lsuTranslationEnable;
  wire                AlignerPlugin_api_singleFetch;
  wire                AlignerPlugin_api_downMoving;
  wire                AlignerPlugin_api_haltIt;
  reg                 DispatchPlugin_api_haltDispatch;
  wire                execute_freeze_valid;
  wire       [0:0]    execute_lane0_api_hartsInflight;
  wire                toplevel_execute_lane0_ctrls_2_upIsCancel;
  wire                toplevel_execute_lane0_ctrls_2_downIsCancel;
  wire                CsrRamPlugin_api_holdRead;
  wire                CsrRamPlugin_api_holdWrite;
  reg                 CsrAccessPlugin_bus_decode_exception;
  wire                CsrAccessPlugin_bus_decode_read;
  wire                CsrAccessPlugin_bus_decode_write;
  wire       [11:0]   CsrAccessPlugin_bus_decode_address;
  reg                 CsrAccessPlugin_bus_decode_trap;
  wire                PrivilegedPlugin_api_lsuTriggerBus_load;
  wire                PrivilegedPlugin_api_lsuTriggerBus_store;
  reg                 TrapPlugin_api_harts_0_redo;
  reg                 TrapPlugin_api_harts_0_askWake;
  reg                 TrapPlugin_api_harts_0_rvTrap;
  wire                TrapPlugin_api_harts_0_fsmBusy;
  wire       [0:0]    execute_lane1_api_hartsInflight;
  wire                toplevel_execute_lane1_ctrls_2_upIsCancel;
  wire                toplevel_execute_lane1_ctrls_2_downIsCancel;
  reg                 MmuPlugin_logic_accessBus_cmd_valid;
  wire                MmuPlugin_logic_accessBus_cmd_ready;
  wire       [31:0]   MmuPlugin_logic_accessBus_cmd_payload_address;
  wire       [1:0]    MmuPlugin_logic_accessBus_cmd_payload_size;
  wire                MmuPlugin_logic_accessBus_rsp_valid;
  wire       [31:0]   MmuPlugin_logic_accessBus_rsp_payload_data;
  reg                 MmuPlugin_logic_accessBus_rsp_payload_error;
  reg                 MmuPlugin_logic_accessBus_rsp_payload_redo;
  wire                MmuPlugin_logic_accessBus_rsp_payload_waitAny;
  reg        [0:0]    MmuPlugin_logic_satp_mode;
  reg        [19:0]   MmuPlugin_logic_satp_ppn;
  reg                 MmuPlugin_logic_status_mxr;
  reg                 MmuPlugin_logic_status_sum;
  reg                 MmuPlugin_logic_status_mprv;
  wire                BtbPlugin_logic_pcPort_valid;
  wire                BtbPlugin_logic_pcPort_payload_fault;
  wire       [31:0]   BtbPlugin_logic_pcPort_payload_pc;
  wire                PcPlugin_logic_harts_0_aggregator_sortedByPriority_5_laneValid;
  wire                BtbPlugin_logic_historyPort_valid;
  wire       [11:0]   BtbPlugin_logic_historyPort_payload_history;
  wire                BtbPlugin_logic_flushPort_valid;
  wire                BtbPlugin_logic_flushPort_payload_self;
  wire                FetchL1Plugin_logic_bus_cmd_valid;
  wire                FetchL1Plugin_logic_bus_cmd_ready;
  wire       [31:0]   FetchL1Plugin_logic_bus_cmd_payload_address;
  wire                FetchL1Plugin_logic_bus_cmd_payload_io;
  wire                FetchL1Plugin_logic_bus_rsp_valid;
  wire                FetchL1Plugin_logic_bus_rsp_ready;
  wire       [63:0]   FetchL1Plugin_logic_bus_rsp_payload_data;
  wire                FetchL1Plugin_logic_bus_rsp_payload_error;
  reg                 FetchL1Plugin_logic_trapPort_valid;
  reg                 FetchL1Plugin_logic_trapPort_payload_exception;
  wire       [31:0]   FetchL1Plugin_logic_trapPort_payload_tval;
  wire       [0:0]    decode_logic_trapPending;
  reg                 DecoderPlugin_logic_forgetPort_valid;
  reg        [31:0]   DecoderPlugin_logic_forgetPort_payload_pcOnLastSlice;
  wire       [0:0]    DispatchPlugin_logic_trapPendings;
  wire       [0:0]    execute_lane0_logic_trapPending;
  wire                early0_IntAluPlugin_logic_wb_valid;
  wire       [31:0]   early0_IntAluPlugin_logic_wb_payload;
  (* keep , syn_keep *) reg        [31:0]   early0_IntAluPlugin_logic_alu_bitwise /* synthesis syn_keep = 1 */ ;
  wire       [31:0]   early0_IntAluPlugin_logic_alu_result;
  wire                early0_BarrelShifterPlugin_logic_wb_valid;
  wire       [31:0]   early0_BarrelShifterPlugin_logic_wb_payload;
  wire       [4:0]    early0_BarrelShifterPlugin_logic_shift_amplitude;
  wire       [31:0]   early0_BarrelShifterPlugin_logic_shift_reversed;
  wire       [31:0]   early0_BarrelShifterPlugin_logic_shift_shifted;
  wire       [31:0]   early0_BarrelShifterPlugin_logic_shift_patched;
  wire                toplevel_execute_lane0_ctrls_3_upIsCancel;
  wire                toplevel_execute_lane0_ctrls_3_downIsCancel;
  wire                early0_BranchPlugin_logic_wb_valid;
  wire       [31:0]   early0_BranchPlugin_logic_wb_payload;
  wire                early0_BranchPlugin_logic_pcPort_valid;
  wire                early0_BranchPlugin_logic_pcPort_payload_fault;
  wire       [31:0]   early0_BranchPlugin_logic_pcPort_payload_pc;
  wire       [0:0]    early0_BranchPlugin_logic_pcPort_payload_laneAge;
  wire                PcPlugin_logic_harts_0_aggregator_sortedByPriority_3_laneValid;
  wire                early0_BranchPlugin_logic_historyPort_valid;
  wire       [11:0]   early0_BranchPlugin_logic_historyPort_payload_history;
  wire       [0:0]    early0_BranchPlugin_logic_historyPort_payload_age;
  wire                early0_BranchPlugin_logic_flushPort_valid;
  reg                 LsuPlugin_logic_trapPort_valid;
  reg                 LsuPlugin_logic_trapPort_payload_exception;
  wire       [31:0]   LsuPlugin_logic_trapPort_payload_tval;
  wire                LsuL1_lockPort_valid;
  wire       [31:0]   LsuL1_lockPort_address;
  reg                 LsuL1_ackUnlock;
  wire                early0_MulPlugin_logic_formatBus_valid;
  wire       [31:0]   early0_MulPlugin_logic_formatBus_payload;
  reg        [60:0]   _zz_toplevel_execute_ctrl3_down_early0_MulPlugin_logic_steps_0_adders_0_lane0;
  reg        [60:0]   _zz_toplevel_execute_ctrl3_down_early0_MulPlugin_logic_steps_0_adders_0_lane0_1;
  reg        [60:0]   _zz_toplevel_execute_ctrl3_down_early0_MulPlugin_logic_steps_0_adders_0_lane0_2;
  reg        [2:0]    _zz_toplevel_execute_ctrl3_down_early0_MulPlugin_logic_steps_0_adders_1_lane0;
  reg        [2:0]    _zz_toplevel_execute_ctrl3_down_early0_MulPlugin_logic_steps_0_adders_1_lane0_1;
  reg        [2:0]    _zz_toplevel_execute_ctrl3_down_early0_MulPlugin_logic_steps_0_adders_1_lane0_2;
  wire                toplevel_execute_lane0_ctrls_4_upIsCancel;
  wire                toplevel_execute_lane0_ctrls_4_downIsCancel;
  reg        [65:0]   _zz_toplevel_execute_ctrl4_down_early0_MulPlugin_logic_steps_1_adders_0_lane0;
  reg        [65:0]   _zz_toplevel_execute_ctrl4_down_early0_MulPlugin_logic_steps_1_adders_0_lane0_1;
  reg                 early0_MulPlugin_logic_writeback_buffer_valid;
  wire                when_MulPlugin_l195;
  reg        [31:0]   early0_MulPlugin_logic_writeback_buffer_data;
  wire                early0_DivPlugin_logic_formatBus_valid;
  wire       [31:0]   early0_DivPlugin_logic_formatBus_payload;
  reg                 early0_DivPlugin_logic_processing_divRevertResult;
  reg                 early0_DivPlugin_logic_processing_cmdSent;
  wire                early0_DivPlugin_logic_processing_div_io_cmd_fire;
  wire                early0_DivPlugin_logic_processing_request;
  wire       [31:0]   early0_DivPlugin_logic_processing_a;
  wire       [31:0]   early0_DivPlugin_logic_processing_b;
  reg        [31:0]   early0_DivPlugin_logic_processing_a_delay_1;
  reg        [31:0]   early0_DivPlugin_logic_processing_b_delay_1;
  reg                 early0_DivPlugin_logic_processing_relaxer_hadRequest;
  wire                when_DivPlugin_l118;
  reg                 early0_DivPlugin_logic_processing_unscheduleRequest;
  wire                early0_DivPlugin_logic_processing_freeze;
  wire       [31:0]   early0_DivPlugin_logic_processing_selected;
  wire       [31:0]   _zz_toplevel_execute_ctrl2_down_DivPlugin_DIV_RESULT_lane0;
  wire                CsrAccessPlugin_logic_wbWi_valid;
  wire       [31:0]   CsrAccessPlugin_logic_wbWi_payload;
  reg                 CsrAccessPlugin_logic_flushPort_valid;
  reg                 TrapPlugin_logic_fetchL1Invalidate_0_cmd_valid;
  reg                 TrapPlugin_logic_fetchL1Invalidate_0_cmd_ready;
  reg                 TrapPlugin_logic_lsuL1Invalidate_0_cmd_valid;
  wire                TrapPlugin_logic_lsuL1Invalidate_0_cmd_ready;
  reg                 early0_EnvPlugin_logic_trapPort_valid;
  reg                 early0_EnvPlugin_logic_trapPort_payload_exception;
  wire       [31:0]   early0_EnvPlugin_logic_trapPort_payload_tval;
  reg        [3:0]    early0_EnvPlugin_logic_trapPort_payload_code;
  reg        [2:0]    early0_EnvPlugin_logic_trapPort_payload_arg;
  wire       [0:0]    early0_EnvPlugin_logic_trapPort_payload_laneAge;
  reg                 early0_EnvPlugin_logic_flushPort_valid;
  wire                late0_IntAluPlugin_logic_wb_valid;
  wire       [31:0]   late0_IntAluPlugin_logic_wb_payload;
  (* keep , syn_keep *) reg        [31:0]   late0_IntAluPlugin_logic_alu_bitwise /* synthesis syn_keep = 1 */ ;
  wire       [31:0]   late0_IntAluPlugin_logic_alu_result;
  wire                late0_BarrelShifterPlugin_logic_wb_valid;
  wire       [31:0]   late0_BarrelShifterPlugin_logic_wb_payload;
  wire       [4:0]    late0_BarrelShifterPlugin_logic_shift_amplitude;
  wire       [31:0]   late0_BarrelShifterPlugin_logic_shift_reversed;
  wire       [31:0]   late0_BarrelShifterPlugin_logic_shift_shifted;
  wire       [31:0]   late0_BarrelShifterPlugin_logic_shift_patched;
  wire                late0_BranchPlugin_logic_wb_valid;
  wire       [31:0]   late0_BranchPlugin_logic_wb_payload;
  wire                late0_BranchPlugin_logic_pcPort_valid;
  wire                late0_BranchPlugin_logic_pcPort_payload_fault;
  wire       [31:0]   late0_BranchPlugin_logic_pcPort_payload_pc;
  wire       [0:0]    late0_BranchPlugin_logic_pcPort_payload_laneAge;
  wire                PcPlugin_logic_harts_0_aggregator_sortedByPriority_1_laneValid;
  wire                late0_BranchPlugin_logic_historyPort_valid;
  wire       [11:0]   late0_BranchPlugin_logic_historyPort_payload_history;
  wire       [0:0]    late0_BranchPlugin_logic_historyPort_payload_age;
  wire                late0_BranchPlugin_logic_flushPort_valid;
  wire       [0:0]    execute_lane1_logic_trapPending;
  wire                early1_IntAluPlugin_logic_wb_valid;
  wire       [31:0]   early1_IntAluPlugin_logic_wb_payload;
  (* keep , syn_keep *) reg        [31:0]   early1_IntAluPlugin_logic_alu_bitwise /* synthesis syn_keep = 1 */ ;
  wire       [31:0]   early1_IntAluPlugin_logic_alu_result;
  wire                early1_BarrelShifterPlugin_logic_wb_valid;
  wire       [31:0]   early1_BarrelShifterPlugin_logic_wb_payload;
  wire       [4:0]    early1_BarrelShifterPlugin_logic_shift_amplitude;
  wire       [31:0]   early1_BarrelShifterPlugin_logic_shift_reversed;
  wire       [31:0]   early1_BarrelShifterPlugin_logic_shift_shifted;
  wire       [31:0]   early1_BarrelShifterPlugin_logic_shift_patched;
  wire                toplevel_execute_lane1_ctrls_3_upIsCancel;
  wire                toplevel_execute_lane1_ctrls_3_downIsCancel;
  wire                early1_BranchPlugin_logic_wb_valid;
  wire       [31:0]   early1_BranchPlugin_logic_wb_payload;
  wire                early1_BranchPlugin_logic_pcPort_valid;
  wire                early1_BranchPlugin_logic_pcPort_payload_fault;
  wire       [31:0]   early1_BranchPlugin_logic_pcPort_payload_pc;
  wire       [0:0]    early1_BranchPlugin_logic_pcPort_payload_laneAge;
  wire                PcPlugin_logic_harts_0_aggregator_sortedByPriority_4_laneValid;
  wire                early1_BranchPlugin_logic_historyPort_valid;
  wire       [11:0]   early1_BranchPlugin_logic_historyPort_payload_history;
  wire       [0:0]    early1_BranchPlugin_logic_historyPort_payload_age;
  wire                early1_BranchPlugin_logic_flushPort_valid;
  wire                late1_IntAluPlugin_logic_wb_valid;
  wire       [31:0]   late1_IntAluPlugin_logic_wb_payload;
  wire                toplevel_execute_lane1_ctrls_4_upIsCancel;
  wire                toplevel_execute_lane1_ctrls_4_downIsCancel;
  (* keep , syn_keep *) reg        [31:0]   late1_IntAluPlugin_logic_alu_bitwise /* synthesis syn_keep = 1 */ ;
  wire       [31:0]   late1_IntAluPlugin_logic_alu_result;
  wire                late1_BarrelShifterPlugin_logic_wb_valid;
  wire       [31:0]   late1_BarrelShifterPlugin_logic_wb_payload;
  wire       [4:0]    late1_BarrelShifterPlugin_logic_shift_amplitude;
  wire       [31:0]   late1_BarrelShifterPlugin_logic_shift_reversed;
  wire       [31:0]   late1_BarrelShifterPlugin_logic_shift_shifted;
  wire       [31:0]   late1_BarrelShifterPlugin_logic_shift_patched;
  wire                late1_BranchPlugin_logic_wb_valid;
  wire       [31:0]   late1_BranchPlugin_logic_wb_payload;
  wire                late1_BranchPlugin_logic_pcPort_valid;
  wire                late1_BranchPlugin_logic_pcPort_payload_fault;
  wire       [31:0]   late1_BranchPlugin_logic_pcPort_payload_pc;
  wire       [0:0]    late1_BranchPlugin_logic_pcPort_payload_laneAge;
  wire                PcPlugin_logic_harts_0_aggregator_sortedByPriority_2_laneValid;
  wire                late1_BranchPlugin_logic_historyPort_valid;
  wire       [11:0]   late1_BranchPlugin_logic_historyPort_payload_history;
  wire       [0:0]    late1_BranchPlugin_logic_historyPort_payload_age;
  wire                late1_BranchPlugin_logic_flushPort_valid;
  wire                WhiteboxerPlugin_logic_fetch_fire;
  wire       [31:0]   PrivilegedPlugin_api_lsuTriggerBus_virtual;
  wire       [1:0]    PrivilegedPlugin_api_lsuTriggerBus_size;
  wire                PrivilegedPlugin_api_harts_0_allowInterrupts;
  wire                PrivilegedPlugin_api_harts_0_allowException;
  wire                PrivilegedPlugin_api_harts_0_allowEbreakException;
  wire                PrivilegedPlugin_api_harts_0_fpuEnable;
  reg        [31:0]   early0_BranchPlugin_pcCalc_target_a;
  reg        [31:0]   early0_BranchPlugin_pcCalc_target_b;
  wire       [1:0]    early0_BranchPlugin_pcCalc_slices;
  reg        [31:0]   early1_BranchPlugin_pcCalc_target_a;
  reg        [31:0]   early1_BranchPlugin_pcCalc_target_b;
  wire       [1:0]    early1_BranchPlugin_pcCalc_slices;
  wire       [3:0]    AlignerPlugin_logic_maskGen_frontMasks_0;
  wire       [3:0]    AlignerPlugin_logic_maskGen_frontMasks_1;
  wire       [3:0]    AlignerPlugin_logic_maskGen_frontMasks_2;
  wire       [3:0]    AlignerPlugin_logic_maskGen_frontMasks_3;
  wire       [3:0]    AlignerPlugin_logic_maskGen_backMasks_0;
  wire       [3:0]    AlignerPlugin_logic_maskGen_backMasks_1;
  wire       [3:0]    AlignerPlugin_logic_maskGen_backMasks_2;
  wire       [3:0]    AlignerPlugin_logic_maskGen_backMasks_3;
  wire       [15:0]   AlignerPlugin_logic_slices_data_0;
  wire       [15:0]   AlignerPlugin_logic_slices_data_1;
  wire       [15:0]   AlignerPlugin_logic_slices_data_2;
  wire       [15:0]   AlignerPlugin_logic_slices_data_3;
  wire       [15:0]   AlignerPlugin_logic_slices_data_4;
  wire       [15:0]   AlignerPlugin_logic_slices_data_5;
  wire       [15:0]   AlignerPlugin_logic_slices_data_6;
  wire       [15:0]   AlignerPlugin_logic_slices_data_7;
  wire       [7:0]    AlignerPlugin_logic_slices_mask;
  wire       [7:0]    AlignerPlugin_logic_slices_last;
  wire       [31:0]   AlignerPlugin_logic_slicesInstructions_0;
  wire       [31:0]   AlignerPlugin_logic_slicesInstructions_1;
  wire       [31:0]   AlignerPlugin_logic_slicesInstructions_2;
  wire       [31:0]   AlignerPlugin_logic_slicesInstructions_3;
  wire       [31:0]   AlignerPlugin_logic_slicesInstructions_4;
  wire       [31:0]   AlignerPlugin_logic_slicesInstructions_5;
  wire       [31:0]   AlignerPlugin_logic_slicesInstructions_6;
  wire       [31:0]   AlignerPlugin_logic_slicesInstructions_7;
  reg        [7:0]    AlignerPlugin_logic_scanners_0_usageMask;
  wire                AlignerPlugin_logic_scanners_0_checker_0_required;
  wire                AlignerPlugin_logic_scanners_0_checker_0_last;
  wire                AlignerPlugin_logic_scanners_0_checker_0_redo;
  wire                AlignerPlugin_logic_scanners_0_checker_0_present;
  wire                AlignerPlugin_logic_scanners_0_checker_0_valid;
  wire                AlignerPlugin_logic_scanners_0_checker_1_required;
  wire                AlignerPlugin_logic_scanners_0_checker_1_last;
  wire                AlignerPlugin_logic_scanners_0_checker_1_redo;
  wire                AlignerPlugin_logic_scanners_0_checker_1_present;
  wire                AlignerPlugin_logic_scanners_0_checker_1_valid;
  wire                AlignerPlugin_logic_scanners_0_redo;
  wire                AlignerPlugin_logic_scanners_0_valid;
  reg        [7:0]    AlignerPlugin_logic_scanners_1_usageMask;
  wire                AlignerPlugin_logic_scanners_1_checker_0_required;
  wire                AlignerPlugin_logic_scanners_1_checker_0_last;
  wire                AlignerPlugin_logic_scanners_1_checker_0_redo;
  wire                AlignerPlugin_logic_scanners_1_checker_0_present;
  wire                AlignerPlugin_logic_scanners_1_checker_0_valid;
  wire                AlignerPlugin_logic_scanners_1_checker_1_required;
  wire                AlignerPlugin_logic_scanners_1_checker_1_last;
  wire                AlignerPlugin_logic_scanners_1_checker_1_redo;
  wire                AlignerPlugin_logic_scanners_1_checker_1_present;
  wire                AlignerPlugin_logic_scanners_1_checker_1_valid;
  wire                AlignerPlugin_logic_scanners_1_redo;
  wire                AlignerPlugin_logic_scanners_1_valid;
  reg        [7:0]    AlignerPlugin_logic_scanners_2_usageMask;
  wire                AlignerPlugin_logic_scanners_2_checker_0_required;
  wire                AlignerPlugin_logic_scanners_2_checker_0_last;
  wire                AlignerPlugin_logic_scanners_2_checker_0_redo;
  wire                AlignerPlugin_logic_scanners_2_checker_0_present;
  wire                AlignerPlugin_logic_scanners_2_checker_0_valid;
  wire                AlignerPlugin_logic_scanners_2_checker_1_required;
  wire                AlignerPlugin_logic_scanners_2_checker_1_last;
  wire                AlignerPlugin_logic_scanners_2_checker_1_redo;
  wire                AlignerPlugin_logic_scanners_2_checker_1_present;
  wire                AlignerPlugin_logic_scanners_2_checker_1_valid;
  wire                AlignerPlugin_logic_scanners_2_redo;
  wire                AlignerPlugin_logic_scanners_2_valid;
  reg        [7:0]    AlignerPlugin_logic_scanners_3_usageMask;
  wire                AlignerPlugin_logic_scanners_3_checker_0_required;
  wire                AlignerPlugin_logic_scanners_3_checker_0_last;
  wire                AlignerPlugin_logic_scanners_3_checker_0_redo;
  wire                AlignerPlugin_logic_scanners_3_checker_0_present;
  wire                AlignerPlugin_logic_scanners_3_checker_0_valid;
  wire                AlignerPlugin_logic_scanners_3_checker_1_required;
  wire                AlignerPlugin_logic_scanners_3_checker_1_last;
  wire                AlignerPlugin_logic_scanners_3_checker_1_redo;
  wire                AlignerPlugin_logic_scanners_3_checker_1_present;
  wire                AlignerPlugin_logic_scanners_3_checker_1_valid;
  wire                AlignerPlugin_logic_scanners_3_redo;
  wire                AlignerPlugin_logic_scanners_3_valid;
  reg        [7:0]    AlignerPlugin_logic_scanners_4_usageMask;
  wire                AlignerPlugin_logic_scanners_4_checker_0_required;
  wire                AlignerPlugin_logic_scanners_4_checker_0_last;
  wire                AlignerPlugin_logic_scanners_4_checker_0_redo;
  wire                AlignerPlugin_logic_scanners_4_checker_0_present;
  wire                AlignerPlugin_logic_scanners_4_checker_0_valid;
  wire                AlignerPlugin_logic_scanners_4_checker_1_required;
  wire                AlignerPlugin_logic_scanners_4_checker_1_last;
  wire                AlignerPlugin_logic_scanners_4_checker_1_redo;
  wire                AlignerPlugin_logic_scanners_4_checker_1_present;
  wire                AlignerPlugin_logic_scanners_4_checker_1_valid;
  wire                AlignerPlugin_logic_scanners_4_redo;
  wire                AlignerPlugin_logic_scanners_4_valid;
  reg        [7:0]    AlignerPlugin_logic_scanners_5_usageMask;
  wire                AlignerPlugin_logic_scanners_5_checker_0_required;
  wire                AlignerPlugin_logic_scanners_5_checker_0_last;
  wire                AlignerPlugin_logic_scanners_5_checker_0_redo;
  wire                AlignerPlugin_logic_scanners_5_checker_0_present;
  wire                AlignerPlugin_logic_scanners_5_checker_0_valid;
  wire                AlignerPlugin_logic_scanners_5_checker_1_required;
  wire                AlignerPlugin_logic_scanners_5_checker_1_last;
  wire                AlignerPlugin_logic_scanners_5_checker_1_redo;
  wire                AlignerPlugin_logic_scanners_5_checker_1_present;
  wire                AlignerPlugin_logic_scanners_5_checker_1_valid;
  wire                AlignerPlugin_logic_scanners_5_redo;
  wire                AlignerPlugin_logic_scanners_5_valid;
  reg        [7:0]    AlignerPlugin_logic_scanners_6_usageMask;
  wire                AlignerPlugin_logic_scanners_6_checker_0_required;
  wire                AlignerPlugin_logic_scanners_6_checker_0_last;
  wire                AlignerPlugin_logic_scanners_6_checker_0_redo;
  wire                AlignerPlugin_logic_scanners_6_checker_0_present;
  wire                AlignerPlugin_logic_scanners_6_checker_0_valid;
  wire                AlignerPlugin_logic_scanners_6_checker_1_required;
  wire                AlignerPlugin_logic_scanners_6_checker_1_last;
  wire                AlignerPlugin_logic_scanners_6_checker_1_redo;
  wire                AlignerPlugin_logic_scanners_6_checker_1_present;
  wire                AlignerPlugin_logic_scanners_6_checker_1_valid;
  wire                AlignerPlugin_logic_scanners_6_redo;
  wire                AlignerPlugin_logic_scanners_6_valid;
  reg        [7:0]    AlignerPlugin_logic_scanners_7_usageMask;
  wire                AlignerPlugin_logic_scanners_7_checker_0_required;
  wire                AlignerPlugin_logic_scanners_7_checker_0_last;
  wire                AlignerPlugin_logic_scanners_7_checker_0_redo;
  wire                AlignerPlugin_logic_scanners_7_checker_0_present;
  wire                AlignerPlugin_logic_scanners_7_checker_0_valid;
  wire                AlignerPlugin_logic_scanners_7_checker_1_required;
  wire                AlignerPlugin_logic_scanners_7_checker_1_last;
  wire                AlignerPlugin_logic_scanners_7_checker_1_redo;
  wire                AlignerPlugin_logic_scanners_7_checker_1_present;
  wire                AlignerPlugin_logic_scanners_7_checker_1_valid;
  wire                AlignerPlugin_logic_scanners_7_redo;
  wire                AlignerPlugin_logic_scanners_7_valid;
  wire       [7:0]    AlignerPlugin_logic_usedMask_0;
  wire       [7:0]    AlignerPlugin_logic_usedMask_1;
  wire       [7:0]    AlignerPlugin_logic_usedMask_2;
  wire                AlignerPlugin_logic_extractors_0_first;
  wire       [7:0]    AlignerPlugin_logic_extractors_0_usableMask;
  wire       [7:0]    _zz_AlignerPlugin_logic_extractors_0_usableMask_bools_0;
  wire                AlignerPlugin_logic_extractors_0_usableMask_bools_0;
  wire                AlignerPlugin_logic_extractors_0_usableMask_bools_1;
  wire                AlignerPlugin_logic_extractors_0_usableMask_bools_2;
  wire                AlignerPlugin_logic_extractors_0_usableMask_bools_3;
  wire                AlignerPlugin_logic_extractors_0_usableMask_bools_4;
  wire                AlignerPlugin_logic_extractors_0_usableMask_bools_5;
  wire                AlignerPlugin_logic_extractors_0_usableMask_bools_6;
  wire                AlignerPlugin_logic_extractors_0_usableMask_bools_7;
  reg        [7:0]    _zz_AlignerPlugin_logic_extractors_0_slicesOh;
  wire                AlignerPlugin_logic_extractors_0_usableMask_range_0_to_1;
  wire                AlignerPlugin_logic_extractors_0_usableMask_range_0_to_2;
  wire                AlignerPlugin_logic_extractors_0_usableMask_range_0_to_3;
  wire                AlignerPlugin_logic_extractors_0_usableMask_range_4_to_5;
  wire                AlignerPlugin_logic_extractors_0_usableMask_range_4_to_6;
  wire       [7:0]    AlignerPlugin_logic_extractors_0_slicesOh;
  wire                _zz_AlignerPlugin_logic_extractors_0_redo;
  wire                _zz_AlignerPlugin_logic_extractors_0_redo_1;
  wire                _zz_AlignerPlugin_logic_extractors_0_redo_2;
  wire                _zz_AlignerPlugin_logic_extractors_0_redo_3;
  wire                _zz_AlignerPlugin_logic_extractors_0_redo_4;
  wire                _zz_AlignerPlugin_logic_extractors_0_redo_5;
  wire                _zz_AlignerPlugin_logic_extractors_0_redo_6;
  wire                _zz_AlignerPlugin_logic_extractors_0_redo_7;
  reg                 AlignerPlugin_logic_extractors_0_redo;
  wire       [1:0]    AlignerPlugin_logic_extractors_0_localMask;
  wire       [7:0]    AlignerPlugin_logic_extractors_0_usageMask;
  reg                 AlignerPlugin_logic_extractors_0_valid;
  reg        [31:0]   AlignerPlugin_logic_extractors_0_ctx_pc;
  wire       [31:0]   AlignerPlugin_logic_extractors_0_ctx_instruction;
  wire       [9:0]    AlignerPlugin_logic_extractors_0_ctx_hm_Fetch_ID;
  wire       [1:0]    AlignerPlugin_logic_extractors_0_ctx_hm_GSharePlugin_GSHARE_COUNTER_0;
  wire       [1:0]    AlignerPlugin_logic_extractors_0_ctx_hm_GSharePlugin_GSHARE_COUNTER_1;
  wire       [1:0]    AlignerPlugin_logic_extractors_0_ctx_hm_GSharePlugin_GSHARE_COUNTER_2;
  wire       [1:0]    AlignerPlugin_logic_extractors_0_ctx_hm_GSharePlugin_GSHARE_COUNTER_3;
  wire       [11:0]   AlignerPlugin_logic_extractors_0_ctx_hm_Prediction_BRANCH_HISTORY;
  wire       [3:0]    AlignerPlugin_logic_extractors_0_ctx_hm_Prediction_WORD_SLICES_BRANCH;
  wire       [3:0]    AlignerPlugin_logic_extractors_0_ctx_hm_Prediction_WORD_SLICES_TAKEN;
  wire       [31:0]   AlignerPlugin_logic_extractors_0_ctx_hm_Prediction_WORD_JUMP_PC;
  wire                AlignerPlugin_logic_extractors_0_ctx_hm_Prediction_WORD_JUMPED;
  wire       [1:0]    AlignerPlugin_logic_extractors_0_ctx_hm_Prediction_WORD_JUMP_SLICE;
  wire                AlignerPlugin_logic_extractors_0_ctx_trap;
  wire                when_AlignerPlugin_l163;
  wire                AlignerPlugin_logic_extractors_1_first;
  wire       [6:0]    AlignerPlugin_logic_extractors_1_usableMask;
  wire       [6:0]    _zz_AlignerPlugin_logic_extractors_1_usableMask_bools_0;
  wire                AlignerPlugin_logic_extractors_1_usableMask_bools_0;
  wire                AlignerPlugin_logic_extractors_1_usableMask_bools_1;
  wire                AlignerPlugin_logic_extractors_1_usableMask_bools_2;
  wire                AlignerPlugin_logic_extractors_1_usableMask_bools_3;
  wire                AlignerPlugin_logic_extractors_1_usableMask_bools_4;
  wire                AlignerPlugin_logic_extractors_1_usableMask_bools_5;
  wire                AlignerPlugin_logic_extractors_1_usableMask_bools_6;
  reg        [6:0]    _zz_AlignerPlugin_logic_extractors_1_slicesOh;
  wire                AlignerPlugin_logic_extractors_1_usableMask_range_0_to_1;
  wire                AlignerPlugin_logic_extractors_1_usableMask_range_0_to_2;
  wire                AlignerPlugin_logic_extractors_1_usableMask_range_0_to_3;
  wire                AlignerPlugin_logic_extractors_1_usableMask_range_4_to_5;
  wire       [6:0]    AlignerPlugin_logic_extractors_1_slicesOh;
  wire                _zz_AlignerPlugin_logic_extractors_1_redo;
  wire                _zz_AlignerPlugin_logic_extractors_1_redo_1;
  wire                _zz_AlignerPlugin_logic_extractors_1_redo_2;
  wire                _zz_AlignerPlugin_logic_extractors_1_redo_3;
  wire                _zz_AlignerPlugin_logic_extractors_1_redo_4;
  wire                _zz_AlignerPlugin_logic_extractors_1_redo_5;
  wire                _zz_AlignerPlugin_logic_extractors_1_redo_6;
  reg                 AlignerPlugin_logic_extractors_1_redo;
  wire       [1:0]    AlignerPlugin_logic_extractors_1_localMask;
  wire       [7:0]    AlignerPlugin_logic_extractors_1_usageMask;
  reg                 AlignerPlugin_logic_extractors_1_valid;
  reg        [31:0]   AlignerPlugin_logic_extractors_1_ctx_pc;
  wire       [31:0]   AlignerPlugin_logic_extractors_1_ctx_instruction;
  wire       [9:0]    AlignerPlugin_logic_extractors_1_ctx_hm_Fetch_ID;
  wire       [1:0]    AlignerPlugin_logic_extractors_1_ctx_hm_GSharePlugin_GSHARE_COUNTER_0;
  wire       [1:0]    AlignerPlugin_logic_extractors_1_ctx_hm_GSharePlugin_GSHARE_COUNTER_1;
  wire       [1:0]    AlignerPlugin_logic_extractors_1_ctx_hm_GSharePlugin_GSHARE_COUNTER_2;
  wire       [1:0]    AlignerPlugin_logic_extractors_1_ctx_hm_GSharePlugin_GSHARE_COUNTER_3;
  wire       [11:0]   AlignerPlugin_logic_extractors_1_ctx_hm_Prediction_BRANCH_HISTORY;
  wire       [3:0]    AlignerPlugin_logic_extractors_1_ctx_hm_Prediction_WORD_SLICES_BRANCH;
  wire       [3:0]    AlignerPlugin_logic_extractors_1_ctx_hm_Prediction_WORD_SLICES_TAKEN;
  wire       [31:0]   AlignerPlugin_logic_extractors_1_ctx_hm_Prediction_WORD_JUMP_PC;
  wire                AlignerPlugin_logic_extractors_1_ctx_hm_Prediction_WORD_JUMPED;
  wire       [1:0]    AlignerPlugin_logic_extractors_1_ctx_hm_Prediction_WORD_JUMP_SLICE;
  wire                AlignerPlugin_logic_extractors_1_ctx_trap;
  wire                when_AlignerPlugin_l163_1;
  reg        [9:0]    AlignerPlugin_logic_feeder_harts_0_dopId;
  wire                when_AlignerPlugin_l173;
  wire                AlignerPlugin_logic_feeder_lanes_0_valid;
  wire                AlignerPlugin_logic_feeder_lanes_0_isRvc;
  reg        [31:0]   AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst;
  reg                 AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_illegal;
  wire       [4:0]    _zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst;
  wire       [4:0]    _zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_1;
  wire       [11:0]   _zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_2;
  wire       [11:0]   _zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_3;
  wire                _zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_4;
  reg        [11:0]   _zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_5;
  wire                _zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_6;
  reg        [9:0]    _zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_7;
  wire       [20:0]   _zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_8;
  wire                _zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_9;
  reg        [14:0]   _zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_10;
  wire                _zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_11;
  reg        [2:0]    _zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_12;
  wire                _zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_13;
  reg        [9:0]    _zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_14;
  wire       [20:0]   _zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_15;
  wire                _zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_16;
  reg        [4:0]    _zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_17;
  wire       [12:0]   _zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_18;
  wire       [4:0]    _zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_19;
  wire       [4:0]    _zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_20;
  wire       [4:0]    _zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_21;
  wire       [4:0]    switch_Rvc_l52;
  wire                when_Rvc_l56;
  wire                when_Rvc_l77;
  wire       [31:0]   _zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_22;
  wire                when_Rvc_l98;
  wire                when_Rvc_l111;
  wire       [1:0]    _zz_toplevel_decode_ctrls_0_up_Decode_INSTRUCTION_SLICE_COUNT_0;
  wire       [1:0]    _zz_toplevel_decode_ctrls_0_up_Decode_INSTRUCTION_SLICE_COUNT_0_1;
  wire                _zz_toplevel_decode_ctrls_0_up_Decode_INSTRUCTION_SLICE_COUNT_0_2;
  reg        [1:0]    _zz_toplevel_decode_ctrls_0_up_Decode_INSTRUCTION_SLICE_COUNT_0_3;
  wire       [1:0]    _zz_toplevel_decode_ctrls_0_up_Decode_INSTRUCTION_SLICE_COUNT_0_4;
  wire                _zz_toplevel_decode_ctrls_0_up_Decode_INSTRUCTION_SLICE_COUNT_0_5;
  wire       [1:0]    AlignerPlugin_logic_feeder_lanes_0_onBtb_pcLastSlice;
  wire                AlignerPlugin_logic_feeder_lanes_0_onBtb_didPrediction;
  wire                AlignerPlugin_logic_feeder_lanes_1_valid;
  wire                AlignerPlugin_logic_feeder_lanes_1_isRvc;
  reg        [31:0]   AlignerPlugin_logic_feeder_lanes_1_withRvc_dec_inst;
  reg                 AlignerPlugin_logic_feeder_lanes_1_withRvc_dec_illegal;
  wire       [4:0]    _zz_AlignerPlugin_logic_feeder_lanes_1_withRvc_dec_inst;
  wire       [4:0]    _zz_AlignerPlugin_logic_feeder_lanes_1_withRvc_dec_inst_1;
  wire       [11:0]   _zz_AlignerPlugin_logic_feeder_lanes_1_withRvc_dec_inst_2;
  wire       [11:0]   _zz_AlignerPlugin_logic_feeder_lanes_1_withRvc_dec_inst_3;
  wire                _zz_AlignerPlugin_logic_feeder_lanes_1_withRvc_dec_inst_4;
  reg        [11:0]   _zz_AlignerPlugin_logic_feeder_lanes_1_withRvc_dec_inst_5;
  wire                _zz_AlignerPlugin_logic_feeder_lanes_1_withRvc_dec_inst_6;
  reg        [9:0]    _zz_AlignerPlugin_logic_feeder_lanes_1_withRvc_dec_inst_7;
  wire       [20:0]   _zz_AlignerPlugin_logic_feeder_lanes_1_withRvc_dec_inst_8;
  wire                _zz_AlignerPlugin_logic_feeder_lanes_1_withRvc_dec_inst_9;
  reg        [14:0]   _zz_AlignerPlugin_logic_feeder_lanes_1_withRvc_dec_inst_10;
  wire                _zz_AlignerPlugin_logic_feeder_lanes_1_withRvc_dec_inst_11;
  reg        [2:0]    _zz_AlignerPlugin_logic_feeder_lanes_1_withRvc_dec_inst_12;
  wire                _zz_AlignerPlugin_logic_feeder_lanes_1_withRvc_dec_inst_13;
  reg        [9:0]    _zz_AlignerPlugin_logic_feeder_lanes_1_withRvc_dec_inst_14;
  wire       [20:0]   _zz_AlignerPlugin_logic_feeder_lanes_1_withRvc_dec_inst_15;
  wire                _zz_AlignerPlugin_logic_feeder_lanes_1_withRvc_dec_inst_16;
  reg        [4:0]    _zz_AlignerPlugin_logic_feeder_lanes_1_withRvc_dec_inst_17;
  wire       [12:0]   _zz_AlignerPlugin_logic_feeder_lanes_1_withRvc_dec_inst_18;
  wire       [4:0]    _zz_AlignerPlugin_logic_feeder_lanes_1_withRvc_dec_inst_19;
  wire       [4:0]    _zz_AlignerPlugin_logic_feeder_lanes_1_withRvc_dec_inst_20;
  wire       [4:0]    _zz_AlignerPlugin_logic_feeder_lanes_1_withRvc_dec_inst_21;
  wire       [4:0]    switch_Rvc_l52_1;
  wire                when_Rvc_l56_1;
  wire                when_Rvc_l77_1;
  wire       [31:0]   _zz_AlignerPlugin_logic_feeder_lanes_1_withRvc_dec_inst_22;
  wire                when_Rvc_l98_1;
  wire                when_Rvc_l111_1;
  wire       [1:0]    _zz_toplevel_decode_ctrls_0_up_Decode_INSTRUCTION_SLICE_COUNT_1;
  wire       [1:0]    _zz_toplevel_decode_ctrls_0_up_Decode_INSTRUCTION_SLICE_COUNT_1_1;
  wire                _zz_toplevel_decode_ctrls_0_up_Decode_INSTRUCTION_SLICE_COUNT_1_2;
  reg        [1:0]    _zz_toplevel_decode_ctrls_0_up_Decode_INSTRUCTION_SLICE_COUNT_1_3;
  wire       [1:0]    _zz_toplevel_decode_ctrls_0_up_Decode_INSTRUCTION_SLICE_COUNT_1_4;
  wire                _zz_toplevel_decode_ctrls_0_up_Decode_INSTRUCTION_SLICE_COUNT_1_5;
  wire       [1:0]    AlignerPlugin_logic_feeder_lanes_1_onBtb_pcLastSlice;
  wire                AlignerPlugin_logic_feeder_lanes_1_onBtb_didPrediction;
  reg        [63:0]   AlignerPlugin_logic_buffer_data;
  reg        [3:0]    AlignerPlugin_logic_buffer_mask;
  reg        [3:0]    AlignerPlugin_logic_buffer_last;
  reg        [31:0]   AlignerPlugin_logic_buffer_pc;
  reg                 AlignerPlugin_logic_buffer_trap;
  reg        [9:0]    AlignerPlugin_logic_buffer_hm_Fetch_ID;
  reg        [1:0]    AlignerPlugin_logic_buffer_hm_GSharePlugin_GSHARE_COUNTER_0;
  reg        [1:0]    AlignerPlugin_logic_buffer_hm_GSharePlugin_GSHARE_COUNTER_1;
  reg        [1:0]    AlignerPlugin_logic_buffer_hm_GSharePlugin_GSHARE_COUNTER_2;
  reg        [1:0]    AlignerPlugin_logic_buffer_hm_GSharePlugin_GSHARE_COUNTER_3;
  reg        [11:0]   AlignerPlugin_logic_buffer_hm_Prediction_BRANCH_HISTORY;
  reg        [3:0]    AlignerPlugin_logic_buffer_hm_Prediction_WORD_SLICES_BRANCH;
  reg        [3:0]    AlignerPlugin_logic_buffer_hm_Prediction_WORD_SLICES_TAKEN;
  reg        [31:0]   AlignerPlugin_logic_buffer_hm_Prediction_WORD_JUMP_PC;
  reg                 AlignerPlugin_logic_buffer_hm_Prediction_WORD_JUMPED;
  reg        [1:0]    AlignerPlugin_logic_buffer_hm_Prediction_WORD_JUMP_SLICE;
  wire       [127:0]  _zz_AlignerPlugin_logic_slices_data_0;
  wire                when_AlignerPlugin_l243;
  wire                when_AlignerPlugin_l244;
  wire                when_AlignerPlugin_l244_1;
  wire                AlignerPlugin_logic_buffer_downFire;
  wire       [7:0]    AlignerPlugin_logic_buffer_usedMask;
  wire                AlignerPlugin_logic_buffer_haltUp;
  wire                when_AlignerPlugin_l259;
  reg        [3:0]    CsrAccessPlugin_bus_decode_trapCode;
  wire                CsrAccessPlugin_bus_read_valid;
  wire                CsrAccessPlugin_bus_read_moving;
  wire       [11:0]   CsrAccessPlugin_bus_read_address;
  reg                 CsrAccessPlugin_bus_read_halt;
  reg        [31:0]   CsrAccessPlugin_bus_read_toWriteBits;
  wire       [31:0]   CsrAccessPlugin_bus_read_data;
  wire                CsrAccessPlugin_bus_write_valid;
  wire                CsrAccessPlugin_bus_write_moving;
  reg                 CsrAccessPlugin_bus_write_halt;
  reg        [31:0]   CsrAccessPlugin_bus_write_bits;
  wire       [11:0]   CsrAccessPlugin_bus_write_address;
  reg        [3:0]    FetchL1Plugin_logic_trapPort_payload_code;
  reg        [2:0]    FetchL1Plugin_logic_trapPort_payload_arg;
  reg                 FetchL1Plugin_logic_banks_0_write_valid;
  reg        [8:0]    FetchL1Plugin_logic_banks_0_write_payload_address;
  reg        [63:0]   FetchL1Plugin_logic_banks_0_write_payload_data;
  wire                FetchL1Plugin_logic_banks_0_read_cmd_valid;
  wire       [8:0]    FetchL1Plugin_logic_banks_0_read_cmd_payload;
  (* keep , syn_keep *) wire       [63:0]   FetchL1Plugin_logic_banks_0_read_rsp /* synthesis syn_keep = 1 */ ;
  reg                 FetchL1Plugin_logic_banks_1_write_valid;
  reg        [8:0]    FetchL1Plugin_logic_banks_1_write_payload_address;
  reg        [63:0]   FetchL1Plugin_logic_banks_1_write_payload_data;
  wire                FetchL1Plugin_logic_banks_1_read_cmd_valid;
  wire       [8:0]    FetchL1Plugin_logic_banks_1_read_cmd_payload;
  (* keep , syn_keep *) wire       [63:0]   FetchL1Plugin_logic_banks_1_read_rsp /* synthesis syn_keep = 1 */ ;
  reg        [1:0]    FetchL1Plugin_logic_waysWrite_mask;
  reg        [5:0]    FetchL1Plugin_logic_waysWrite_address;
  reg                 FetchL1Plugin_logic_waysWrite_tag_loaded;
  reg                 FetchL1Plugin_logic_waysWrite_tag_error;
  reg        [19:0]   FetchL1Plugin_logic_waysWrite_tag_address;
  wire                FetchL1Plugin_logic_ways_0_read_cmd_valid;
  wire       [5:0]    FetchL1Plugin_logic_ways_0_read_cmd_payload;
  (* keep , syn_keep *) wire                FetchL1Plugin_logic_ways_0_read_rsp_loaded /* synthesis syn_keep = 1 */ ;
  (* keep , syn_keep *) wire                FetchL1Plugin_logic_ways_0_read_rsp_error /* synthesis syn_keep = 1 */ ;
  (* keep , syn_keep *) wire       [19:0]   FetchL1Plugin_logic_ways_0_read_rsp_address /* synthesis syn_keep = 1 */ ;
  wire       [21:0]   _zz_FetchL1Plugin_logic_ways_0_read_rsp_loaded;
  wire                FetchL1Plugin_logic_ways_1_read_cmd_valid;
  wire       [5:0]    FetchL1Plugin_logic_ways_1_read_cmd_payload;
  (* keep , syn_keep *) wire                FetchL1Plugin_logic_ways_1_read_rsp_loaded /* synthesis syn_keep = 1 */ ;
  (* keep , syn_keep *) wire                FetchL1Plugin_logic_ways_1_read_rsp_error /* synthesis syn_keep = 1 */ ;
  (* keep , syn_keep *) wire       [19:0]   FetchL1Plugin_logic_ways_1_read_rsp_address /* synthesis syn_keep = 1 */ ;
  wire       [21:0]   _zz_FetchL1Plugin_logic_ways_1_read_rsp_loaded;
  reg                 FetchL1Plugin_logic_plru_write_valid;
  reg        [5:0]    FetchL1Plugin_logic_plru_write_payload_address;
  reg        [0:0]    FetchL1Plugin_logic_plru_write_payload_data_0;
  wire                FetchL1Plugin_logic_plru_read_cmd_valid;
  wire       [5:0]    FetchL1Plugin_logic_plru_read_cmd_payload;
  (* keep , syn_keep *) wire       [0:0]    FetchL1Plugin_logic_plru_read_rsp_0 /* synthesis syn_keep = 1 */ ;
  wire                FetchL1Plugin_logic_invalidate_cmd_valid;
  wire                FetchL1Plugin_logic_invalidate_cmd_ready;
  reg                 FetchL1Plugin_logic_invalidate_canStart;
  reg        [6:0]    FetchL1Plugin_logic_invalidate_counter;
  wire       [6:0]    FetchL1Plugin_logic_invalidate_counterIncr;
  wire                FetchL1Plugin_logic_invalidate_done;
  wire                FetchL1Plugin_logic_invalidate_last;
  reg                 FetchL1Plugin_logic_invalidate_firstEver;
  wire                when_FetchL1Plugin_l220;
  wire                when_FetchL1Plugin_l227;
  wire                when_FetchL1Plugin_l232;
  wire                fetch_logic_ctrls_0_haltRequest_FetchL1Plugin_l233;
  reg                 FetchL1Plugin_logic_refill_start_valid;
  wire       [31:0]   FetchL1Plugin_logic_refill_start_address;
  wire       [0:0]    FetchL1Plugin_logic_refill_start_wayToAllocate;
  wire                FetchL1Plugin_logic_refill_start_isIo;
  reg                 FetchL1Plugin_logic_refill_slots_0_valid;
  reg                 FetchL1Plugin_logic_refill_slots_0_cmdSent;
  (* keep , syn_keep *) reg        [31:0]   FetchL1Plugin_logic_refill_slots_0_address /* synthesis syn_keep = 1 */ ;
  reg                 FetchL1Plugin_logic_refill_slots_0_isIo;
  reg        [0:0]    FetchL1Plugin_logic_refill_slots_0_wayToAllocate;
  reg        [0:0]    FetchL1Plugin_logic_refill_slots_0_priority;
  wire                FetchL1Plugin_logic_refill_slots_0_askCmd;
  reg        [31:0]   FetchL1Plugin_logic_refill_pushCounter;
  wire                FetchL1Plugin_logic_refill_hazard;
  wire                when_FetchL1Plugin_l271;
  wire                when_FetchL1Plugin_l293;
  wire       [0:0]    FetchL1Plugin_logic_refill_onCmd_oh;
  (* keep , syn_keep *) reg        [2:0]    FetchL1Plugin_logic_refill_onRsp_wordIndex /* synthesis syn_keep = 1 */ ;
  wire                FetchL1Plugin_logic_refill_onRsp_holdHarts;
  wire                fetch_logic_ctrls_0_haltRequest_FetchL1Plugin_l317;
  reg                 FetchL1Plugin_logic_refill_onRsp_firstCycle;
  wire                FetchL1Plugin_logic_bus_rsp_fire;
  wire       [0:0]    FetchL1Plugin_logic_refill_onRsp_wayToAllocate;
  wire       [31:0]   FetchL1Plugin_logic_refill_onRsp_address;
  wire                when_FetchL1Plugin_l324;
  wire                when_FetchL1Plugin_l350;
  wire                FetchL1Plugin_logic_cmd_doIt;
  wire                FetchL1Plugin_logic_hits_w_0_indirect_wayTlbHits_0;
  wire                FetchL1Plugin_logic_hits_w_0_indirect_wayTlbHits_1;
  wire                FetchL1Plugin_logic_hits_w_0_indirect_wayTlbHits_2;
  wire                FetchL1Plugin_logic_hits_w_0_indirect_translatedHits;
  wire                FetchL1Plugin_logic_hits_w_0_indirect_bypassHits;
  wire                FetchL1Plugin_logic_hits_w_1_indirect_wayTlbHits_0;
  wire                FetchL1Plugin_logic_hits_w_1_indirect_wayTlbHits_1;
  wire                FetchL1Plugin_logic_hits_w_1_indirect_wayTlbHits_2;
  wire                FetchL1Plugin_logic_hits_w_1_indirect_translatedHits;
  wire                FetchL1Plugin_logic_hits_w_1_indirect_bypassHits;
  wire       [31:0]   FetchL1Plugin_logic_ctrl_pmaPort_cmd_address;
  wire                FetchL1Plugin_logic_ctrl_pmaPort_rsp_fault;
  wire                FetchL1Plugin_logic_ctrl_pmaPort_rsp_io;
  wire       [0:0]    FetchL1Plugin_logic_ctrl_plruLogic_core_io_context_state_0;
  wire       [0:0]    FetchL1Plugin_logic_ctrl_plruLogic_core_io_evict_id;
  wire       [0:0]    FetchL1Plugin_logic_ctrl_plruLogic_core_io_update_id;
  wire       [0:0]    FetchL1Plugin_logic_ctrl_plruLogic_core_io_update_state_0;
  wire                FetchL1Plugin_logic_ctrl_plruLogic_core_evict_sel_0;
  wire                FetchL1Plugin_logic_ctrl_plruLogic_core_evict_logic_0_state;
  wire                FetchL1Plugin_logic_ctrl_plruLogic_buffer_valid;
  wire       [5:0]    FetchL1Plugin_logic_ctrl_plruLogic_buffer_payload_address;
  wire       [0:0]    FetchL1Plugin_logic_ctrl_plruLogic_buffer_payload_data_0;
  reg                 FetchL1Plugin_logic_ctrl_plruLogic_buffer_regNext_valid;
  reg        [5:0]    FetchL1Plugin_logic_ctrl_plruLogic_buffer_regNext_payload_address;
  reg        [0:0]    FetchL1Plugin_logic_ctrl_plruLogic_buffer_regNext_payload_data_0;
  wire                FetchL1Plugin_logic_ctrl_dataAccessFault;
  reg                 FetchL1Plugin_logic_ctrl_trapSent;
  reg                 FetchL1Plugin_logic_ctrl_allowRefill;
  wire                when_FetchL1Plugin_l483;
  wire                when_FetchL1Plugin_l489;
  wire                when_FetchL1Plugin_l496;
  wire                when_FetchL1Plugin_l529;
  wire                when_FetchL1Plugin_l542;
  wire                when_FetchL1Plugin_l546;
  reg                 FetchL1Plugin_logic_ctrl_firstCycle;
  wire                when_FetchL1Plugin_l550;
  wire                when_FetchL1Plugin_l567;
  reg        [9:0]    FetchL1Plugin_logic_initializer_counter;
  wire                FetchL1Plugin_logic_initializer_busy;
  reg        [3:0]    LsuPlugin_logic_trapPort_payload_code;
  reg        [2:0]    LsuPlugin_logic_trapPort_payload_arg;
  wire       [0:0]    LsuPlugin_logic_trapPort_payload_laneAge;
  reg                 LsuPlugin_logic_flushPort_valid;
  wire       [15:0]   LsuPlugin_logic_flushPort_payload_uopId;
  wire       [0:0]    LsuPlugin_logic_flushPort_payload_laneAge;
  wire                LsuPlugin_logic_flushPort_payload_self;
  wire                LsuPlugin_logic_commitProbe_valid;
  wire       [31:0]   LsuPlugin_logic_commitProbe_payload_pc;
  wire       [31:0]   LsuPlugin_logic_commitProbe_payload_address;
  wire                LsuPlugin_logic_commitProbe_payload_load;
  wire                LsuPlugin_logic_commitProbe_payload_store;
  wire                LsuPlugin_logic_commitProbe_payload_trap;
  wire                LsuPlugin_logic_commitProbe_payload_io;
  wire                LsuPlugin_logic_commitProbe_payload_prefetchFailed;
  wire                LsuPlugin_logic_commitProbe_payload_miss;
  wire                LsuPlugin_logic_iwb_valid;
  reg        [31:0]   LsuPlugin_logic_iwb_payload;
  wire                toplevel_execute_lane0_ctrls_0_upIsCancel;
  wire                toplevel_execute_lane0_ctrls_0_downIsCancel;
  wire                LsuPlugin_logic_bus_cmd_valid;
  wire                LsuPlugin_logic_bus_cmd_ready;
  wire                LsuPlugin_logic_bus_cmd_payload_write;
  wire       [31:0]   LsuPlugin_logic_bus_cmd_payload_address;
  wire       [31:0]   LsuPlugin_logic_bus_cmd_payload_data;
  wire       [1:0]    LsuPlugin_logic_bus_cmd_payload_size;
  wire       [3:0]    LsuPlugin_logic_bus_cmd_payload_mask;
  wire                LsuPlugin_logic_bus_cmd_payload_io;
  wire                LsuPlugin_logic_bus_cmd_payload_fromHart;
  wire       [15:0]   LsuPlugin_logic_bus_cmd_payload_uopId;
  wire                LsuPlugin_logic_bus_rsp_valid;
  wire                LsuPlugin_logic_bus_rsp_payload_error;
  wire       [31:0]   LsuPlugin_logic_bus_rsp_payload_data;
  wire                LsuPlugin_logic_flusher_wantExit;
  reg                 LsuPlugin_logic_flusher_wantStart;
  wire                LsuPlugin_logic_flusher_wantKill;
  reg        [6:0]    LsuPlugin_logic_flusher_cmdCounter;
  wire                LsuPlugin_logic_flusher_inflight;
  reg                 PrivilegedPlugin_logic_harts_0_xretAwayFromMachine;
  wire       [1:0]    PrivilegedPlugin_logic_harts_0_commitMask;
  reg                 PrivilegedPlugin_logic_harts_0_int_pending;
  reg        [1:0]    PrivilegedPlugin_logic_harts_0_privilege;
  wire                PrivilegedPlugin_logic_harts_0_withMachinePrivilege;
  wire                PrivilegedPlugin_logic_harts_0_withSupervisorPrivilege;
  wire                PrivilegedPlugin_logic_harts_0_hartRunning;
  wire                PrivilegedPlugin_logic_harts_0_debugMode;
  wire                when_CsrService_l188;
  reg                 PrivilegedPlugin_logic_harts_0_m_status_mie;
  reg                 PrivilegedPlugin_logic_harts_0_m_status_mpie;
  reg        [1:0]    PrivilegedPlugin_logic_harts_0_m_status_mpp;
  reg        [1:0]    PrivilegedPlugin_logic_harts_0_m_status_fs;
  reg                 PrivilegedPlugin_logic_harts_0_m_status_sd;
  reg                 PrivilegedPlugin_logic_harts_0_m_status_tsr;
  reg                 PrivilegedPlugin_logic_harts_0_m_status_tvm;
  reg                 PrivilegedPlugin_logic_harts_0_m_status_tw;
  wire                when_PrivilegedPlugin_l533;
  wire                _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue;
  wire                _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_1;
  wire                when_CsrService_l166;
  reg                 PrivilegedPlugin_logic_harts_0_m_cause_interrupt;
  reg        [3:0]    PrivilegedPlugin_logic_harts_0_m_cause_code;
  wire                _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_2;
  reg                 PrivilegedPlugin_logic_harts_0_m_ip_meip;
  reg                 PrivilegedPlugin_logic_harts_0_m_ip_mtip;
  reg                 PrivilegedPlugin_logic_harts_0_m_ip_msip;
  wire                _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_3;
  reg                 PrivilegedPlugin_logic_harts_0_m_ie_meie;
  reg                 PrivilegedPlugin_logic_harts_0_m_ie_mtie;
  reg                 PrivilegedPlugin_logic_harts_0_m_ie_msie;
  wire                _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_4;
  reg                 PrivilegedPlugin_logic_harts_0_m_edeleg_iam;
  reg                 PrivilegedPlugin_logic_harts_0_m_edeleg_bp;
  reg                 PrivilegedPlugin_logic_harts_0_m_edeleg_eu;
  reg                 PrivilegedPlugin_logic_harts_0_m_edeleg_es;
  reg                 PrivilegedPlugin_logic_harts_0_m_edeleg_ipf;
  reg                 PrivilegedPlugin_logic_harts_0_m_edeleg_lpf;
  reg                 PrivilegedPlugin_logic_harts_0_m_edeleg_spf;
  wire                _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_5;
  reg                 PrivilegedPlugin_logic_harts_0_m_ideleg_st;
  reg                 PrivilegedPlugin_logic_harts_0_m_ideleg_se;
  reg                 PrivilegedPlugin_logic_harts_0_m_ideleg_ss;
  wire                _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_6;
  wire                _zz_when_TrapPlugin_l195;
  wire                _zz_when_TrapPlugin_l195_1;
  wire                _zz_when_TrapPlugin_l195_2;
  reg                 PrivilegedPlugin_logic_harts_0_s_cause_interrupt;
  reg        [3:0]    PrivilegedPlugin_logic_harts_0_s_cause_code;
  wire                _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_7;
  reg                 PrivilegedPlugin_logic_harts_0_s_status_sie;
  reg                 PrivilegedPlugin_logic_harts_0_s_status_spie;
  reg        [0:0]    PrivilegedPlugin_logic_harts_0_s_status_spp;
  wire                _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_8;
  wire                _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_9;
  reg                 PrivilegedPlugin_logic_harts_0_s_ip_seipSoft;
  reg                 PrivilegedPlugin_logic_harts_0_s_ip_seipInput;
  wire                PrivilegedPlugin_logic_harts_0_s_ip_seipOr;
  reg                 PrivilegedPlugin_logic_harts_0_s_ip_stip;
  reg                 PrivilegedPlugin_logic_harts_0_s_ip_ssip;
  wire                PrivilegedPlugin_logic_harts_0_s_ip_seipMasked;
  wire                PrivilegedPlugin_logic_harts_0_s_ip_stipMasked;
  wire                PrivilegedPlugin_logic_harts_0_s_ip_ssipMasked;
  reg                 PrivilegedPlugin_logic_harts_0_s_ie_seie;
  reg                 PrivilegedPlugin_logic_harts_0_s_ie_stie;
  reg                 PrivilegedPlugin_logic_harts_0_s_ie_ssie;
  wire                _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_10;
  wire                _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_11;
  wire                _zz_when_TrapPlugin_l195_3;
  wire                _zz_when_TrapPlugin_l195_4;
  wire                _zz_when_TrapPlugin_l195_5;
  wire       [1:0]    PrivilegedPlugin_logic_defaultTrap_csrPrivilege;
  wire                PrivilegedPlugin_logic_defaultTrap_csrReadOnly;
  wire                when_PrivilegedPlugin_l679;
  reg                 GSharePlugin_logic_mem_write_valid;
  reg        [11:0]   GSharePlugin_logic_mem_write_payload_address;
  reg        [1:0]    GSharePlugin_logic_mem_write_payload_data_0;
  reg        [1:0]    GSharePlugin_logic_mem_write_payload_data_1;
  reg        [1:0]    GSharePlugin_logic_mem_write_payload_data_2;
  reg        [1:0]    GSharePlugin_logic_mem_write_payload_data_3;
  wire       [11:0]   _zz_fetch_logic_ctrls_0_down_GSharePlugin_logic_HASH;
  wire       [7:0]    _zz_fetch_logic_ctrls_1_down_GSharePlugin_GSHARE_COUNTER_0;
  wire                when_GSharePlugin_l82;
  reg        [1:0]    BtbPlugin_logic_ras_ptr_push;
  reg        [1:0]    BtbPlugin_logic_ras_ptr_pop;
  reg                 BtbPlugin_logic_ras_ptr_pushIt;
  reg                 BtbPlugin_logic_ras_ptr_popIt;
  wire                BtbPlugin_logic_ras_readIt;
  reg        [30:0]   BtbPlugin_logic_ras_read;
  reg                 BtbPlugin_logic_ras_write_valid;
  reg        [1:0]    BtbPlugin_logic_ras_write_payload_address;
  reg        [30:0]   BtbPlugin_logic_ras_write_payload_data;
  wire       [9:0]    WhiteboxerPlugin_logic_fetch_fetchId;
  wire                WhiteboxerPlugin_logic_decodes_0_fire;
  reg                 toplevel_decode_ctrls_0_up_LANE_SEL_0_regNext;
  wire                when_CtrlLaneApi_l46;
  wire                WhiteboxerPlugin_logic_decodes_0_spawn;
  wire       [63:0]   WhiteboxerPlugin_logic_decodes_0_pc;
  wire       [9:0]    WhiteboxerPlugin_logic_decodes_0_fetchId;
  wire       [9:0]    WhiteboxerPlugin_logic_decodes_0_decodeId;
  wire                WhiteboxerPlugin_logic_decodes_1_fire;
  reg                 toplevel_decode_ctrls_0_up_LANE_SEL_1_regNext;
  wire                when_CtrlLaneApi_l46_1;
  wire                WhiteboxerPlugin_logic_decodes_1_spawn;
  wire       [63:0]   WhiteboxerPlugin_logic_decodes_1_pc;
  wire       [9:0]    WhiteboxerPlugin_logic_decodes_1_fetchId;
  wire       [9:0]    WhiteboxerPlugin_logic_decodes_1_decodeId;
  wire       [15:0]   early0_BranchPlugin_logic_flushPort_payload_uopId;
  wire       [0:0]    early0_BranchPlugin_logic_flushPort_payload_laneAge;
  wire                early0_BranchPlugin_logic_flushPort_payload_self;
  wire                early0_BranchPlugin_logic_alu_expectedMsb;
  wire       [2:0]    switch_Misc_l241;
  reg                 _zz_toplevel_execute_ctrl3_down_early0_BranchPlugin_logic_jumpLogic_COND_lane0;
  reg                 _zz_toplevel_execute_ctrl3_down_early0_BranchPlugin_logic_jumpLogic_COND_lane0_1;
  wire                early0_BranchPlugin_logic_jumpLogic_wrongCond;
  wire                early0_BranchPlugin_logic_jumpLogic_needFix;
  wire                early0_BranchPlugin_logic_jumpLogic_doIt;
  wire       [11:0]   early0_BranchPlugin_logic_jumpLogic_history_fetched;
  wire       [11:0]   early0_BranchPlugin_logic_jumpLogic_history_next;
  wire       [1:0]    early0_BranchPlugin_logic_jumpLogic_history_fromFetch_slice;
  wire       [11:0]   early0_BranchPlugin_logic_jumpLogic_history_fromFetch_shifter;
  wire                when_BranchPlugin_l206;
  wire                when_BranchPlugin_l206_1;
  wire                when_BranchPlugin_l206_2;
  wire                when_BranchPlugin_l210;
  wire                early0_BranchPlugin_logic_jumpLogic_rdLink;
  wire                early0_BranchPlugin_logic_jumpLogic_rs1Link;
  wire                early0_BranchPlugin_logic_jumpLogic_rdEquRs1;
  wire       [15:0]   CsrAccessPlugin_logic_flushPort_payload_uopId;
  wire       [0:0]    CsrAccessPlugin_logic_flushPort_payload_laneAge;
  wire                CsrAccessPlugin_logic_flushPort_payload_self;
  reg                 CsrAccessPlugin_logic_trapPort_valid;
  reg                 CsrAccessPlugin_logic_trapPort_payload_exception;
  wire       [31:0]   CsrAccessPlugin_logic_trapPort_payload_tval;
  reg        [3:0]    CsrAccessPlugin_logic_trapPort_payload_code;
  wire       [2:0]    CsrAccessPlugin_logic_trapPort_payload_arg;
  wire       [0:0]    CsrAccessPlugin_logic_trapPort_payload_laneAge;
  wire       [15:0]   early0_EnvPlugin_logic_flushPort_payload_uopId;
  wire       [0:0]    early0_EnvPlugin_logic_flushPort_payload_laneAge;
  wire                early0_EnvPlugin_logic_flushPort_payload_self;
  wire       [1:0]    early0_EnvPlugin_logic_exe_privilege;
  wire       [1:0]    early0_EnvPlugin_logic_exe_xretPriv;
  reg                 early0_EnvPlugin_logic_exe_commit;
  wire                early0_EnvPlugin_logic_exe_retKo;
  wire                early0_EnvPlugin_logic_exe_vmaKo;
  wire                when_EnvPlugin_l83;
  wire                when_EnvPlugin_l92;
  wire                when_EnvPlugin_l107;
  wire                when_EnvPlugin_l116;
  wire                when_EnvPlugin_l120;
  wire       [15:0]   late0_BranchPlugin_logic_flushPort_payload_uopId;
  wire       [0:0]    late0_BranchPlugin_logic_flushPort_payload_laneAge;
  wire                late0_BranchPlugin_logic_flushPort_payload_self;
  wire       [15:0]   early1_BranchPlugin_logic_flushPort_payload_uopId;
  wire       [0:0]    early1_BranchPlugin_logic_flushPort_payload_laneAge;
  wire                early1_BranchPlugin_logic_flushPort_payload_self;
  wire                early1_BranchPlugin_logic_alu_expectedMsb;
  wire       [2:0]    switch_Misc_l241_1;
  reg                 _zz_toplevel_execute_ctrl3_down_early1_BranchPlugin_logic_jumpLogic_COND_lane1;
  reg                 _zz_toplevel_execute_ctrl3_down_early1_BranchPlugin_logic_jumpLogic_COND_lane1_1;
  wire                early1_BranchPlugin_logic_jumpLogic_wrongCond;
  wire                early1_BranchPlugin_logic_jumpLogic_needFix;
  wire                early1_BranchPlugin_logic_jumpLogic_doIt;
  wire       [11:0]   early1_BranchPlugin_logic_jumpLogic_history_fetched;
  wire       [11:0]   early1_BranchPlugin_logic_jumpLogic_history_next;
  wire       [1:0]    early1_BranchPlugin_logic_jumpLogic_history_fromFetch_slice;
  wire       [11:0]   early1_BranchPlugin_logic_jumpLogic_history_fromFetch_shifter;
  wire                when_BranchPlugin_l206_3;
  wire                when_BranchPlugin_l206_4;
  wire                when_BranchPlugin_l206_5;
  wire                when_BranchPlugin_l210_1;
  wire                early1_BranchPlugin_logic_jumpLogic_rdLink;
  wire                early1_BranchPlugin_logic_jumpLogic_rs1Link;
  wire                early1_BranchPlugin_logic_jumpLogic_rdEquRs1;
  wire       [15:0]   late1_BranchPlugin_logic_flushPort_payload_uopId;
  wire       [0:0]    late1_BranchPlugin_logic_flushPort_payload_laneAge;
  wire                late1_BranchPlugin_logic_flushPort_payload_self;
  wire                _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_12;
  wire       [0:0]    MmuPlugin_logic_satpModeWrite;
  wire                toplevel_execute_lane0_ctrls_1_upIsCancel;
  wire                toplevel_execute_lane0_ctrls_1_downIsCancel;
  reg        [31:0]   _zz_toplevel_execute_ctrl1_down_early0_SrcPlugin_SRC1_lane0;
  reg        [31:0]   _zz_toplevel_execute_ctrl1_down_early0_SrcPlugin_SRC2_lane0;
  reg        [31:0]   early0_SrcPlugin_logic_addsub_combined_rs2Patched;
  wire                lane0_IntFormatPlugin_logic_stages_0_wb_valid;
  wire       [31:0]   lane0_IntFormatPlugin_logic_stages_0_wb_payload;
  wire       [0:0]    lane0_IntFormatPlugin_logic_stages_0_hits;
  wire       [31:0]   lane0_IntFormatPlugin_logic_stages_0_raw;
  wire                lane0_IntFormatPlugin_logic_stages_1_wb_valid;
  wire       [31:0]   lane0_IntFormatPlugin_logic_stages_1_wb_payload;
  wire       [2:0]    lane0_IntFormatPlugin_logic_stages_1_hits;
  wire       [31:0]   lane0_IntFormatPlugin_logic_stages_1_raw;
  wire                lane0_IntFormatPlugin_logic_stages_2_wb_valid;
  reg        [31:0]   lane0_IntFormatPlugin_logic_stages_2_wb_payload;
  wire       [3:0]    lane0_IntFormatPlugin_logic_stages_2_hits;
  wire       [31:0]   lane0_IntFormatPlugin_logic_stages_2_raw;
  wire                lane0_IntFormatPlugin_logic_stages_2_segments_0_sign_sels_0;
  reg                 _zz_lane0_IntFormatPlugin_logic_stages_2_segments_0_sign_value;
  wire                lane0_IntFormatPlugin_logic_stages_2_segments_0_sign_value;
  wire                lane0_IntFormatPlugin_logic_stages_2_segments_0_doIt;
  wire                lane0_IntFormatPlugin_logic_stages_2_segments_1_sign_sels_0;
  wire                lane0_IntFormatPlugin_logic_stages_2_segments_1_sign_sels_1;
  reg                 _zz_lane0_IntFormatPlugin_logic_stages_2_segments_1_sign_value;
  wire                lane0_IntFormatPlugin_logic_stages_2_segments_1_sign_value;
  wire                lane0_IntFormatPlugin_logic_stages_2_segments_1_doIt;
  reg        [31:0]   _zz_toplevel_execute_ctrl3_down_late0_SrcPlugin_SRC1_lane0;
  reg        [31:0]   _zz_toplevel_execute_ctrl3_down_late0_SrcPlugin_SRC2_lane0;
  reg        [31:0]   late0_SrcPlugin_logic_addsub_combined_rs2Patched;
  wire                toplevel_execute_lane1_ctrls_1_upIsCancel;
  wire                toplevel_execute_lane1_ctrls_1_downIsCancel;
  reg        [31:0]   _zz_toplevel_execute_ctrl1_down_early1_SrcPlugin_SRC1_lane1;
  reg        [31:0]   _zz_toplevel_execute_ctrl1_down_early1_SrcPlugin_SRC2_lane1;
  reg        [31:0]   early1_SrcPlugin_logic_addsub_combined_rs2Patched;
  wire                lane1_IntFormatPlugin_logic_stages_0_wb_valid;
  wire       [31:0]   lane1_IntFormatPlugin_logic_stages_0_wb_payload;
  wire       [0:0]    lane1_IntFormatPlugin_logic_stages_0_hits;
  wire       [31:0]   lane1_IntFormatPlugin_logic_stages_0_raw;
  wire                lane1_IntFormatPlugin_logic_stages_1_wb_valid;
  wire       [31:0]   lane1_IntFormatPlugin_logic_stages_1_wb_payload;
  wire       [0:0]    lane1_IntFormatPlugin_logic_stages_1_hits;
  wire       [31:0]   lane1_IntFormatPlugin_logic_stages_1_raw;
  wire                lane1_IntFormatPlugin_logic_stages_2_wb_valid;
  wire       [31:0]   lane1_IntFormatPlugin_logic_stages_2_wb_payload;
  wire       [1:0]    lane1_IntFormatPlugin_logic_stages_2_hits;
  wire       [31:0]   lane1_IntFormatPlugin_logic_stages_2_raw;
  reg        [31:0]   _zz_toplevel_execute_ctrl3_down_late1_SrcPlugin_SRC1_lane1;
  reg        [31:0]   _zz_toplevel_execute_ctrl3_down_late1_SrcPlugin_SRC2_lane1;
  reg        [31:0]   late1_SrcPlugin_logic_addsub_combined_rs2Patched;
  wire                late0_BranchPlugin_logic_alu_expectedMsb;
  wire       [2:0]    switch_Misc_l241_2;
  reg                 _zz_toplevel_execute_ctrl4_down_late0_BranchPlugin_logic_jumpLogic_COND_lane0;
  reg                 _zz_toplevel_execute_ctrl4_down_late0_BranchPlugin_logic_jumpLogic_COND_lane0_1;
  wire                late0_BranchPlugin_logic_jumpLogic_wrongCond;
  wire                late0_BranchPlugin_logic_jumpLogic_needFix;
  wire                late0_BranchPlugin_logic_jumpLogic_doIt;
  wire       [11:0]   late0_BranchPlugin_logic_jumpLogic_history_fetched;
  wire       [11:0]   late0_BranchPlugin_logic_jumpLogic_history_next;
  wire       [1:0]    late0_BranchPlugin_logic_jumpLogic_history_fromFetch_slice;
  wire       [11:0]   late0_BranchPlugin_logic_jumpLogic_history_fromFetch_shifter;
  wire                when_BranchPlugin_l206_6;
  wire                when_BranchPlugin_l206_7;
  wire                when_BranchPlugin_l206_8;
  wire                when_BranchPlugin_l210_2;
  wire                late0_BranchPlugin_logic_jumpLogic_rdLink;
  wire                late0_BranchPlugin_logic_jumpLogic_rs1Link;
  wire                late0_BranchPlugin_logic_jumpLogic_rdEquRs1;
  wire                late0_BranchPlugin_logic_jumpLogic_learn_valid;
  reg                 late0_BranchPlugin_logic_jumpLogic_learn_ready;
  wire       [31:0]   late0_BranchPlugin_logic_jumpLogic_learn_payload_pcOnLastSlice;
  wire       [31:0]   late0_BranchPlugin_logic_jumpLogic_learn_payload_pcTarget;
  wire                late0_BranchPlugin_logic_jumpLogic_learn_payload_taken;
  wire                late0_BranchPlugin_logic_jumpLogic_learn_payload_isBranch;
  wire                late0_BranchPlugin_logic_jumpLogic_learn_payload_isPush;
  wire                late0_BranchPlugin_logic_jumpLogic_learn_payload_isPop;
  wire                late0_BranchPlugin_logic_jumpLogic_learn_payload_wasWrong;
  wire                late0_BranchPlugin_logic_jumpLogic_learn_payload_badPredictedTarget;
  wire       [11:0]   late0_BranchPlugin_logic_jumpLogic_learn_payload_history;
  wire       [15:0]   late0_BranchPlugin_logic_jumpLogic_learn_payload_uopId;
  wire       [1:0]    late0_BranchPlugin_logic_jumpLogic_learn_payload_ctx_GSharePlugin_GSHARE_COUNTER_0;
  wire       [1:0]    late0_BranchPlugin_logic_jumpLogic_learn_payload_ctx_GSharePlugin_GSHARE_COUNTER_1;
  wire       [1:0]    late0_BranchPlugin_logic_jumpLogic_learn_payload_ctx_GSharePlugin_GSHARE_COUNTER_2;
  wire       [1:0]    late0_BranchPlugin_logic_jumpLogic_learn_payload_ctx_GSharePlugin_GSHARE_COUNTER_3;
  wire                late1_BranchPlugin_logic_alu_expectedMsb;
  wire       [2:0]    switch_Misc_l241_3;
  reg                 _zz_toplevel_execute_ctrl4_down_late1_BranchPlugin_logic_jumpLogic_COND_lane1;
  reg                 _zz_toplevel_execute_ctrl4_down_late1_BranchPlugin_logic_jumpLogic_COND_lane1_1;
  wire                late1_BranchPlugin_logic_jumpLogic_wrongCond;
  wire                late1_BranchPlugin_logic_jumpLogic_needFix;
  wire                late1_BranchPlugin_logic_jumpLogic_doIt;
  wire       [11:0]   late1_BranchPlugin_logic_jumpLogic_history_fetched;
  wire       [11:0]   late1_BranchPlugin_logic_jumpLogic_history_next;
  wire       [1:0]    late1_BranchPlugin_logic_jumpLogic_history_fromFetch_slice;
  wire       [11:0]   late1_BranchPlugin_logic_jumpLogic_history_fromFetch_shifter;
  wire                when_BranchPlugin_l206_9;
  wire                when_BranchPlugin_l206_10;
  wire                when_BranchPlugin_l206_11;
  wire                when_BranchPlugin_l210_3;
  wire                late1_BranchPlugin_logic_jumpLogic_rdLink;
  wire                late1_BranchPlugin_logic_jumpLogic_rs1Link;
  wire                late1_BranchPlugin_logic_jumpLogic_rdEquRs1;
  wire                late1_BranchPlugin_logic_jumpLogic_learn_valid;
  reg                 late1_BranchPlugin_logic_jumpLogic_learn_ready;
  wire       [31:0]   late1_BranchPlugin_logic_jumpLogic_learn_payload_pcOnLastSlice;
  wire       [31:0]   late1_BranchPlugin_logic_jumpLogic_learn_payload_pcTarget;
  wire                late1_BranchPlugin_logic_jumpLogic_learn_payload_taken;
  wire                late1_BranchPlugin_logic_jumpLogic_learn_payload_isBranch;
  wire                late1_BranchPlugin_logic_jumpLogic_learn_payload_isPush;
  wire                late1_BranchPlugin_logic_jumpLogic_learn_payload_isPop;
  wire                late1_BranchPlugin_logic_jumpLogic_learn_payload_wasWrong;
  wire                late1_BranchPlugin_logic_jumpLogic_learn_payload_badPredictedTarget;
  wire       [11:0]   late1_BranchPlugin_logic_jumpLogic_learn_payload_history;
  wire       [15:0]   late1_BranchPlugin_logic_jumpLogic_learn_payload_uopId;
  wire       [1:0]    late1_BranchPlugin_logic_jumpLogic_learn_payload_ctx_GSharePlugin_GSHARE_COUNTER_0;
  wire       [1:0]    late1_BranchPlugin_logic_jumpLogic_learn_payload_ctx_GSharePlugin_GSHARE_COUNTER_1;
  wire       [1:0]    late1_BranchPlugin_logic_jumpLogic_learn_payload_ctx_GSharePlugin_GSHARE_COUNTER_2;
  wire       [1:0]    late1_BranchPlugin_logic_jumpLogic_learn_payload_ctx_GSharePlugin_GSHARE_COUNTER_3;
  wire                LearnPlugin_logic_learn_valid;
  wire       [31:0]   LearnPlugin_logic_learn_payload_pcOnLastSlice;
  wire       [31:0]   LearnPlugin_logic_learn_payload_pcTarget;
  wire                LearnPlugin_logic_learn_payload_taken;
  wire                LearnPlugin_logic_learn_payload_isBranch;
  wire                LearnPlugin_logic_learn_payload_isPush;
  wire                LearnPlugin_logic_learn_payload_isPop;
  wire                LearnPlugin_logic_learn_payload_wasWrong;
  wire                LearnPlugin_logic_learn_payload_badPredictedTarget;
  wire       [11:0]   LearnPlugin_logic_learn_payload_history;
  wire       [15:0]   LearnPlugin_logic_learn_payload_uopId;
  wire       [1:0]    LearnPlugin_logic_learn_payload_ctx_GSharePlugin_GSHARE_COUNTER_0;
  wire       [1:0]    LearnPlugin_logic_learn_payload_ctx_GSharePlugin_GSHARE_COUNTER_1;
  wire       [1:0]    LearnPlugin_logic_learn_payload_ctx_GSharePlugin_GSHARE_COUNTER_2;
  wire       [1:0]    LearnPlugin_logic_learn_payload_ctx_GSharePlugin_GSHARE_COUNTER_3;
  wire                late0_BranchPlugin_logic_jumpLogic_learn_m2sPipe_valid;
  wire                late0_BranchPlugin_logic_jumpLogic_learn_m2sPipe_ready;
  wire       [31:0]   late0_BranchPlugin_logic_jumpLogic_learn_m2sPipe_payload_pcOnLastSlice;
  wire       [31:0]   late0_BranchPlugin_logic_jumpLogic_learn_m2sPipe_payload_pcTarget;
  wire                late0_BranchPlugin_logic_jumpLogic_learn_m2sPipe_payload_taken;
  wire                late0_BranchPlugin_logic_jumpLogic_learn_m2sPipe_payload_isBranch;
  wire                late0_BranchPlugin_logic_jumpLogic_learn_m2sPipe_payload_isPush;
  wire                late0_BranchPlugin_logic_jumpLogic_learn_m2sPipe_payload_isPop;
  wire                late0_BranchPlugin_logic_jumpLogic_learn_m2sPipe_payload_wasWrong;
  wire                late0_BranchPlugin_logic_jumpLogic_learn_m2sPipe_payload_badPredictedTarget;
  wire       [11:0]   late0_BranchPlugin_logic_jumpLogic_learn_m2sPipe_payload_history;
  wire       [15:0]   late0_BranchPlugin_logic_jumpLogic_learn_m2sPipe_payload_uopId;
  wire       [1:0]    late0_BranchPlugin_logic_jumpLogic_learn_m2sPipe_payload_ctx_GSharePlugin_GSHARE_COUNTER_0;
  wire       [1:0]    late0_BranchPlugin_logic_jumpLogic_learn_m2sPipe_payload_ctx_GSharePlugin_GSHARE_COUNTER_1;
  wire       [1:0]    late0_BranchPlugin_logic_jumpLogic_learn_m2sPipe_payload_ctx_GSharePlugin_GSHARE_COUNTER_2;
  wire       [1:0]    late0_BranchPlugin_logic_jumpLogic_learn_m2sPipe_payload_ctx_GSharePlugin_GSHARE_COUNTER_3;
  reg                 late0_BranchPlugin_logic_jumpLogic_learn_rValid;
  reg        [31:0]   late0_BranchPlugin_logic_jumpLogic_learn_rData_pcOnLastSlice;
  reg        [31:0]   late0_BranchPlugin_logic_jumpLogic_learn_rData_pcTarget;
  reg                 late0_BranchPlugin_logic_jumpLogic_learn_rData_taken;
  reg                 late0_BranchPlugin_logic_jumpLogic_learn_rData_isBranch;
  reg                 late0_BranchPlugin_logic_jumpLogic_learn_rData_isPush;
  reg                 late0_BranchPlugin_logic_jumpLogic_learn_rData_isPop;
  reg                 late0_BranchPlugin_logic_jumpLogic_learn_rData_wasWrong;
  reg                 late0_BranchPlugin_logic_jumpLogic_learn_rData_badPredictedTarget;
  reg        [11:0]   late0_BranchPlugin_logic_jumpLogic_learn_rData_history;
  reg        [15:0]   late0_BranchPlugin_logic_jumpLogic_learn_rData_uopId;
  reg        [1:0]    late0_BranchPlugin_logic_jumpLogic_learn_rData_ctx_GSharePlugin_GSHARE_COUNTER_0;
  reg        [1:0]    late0_BranchPlugin_logic_jumpLogic_learn_rData_ctx_GSharePlugin_GSHARE_COUNTER_1;
  reg        [1:0]    late0_BranchPlugin_logic_jumpLogic_learn_rData_ctx_GSharePlugin_GSHARE_COUNTER_2;
  reg        [1:0]    late0_BranchPlugin_logic_jumpLogic_learn_rData_ctx_GSharePlugin_GSHARE_COUNTER_3;
  wire                when_Stream_l393;
  wire                late1_BranchPlugin_logic_jumpLogic_learn_m2sPipe_valid;
  wire                late1_BranchPlugin_logic_jumpLogic_learn_m2sPipe_ready;
  wire       [31:0]   late1_BranchPlugin_logic_jumpLogic_learn_m2sPipe_payload_pcOnLastSlice;
  wire       [31:0]   late1_BranchPlugin_logic_jumpLogic_learn_m2sPipe_payload_pcTarget;
  wire                late1_BranchPlugin_logic_jumpLogic_learn_m2sPipe_payload_taken;
  wire                late1_BranchPlugin_logic_jumpLogic_learn_m2sPipe_payload_isBranch;
  wire                late1_BranchPlugin_logic_jumpLogic_learn_m2sPipe_payload_isPush;
  wire                late1_BranchPlugin_logic_jumpLogic_learn_m2sPipe_payload_isPop;
  wire                late1_BranchPlugin_logic_jumpLogic_learn_m2sPipe_payload_wasWrong;
  wire                late1_BranchPlugin_logic_jumpLogic_learn_m2sPipe_payload_badPredictedTarget;
  wire       [11:0]   late1_BranchPlugin_logic_jumpLogic_learn_m2sPipe_payload_history;
  wire       [15:0]   late1_BranchPlugin_logic_jumpLogic_learn_m2sPipe_payload_uopId;
  wire       [1:0]    late1_BranchPlugin_logic_jumpLogic_learn_m2sPipe_payload_ctx_GSharePlugin_GSHARE_COUNTER_0;
  wire       [1:0]    late1_BranchPlugin_logic_jumpLogic_learn_m2sPipe_payload_ctx_GSharePlugin_GSHARE_COUNTER_1;
  wire       [1:0]    late1_BranchPlugin_logic_jumpLogic_learn_m2sPipe_payload_ctx_GSharePlugin_GSHARE_COUNTER_2;
  wire       [1:0]    late1_BranchPlugin_logic_jumpLogic_learn_m2sPipe_payload_ctx_GSharePlugin_GSHARE_COUNTER_3;
  reg                 late1_BranchPlugin_logic_jumpLogic_learn_rValid;
  reg        [31:0]   late1_BranchPlugin_logic_jumpLogic_learn_rData_pcOnLastSlice;
  reg        [31:0]   late1_BranchPlugin_logic_jumpLogic_learn_rData_pcTarget;
  reg                 late1_BranchPlugin_logic_jumpLogic_learn_rData_taken;
  reg                 late1_BranchPlugin_logic_jumpLogic_learn_rData_isBranch;
  reg                 late1_BranchPlugin_logic_jumpLogic_learn_rData_isPush;
  reg                 late1_BranchPlugin_logic_jumpLogic_learn_rData_isPop;
  reg                 late1_BranchPlugin_logic_jumpLogic_learn_rData_wasWrong;
  reg                 late1_BranchPlugin_logic_jumpLogic_learn_rData_badPredictedTarget;
  reg        [11:0]   late1_BranchPlugin_logic_jumpLogic_learn_rData_history;
  reg        [15:0]   late1_BranchPlugin_logic_jumpLogic_learn_rData_uopId;
  reg        [1:0]    late1_BranchPlugin_logic_jumpLogic_learn_rData_ctx_GSharePlugin_GSHARE_COUNTER_0;
  reg        [1:0]    late1_BranchPlugin_logic_jumpLogic_learn_rData_ctx_GSharePlugin_GSHARE_COUNTER_1;
  reg        [1:0]    late1_BranchPlugin_logic_jumpLogic_learn_rData_ctx_GSharePlugin_GSHARE_COUNTER_2;
  reg        [1:0]    late1_BranchPlugin_logic_jumpLogic_learn_rData_ctx_GSharePlugin_GSHARE_COUNTER_3;
  wire                when_Stream_l393_1;
  wire                streamArbiter_10_io_output_combStage_valid;
  wire                streamArbiter_10_io_output_combStage_ready;
  wire       [31:0]   streamArbiter_10_io_output_combStage_payload_pcOnLastSlice;
  wire       [31:0]   streamArbiter_10_io_output_combStage_payload_pcTarget;
  wire                streamArbiter_10_io_output_combStage_payload_taken;
  wire                streamArbiter_10_io_output_combStage_payload_isBranch;
  wire                streamArbiter_10_io_output_combStage_payload_isPush;
  wire                streamArbiter_10_io_output_combStage_payload_isPop;
  wire                streamArbiter_10_io_output_combStage_payload_wasWrong;
  wire                streamArbiter_10_io_output_combStage_payload_badPredictedTarget;
  wire       [11:0]   streamArbiter_10_io_output_combStage_payload_history;
  wire       [15:0]   streamArbiter_10_io_output_combStage_payload_uopId;
  wire       [1:0]    streamArbiter_10_io_output_combStage_payload_ctx_GSharePlugin_GSHARE_COUNTER_0;
  wire       [1:0]    streamArbiter_10_io_output_combStage_payload_ctx_GSharePlugin_GSHARE_COUNTER_1;
  wire       [1:0]    streamArbiter_10_io_output_combStage_payload_ctx_GSharePlugin_GSHARE_COUNTER_2;
  wire       [1:0]    streamArbiter_10_io_output_combStage_payload_ctx_GSharePlugin_GSHARE_COUNTER_3;
  wire                CsrRamPlugin_setup_initPort_valid;
  wire                CsrRamPlugin_setup_initPort_ready;
  wire       [2:0]    CsrRamPlugin_setup_initPort_address;
  wire       [31:0]   CsrRamPlugin_setup_initPort_data;
  wire       [11:0]   _zz_GSharePlugin_logic_onLearn_hash;
  wire       [11:0]   GSharePlugin_logic_onLearn_hash;
  wire       [1:0]    GSharePlugin_logic_onLearn_updated_0;
  wire       [1:0]    GSharePlugin_logic_onLearn_updated_1;
  wire       [1:0]    GSharePlugin_logic_onLearn_updated_2;
  wire       [1:0]    GSharePlugin_logic_onLearn_updated_3;
  wire       [1:0]    GSharePlugin_logic_onLearn_incrValue;
  reg                 GSharePlugin_logic_onLearn_overflow;
  wire                when_GSharePlugin_l104;
  wire                when_GSharePlugin_l104_1;
  wire                when_GSharePlugin_l104_2;
  wire                when_GSharePlugin_l104_3;
  reg        [12:0]   GSharePlugin_logic_initializer_counter;
  wire                GSharePlugin_logic_initializer_busy;
  wire       [7:0]    _zz_GSharePlugin_logic_mem_write_payload_data_0;
  wire       [15:0]   BtbPlugin_logic_onLearn_hash;
  reg                 BtbPlugin_logic_onLearn_port_valid;
  reg        [7:0]    BtbPlugin_logic_onLearn_port_payload_address;
  reg        [15:0]   BtbPlugin_logic_onLearn_port_payload_data_0_hash;
  reg        [0:0]    BtbPlugin_logic_onLearn_port_payload_data_0_sliceLow;
  wire       [30:0]   BtbPlugin_logic_onLearn_port_payload_data_0_pcTarget;
  reg                 BtbPlugin_logic_onLearn_port_payload_data_0_isBranch;
  reg                 BtbPlugin_logic_onLearn_port_payload_data_0_isPush;
  reg                 BtbPlugin_logic_onLearn_port_payload_data_0_isPop;
  reg        [15:0]   BtbPlugin_logic_onLearn_port_payload_data_1_hash;
  reg        [0:0]    BtbPlugin_logic_onLearn_port_payload_data_1_sliceLow;
  wire       [30:0]   BtbPlugin_logic_onLearn_port_payload_data_1_pcTarget;
  reg                 BtbPlugin_logic_onLearn_port_payload_data_1_isBranch;
  reg                 BtbPlugin_logic_onLearn_port_payload_data_1_isPush;
  reg                 BtbPlugin_logic_onLearn_port_payload_data_1_isPop;
  reg        [1:0]    BtbPlugin_logic_onLearn_port_payload_mask;
  wire                CsrRamPlugin_csrMapper_read_valid;
  wire                CsrRamPlugin_csrMapper_read_ready;
  wire       [2:0]    CsrRamPlugin_csrMapper_read_address;
  wire       [31:0]   CsrRamPlugin_csrMapper_read_data;
  wire                CsrRamPlugin_csrMapper_write_valid;
  wire                CsrRamPlugin_csrMapper_write_ready;
  wire       [2:0]    CsrRamPlugin_csrMapper_write_address;
  wire       [31:0]   CsrRamPlugin_csrMapper_write_data;
  reg        [15:0]   DecoderPlugin_logic_harts_0_uopId;
  wire                when_DecoderPlugin_l135;
  wire       [0:0]    DecoderPlugin_logic_interrupt_async;
  wire                when_DecoderPlugin_l143;
  reg        [0:0]    DecoderPlugin_logic_interrupt_buffered;
  wire                _zz_toplevel_decode_ctrls_1_down_DispatchPlugin_MAY_FLUSH_0;
  wire                _zz_toplevel_decode_ctrls_1_down_DispatchPlugin_logic_LANES_LAYER_HIT_0_0;
  wire                _zz_toplevel_decode_ctrls_1_down_DispatchPlugin_logic_LANES_LAYER_HIT_3_0;
  wire                DecoderPlugin_logic_laneLogic_0_interruptPending;
  reg                 DecoderPlugin_logic_laneLogic_0_trapPort_valid;
  reg                 DecoderPlugin_logic_laneLogic_0_trapPort_payload_exception;
  wire       [31:0]   DecoderPlugin_logic_laneLogic_0_trapPort_payload_tval;
  reg        [3:0]    DecoderPlugin_logic_laneLogic_0_trapPort_payload_code;
  wire       [2:0]    DecoderPlugin_logic_laneLogic_0_trapPort_payload_arg;
  wire       [1:0]    DecoderPlugin_logic_laneLogic_0_trapPort_payload_laneAge;
  wire                _zz_toplevel_decode_ctrls_1_down_DispatchPlugin_logic_LANES_LAYER_HIT_0_0_1;
  wire                DecoderPlugin_logic_laneLogic_0_fixer_isJb;
  wire                DecoderPlugin_logic_laneLogic_0_fixer_doIt;
  wire                DecoderPlugin_logic_laneLogic_0_completionPort_valid;
  wire       [15:0]   DecoderPlugin_logic_laneLogic_0_completionPort_payload_uopId;
  wire                DecoderPlugin_logic_laneLogic_0_completionPort_payload_trap;
  wire                DecoderPlugin_logic_laneLogic_0_completionPort_payload_commit;
  reg                 toplevel_decode_ctrls_1_up_LANE_SEL_0_regNext;
  wire                when_CtrlLaneApi_l46_2;
  wire                when_DecoderPlugin_l216;
  wire                DecoderPlugin_logic_laneLogic_0_flushPort_valid;
  wire       [15:0]   DecoderPlugin_logic_laneLogic_0_flushPort_payload_uopId;
  wire       [0:0]    DecoderPlugin_logic_laneLogic_0_flushPort_payload_laneAge;
  wire                DecoderPlugin_logic_laneLogic_0_flushPort_payload_self;
  wire                when_DecoderPlugin_l234;
  wire       [15:0]   DecoderPlugin_logic_laneLogic_0_uopIdBase;
  wire                _zz_toplevel_decode_ctrls_1_down_DispatchPlugin_MAY_FLUSH_1;
  wire                _zz_toplevel_decode_ctrls_1_down_DispatchPlugin_logic_LANES_LAYER_HIT_0_1;
  wire                _zz_toplevel_decode_ctrls_1_down_DispatchPlugin_logic_LANES_LAYER_HIT_3_1;
  wire                DecoderPlugin_logic_laneLogic_1_interruptPending;
  reg                 DecoderPlugin_logic_laneLogic_1_trapPort_valid;
  reg                 DecoderPlugin_logic_laneLogic_1_trapPort_payload_exception;
  wire       [31:0]   DecoderPlugin_logic_laneLogic_1_trapPort_payload_tval;
  reg        [3:0]    DecoderPlugin_logic_laneLogic_1_trapPort_payload_code;
  wire       [2:0]    DecoderPlugin_logic_laneLogic_1_trapPort_payload_arg;
  wire       [1:0]    DecoderPlugin_logic_laneLogic_1_trapPort_payload_laneAge;
  wire                _zz_toplevel_decode_ctrls_1_down_DispatchPlugin_logic_LANES_LAYER_HIT_0_1_1;
  wire                DecoderPlugin_logic_laneLogic_1_fixer_isJb;
  wire                DecoderPlugin_logic_laneLogic_1_fixer_doIt;
  wire                DecoderPlugin_logic_laneLogic_1_completionPort_valid;
  wire       [15:0]   DecoderPlugin_logic_laneLogic_1_completionPort_payload_uopId;
  wire                DecoderPlugin_logic_laneLogic_1_completionPort_payload_trap;
  wire                DecoderPlugin_logic_laneLogic_1_completionPort_payload_commit;
  reg                 toplevel_decode_ctrls_1_up_LANE_SEL_1_regNext;
  wire                when_CtrlLaneApi_l46_3;
  wire                when_DecoderPlugin_l216_1;
  wire                DecoderPlugin_logic_laneLogic_1_flushPort_valid;
  wire       [15:0]   DecoderPlugin_logic_laneLogic_1_flushPort_payload_uopId;
  wire       [0:0]    DecoderPlugin_logic_laneLogic_1_flushPort_payload_laneAge;
  wire                DecoderPlugin_logic_laneLogic_1_flushPort_payload_self;
  wire                when_DecoderPlugin_l234_1;
  wire       [15:0]   DecoderPlugin_logic_laneLogic_1_uopIdBase;
  wire       [2:0]    CsrRamPlugin_csrMapper_ramAddress;
  wire       [11:0]   _zz_CsrRamPlugin_csrMapper_ramAddress;
  reg                 CsrRamPlugin_csrMapper_withRead;
  wire                when_CsrRamPlugin_l77;
  reg                 CsrRamPlugin_csrMapper_doWrite;
  reg                 CsrRamPlugin_csrMapper_fired;
  wire                when_CsrRamPlugin_l84;
  wire                when_CsrRamPlugin_l88;
  wire       [1:0]    lane0_integer_WriteBackPlugin_logic_stages_0_hits;
  wire       [31:0]   lane0_integer_WriteBackPlugin_logic_stages_0_muxed;
  wire                lane0_integer_WriteBackPlugin_logic_stages_0_write_valid;
  wire       [15:0]   lane0_integer_WriteBackPlugin_logic_stages_0_write_payload_uopId;
  wire       [31:0]   lane0_integer_WriteBackPlugin_logic_stages_0_write_payload_data;
  wire       [0:0]    lane0_integer_WriteBackPlugin_logic_stages_1_hits;
  wire       [31:0]   lane0_integer_WriteBackPlugin_logic_stages_1_muxed;
  wire       [31:0]   lane0_integer_WriteBackPlugin_logic_stages_1_merged;
  wire                lane0_integer_WriteBackPlugin_logic_stages_1_write_valid;
  wire       [15:0]   lane0_integer_WriteBackPlugin_logic_stages_1_write_payload_uopId;
  wire       [31:0]   lane0_integer_WriteBackPlugin_logic_stages_1_write_payload_data;
  wire       [1:0]    lane0_integer_WriteBackPlugin_logic_stages_2_hits;
  wire       [31:0]   lane0_integer_WriteBackPlugin_logic_stages_2_muxed;
  wire       [31:0]   lane0_integer_WriteBackPlugin_logic_stages_2_merged;
  wire                lane0_integer_WriteBackPlugin_logic_stages_2_write_valid;
  wire       [15:0]   lane0_integer_WriteBackPlugin_logic_stages_2_write_payload_uopId;
  wire       [31:0]   lane0_integer_WriteBackPlugin_logic_stages_2_write_payload_data;
  wire                lane0_integer_WriteBackPlugin_logic_write_port_valid;
  wire       [4:0]    lane0_integer_WriteBackPlugin_logic_write_port_address;
  wire       [31:0]   lane0_integer_WriteBackPlugin_logic_write_port_data;
  wire       [15:0]   lane0_integer_WriteBackPlugin_logic_write_port_uopId;
  wire       [1:0]    lane1_integer_WriteBackPlugin_logic_stages_0_hits;
  wire       [31:0]   lane1_integer_WriteBackPlugin_logic_stages_0_muxed;
  wire                lane1_integer_WriteBackPlugin_logic_stages_0_write_valid;
  wire       [15:0]   lane1_integer_WriteBackPlugin_logic_stages_0_write_payload_uopId;
  wire       [31:0]   lane1_integer_WriteBackPlugin_logic_stages_0_write_payload_data;
  wire       [0:0]    lane1_integer_WriteBackPlugin_logic_stages_1_hits;
  wire       [31:0]   lane1_integer_WriteBackPlugin_logic_stages_1_muxed;
  wire       [31:0]   lane1_integer_WriteBackPlugin_logic_stages_1_merged;
  wire                lane1_integer_WriteBackPlugin_logic_stages_1_write_valid;
  wire       [15:0]   lane1_integer_WriteBackPlugin_logic_stages_1_write_payload_uopId;
  wire       [31:0]   lane1_integer_WriteBackPlugin_logic_stages_1_write_payload_data;
  wire       [1:0]    lane1_integer_WriteBackPlugin_logic_stages_2_hits;
  wire       [31:0]   lane1_integer_WriteBackPlugin_logic_stages_2_muxed;
  wire       [31:0]   lane1_integer_WriteBackPlugin_logic_stages_2_merged;
  wire                lane1_integer_WriteBackPlugin_logic_stages_2_write_valid;
  wire       [15:0]   lane1_integer_WriteBackPlugin_logic_stages_2_write_payload_uopId;
  wire       [31:0]   lane1_integer_WriteBackPlugin_logic_stages_2_write_payload_data;
  wire                lane1_integer_WriteBackPlugin_logic_write_port_valid;
  wire       [4:0]    lane1_integer_WriteBackPlugin_logic_write_port_address;
  wire       [31:0]   lane1_integer_WriteBackPlugin_logic_write_port_data;
  wire       [15:0]   lane1_integer_WriteBackPlugin_logic_write_port_uopId;
  reg                 DispatchPlugin_logic_slots_0_ctx_valid;
  reg        [3:0]    DispatchPlugin_logic_slots_0_ctx_laneLayerHits;
  reg        [31:0]   DispatchPlugin_logic_slots_0_ctx_uop;
  reg                 DispatchPlugin_logic_slots_0_ctx_hm_Prediction_ALIGNED_JUMPED;
  reg        [31:0]   DispatchPlugin_logic_slots_0_ctx_hm_Prediction_ALIGNED_JUMPED_PC;
  reg        [3:0]    DispatchPlugin_logic_slots_0_ctx_hm_Prediction_ALIGNED_SLICES_TAKEN;
  reg        [3:0]    DispatchPlugin_logic_slots_0_ctx_hm_Prediction_ALIGNED_SLICES_BRANCH;
  reg        [1:0]    DispatchPlugin_logic_slots_0_ctx_hm_GSharePlugin_GSHARE_COUNTER_0;
  reg        [1:0]    DispatchPlugin_logic_slots_0_ctx_hm_GSharePlugin_GSHARE_COUNTER_1;
  reg        [1:0]    DispatchPlugin_logic_slots_0_ctx_hm_GSharePlugin_GSHARE_COUNTER_2;
  reg        [1:0]    DispatchPlugin_logic_slots_0_ctx_hm_GSharePlugin_GSHARE_COUNTER_3;
  reg        [11:0]   DispatchPlugin_logic_slots_0_ctx_hm_Prediction_BRANCH_HISTORY;
  reg                 DispatchPlugin_logic_slots_0_ctx_hm_DispatchPlugin_FENCE_OLDER;
  reg                 DispatchPlugin_logic_slots_0_ctx_hm_DispatchPlugin_MAY_FLUSH;
  reg                 DispatchPlugin_logic_slots_0_ctx_hm_DispatchPlugin_DONT_FLUSH;
  reg                 DispatchPlugin_logic_slots_0_ctx_hm_DispatchPlugin_DONT_FLUSH_FROM_LANES;
  reg        [0:0]    DispatchPlugin_logic_slots_0_ctx_hm_Decode_INSTRUCTION_SLICE_COUNT;
  reg                 DispatchPlugin_logic_slots_0_ctx_hm_DONT_FLUSH_PRECISE_3;
  reg                 DispatchPlugin_logic_slots_0_ctx_hm_DONT_FLUSH_PRECISE_4;
  reg        [31:0]   DispatchPlugin_logic_slots_0_ctx_hm_PC;
  reg                 DispatchPlugin_logic_slots_0_ctx_hm_TRAP;
  reg        [15:0]   DispatchPlugin_logic_slots_0_ctx_hm_Decode_UOP_ID;
  reg                 DispatchPlugin_logic_slots_0_ctx_hm_RS1_ENABLE;
  reg        [4:0]    DispatchPlugin_logic_slots_0_ctx_hm_RS1_PHYS;
  reg                 DispatchPlugin_logic_slots_0_ctx_hm_RS2_ENABLE;
  reg        [4:0]    DispatchPlugin_logic_slots_0_ctx_hm_RS2_PHYS;
  reg                 DispatchPlugin_logic_slots_0_ctx_hm_RD_ENABLE;
  reg        [4:0]    DispatchPlugin_logic_slots_0_ctx_hm_RD_PHYS;
  reg                 DispatchPlugin_logic_slots_0_ctx_hm_DispatchPlugin_logic_hcs_0_onRs_0_ENABLES_0;
  reg                 DispatchPlugin_logic_slots_0_ctx_hm_DispatchPlugin_logic_hcs_0_onRs_1_ENABLES_0;
  reg                 DispatchPlugin_logic_slots_0_ctx_hm_DispatchPlugin_logic_hcs_1_onRs_0_ENABLES_0;
  reg                 DispatchPlugin_logic_slots_0_ctx_hm_DispatchPlugin_logic_hcs_1_onRs_1_ENABLES_0;
  reg                 DispatchPlugin_logic_slots_0_ctx_hm_DispatchPlugin_logic_hcs_1_onRs_1_ENABLES_1;
  reg                 DispatchPlugin_logic_slots_0_ctx_hm_DispatchPlugin_logic_hcs_2_onRs_0_ENABLES_0;
  reg                 DispatchPlugin_logic_slots_0_ctx_hm_DispatchPlugin_logic_hcs_2_onRs_1_ENABLES_0;
  reg                 DispatchPlugin_logic_slots_0_ctx_hm_DispatchPlugin_logic_hcs_3_onRs_0_ENABLES_0;
  reg                 DispatchPlugin_logic_slots_0_ctx_hm_DispatchPlugin_logic_hcs_3_onRs_1_ENABLES_0;
  wire                DispatchPlugin_logic_candidates_0_ctx_valid;
  wire       [3:0]    DispatchPlugin_logic_candidates_0_ctx_laneLayerHits;
  wire       [31:0]   DispatchPlugin_logic_candidates_0_ctx_uop;
  wire                DispatchPlugin_logic_candidates_0_ctx_hm_Prediction_ALIGNED_JUMPED;
  wire       [31:0]   DispatchPlugin_logic_candidates_0_ctx_hm_Prediction_ALIGNED_JUMPED_PC;
  wire       [3:0]    DispatchPlugin_logic_candidates_0_ctx_hm_Prediction_ALIGNED_SLICES_TAKEN;
  wire       [3:0]    DispatchPlugin_logic_candidates_0_ctx_hm_Prediction_ALIGNED_SLICES_BRANCH;
  wire       [1:0]    DispatchPlugin_logic_candidates_0_ctx_hm_GSharePlugin_GSHARE_COUNTER_0;
  wire       [1:0]    DispatchPlugin_logic_candidates_0_ctx_hm_GSharePlugin_GSHARE_COUNTER_1;
  wire       [1:0]    DispatchPlugin_logic_candidates_0_ctx_hm_GSharePlugin_GSHARE_COUNTER_2;
  wire       [1:0]    DispatchPlugin_logic_candidates_0_ctx_hm_GSharePlugin_GSHARE_COUNTER_3;
  wire       [11:0]   DispatchPlugin_logic_candidates_0_ctx_hm_Prediction_BRANCH_HISTORY;
  wire                DispatchPlugin_logic_candidates_0_ctx_hm_DispatchPlugin_FENCE_OLDER;
  wire                DispatchPlugin_logic_candidates_0_ctx_hm_DispatchPlugin_MAY_FLUSH;
  wire                DispatchPlugin_logic_candidates_0_ctx_hm_DispatchPlugin_DONT_FLUSH;
  wire                DispatchPlugin_logic_candidates_0_ctx_hm_DispatchPlugin_DONT_FLUSH_FROM_LANES;
  wire       [0:0]    DispatchPlugin_logic_candidates_0_ctx_hm_Decode_INSTRUCTION_SLICE_COUNT;
  wire                DispatchPlugin_logic_candidates_0_ctx_hm_DONT_FLUSH_PRECISE_3;
  wire                DispatchPlugin_logic_candidates_0_ctx_hm_DONT_FLUSH_PRECISE_4;
  wire       [31:0]   DispatchPlugin_logic_candidates_0_ctx_hm_PC;
  wire                DispatchPlugin_logic_candidates_0_ctx_hm_TRAP;
  wire       [15:0]   DispatchPlugin_logic_candidates_0_ctx_hm_Decode_UOP_ID;
  wire                DispatchPlugin_logic_candidates_0_ctx_hm_RS1_ENABLE;
  wire       [4:0]    DispatchPlugin_logic_candidates_0_ctx_hm_RS1_PHYS;
  wire                DispatchPlugin_logic_candidates_0_ctx_hm_RS2_ENABLE;
  wire       [4:0]    DispatchPlugin_logic_candidates_0_ctx_hm_RS2_PHYS;
  wire                DispatchPlugin_logic_candidates_0_ctx_hm_RD_ENABLE;
  wire       [4:0]    DispatchPlugin_logic_candidates_0_ctx_hm_RD_PHYS;
  wire                DispatchPlugin_logic_candidates_0_ctx_hm_DispatchPlugin_logic_hcs_0_onRs_0_ENABLES_0;
  wire                DispatchPlugin_logic_candidates_0_ctx_hm_DispatchPlugin_logic_hcs_0_onRs_1_ENABLES_0;
  wire                DispatchPlugin_logic_candidates_0_ctx_hm_DispatchPlugin_logic_hcs_1_onRs_0_ENABLES_0;
  wire                DispatchPlugin_logic_candidates_0_ctx_hm_DispatchPlugin_logic_hcs_1_onRs_1_ENABLES_0;
  wire                DispatchPlugin_logic_candidates_0_ctx_hm_DispatchPlugin_logic_hcs_1_onRs_1_ENABLES_1;
  wire                DispatchPlugin_logic_candidates_0_ctx_hm_DispatchPlugin_logic_hcs_2_onRs_0_ENABLES_0;
  wire                DispatchPlugin_logic_candidates_0_ctx_hm_DispatchPlugin_logic_hcs_2_onRs_1_ENABLES_0;
  wire                DispatchPlugin_logic_candidates_0_ctx_hm_DispatchPlugin_logic_hcs_3_onRs_0_ENABLES_0;
  wire                DispatchPlugin_logic_candidates_0_ctx_hm_DispatchPlugin_logic_hcs_3_onRs_1_ENABLES_0;
  wire                DispatchPlugin_logic_candidates_0_fire;
  wire                DispatchPlugin_logic_candidates_0_cancel;
  reg        [3:0]    DispatchPlugin_logic_candidates_0_rsHazards;
  reg        [3:0]    DispatchPlugin_logic_candidates_0_reservationHazards;
  wire                DispatchPlugin_logic_candidates_0_flushHazards;
  wire                DispatchPlugin_logic_candidates_0_fenceOlderHazards;
  wire       [0:0]    DispatchPlugin_logic_candidates_0_age;
  wire                DispatchPlugin_logic_candidates_0_moving;
  wire                DispatchPlugin_logic_candidates_1_ctx_valid;
  reg        [3:0]    DispatchPlugin_logic_candidates_1_ctx_laneLayerHits;
  wire       [31:0]   DispatchPlugin_logic_candidates_1_ctx_uop;
  wire                DispatchPlugin_logic_candidates_1_ctx_hm_Prediction_ALIGNED_JUMPED;
  wire       [31:0]   DispatchPlugin_logic_candidates_1_ctx_hm_Prediction_ALIGNED_JUMPED_PC;
  wire       [3:0]    DispatchPlugin_logic_candidates_1_ctx_hm_Prediction_ALIGNED_SLICES_TAKEN;
  wire       [3:0]    DispatchPlugin_logic_candidates_1_ctx_hm_Prediction_ALIGNED_SLICES_BRANCH;
  wire       [1:0]    DispatchPlugin_logic_candidates_1_ctx_hm_GSharePlugin_GSHARE_COUNTER_0;
  wire       [1:0]    DispatchPlugin_logic_candidates_1_ctx_hm_GSharePlugin_GSHARE_COUNTER_1;
  wire       [1:0]    DispatchPlugin_logic_candidates_1_ctx_hm_GSharePlugin_GSHARE_COUNTER_2;
  wire       [1:0]    DispatchPlugin_logic_candidates_1_ctx_hm_GSharePlugin_GSHARE_COUNTER_3;
  wire       [11:0]   DispatchPlugin_logic_candidates_1_ctx_hm_Prediction_BRANCH_HISTORY;
  wire                DispatchPlugin_logic_candidates_1_ctx_hm_DispatchPlugin_FENCE_OLDER;
  wire                DispatchPlugin_logic_candidates_1_ctx_hm_DispatchPlugin_MAY_FLUSH;
  wire                DispatchPlugin_logic_candidates_1_ctx_hm_DispatchPlugin_DONT_FLUSH;
  wire                DispatchPlugin_logic_candidates_1_ctx_hm_DispatchPlugin_DONT_FLUSH_FROM_LANES;
  wire       [0:0]    DispatchPlugin_logic_candidates_1_ctx_hm_Decode_INSTRUCTION_SLICE_COUNT;
  wire                DispatchPlugin_logic_candidates_1_ctx_hm_DONT_FLUSH_PRECISE_3;
  wire                DispatchPlugin_logic_candidates_1_ctx_hm_DONT_FLUSH_PRECISE_4;
  wire       [31:0]   DispatchPlugin_logic_candidates_1_ctx_hm_PC;
  wire                DispatchPlugin_logic_candidates_1_ctx_hm_TRAP;
  wire       [15:0]   DispatchPlugin_logic_candidates_1_ctx_hm_Decode_UOP_ID;
  wire                DispatchPlugin_logic_candidates_1_ctx_hm_RS1_ENABLE;
  wire       [4:0]    DispatchPlugin_logic_candidates_1_ctx_hm_RS1_PHYS;
  wire                DispatchPlugin_logic_candidates_1_ctx_hm_RS2_ENABLE;
  wire       [4:0]    DispatchPlugin_logic_candidates_1_ctx_hm_RS2_PHYS;
  wire                DispatchPlugin_logic_candidates_1_ctx_hm_RD_ENABLE;
  wire       [4:0]    DispatchPlugin_logic_candidates_1_ctx_hm_RD_PHYS;
  wire                DispatchPlugin_logic_candidates_1_ctx_hm_DispatchPlugin_logic_hcs_0_onRs_0_ENABLES_0;
  wire                DispatchPlugin_logic_candidates_1_ctx_hm_DispatchPlugin_logic_hcs_0_onRs_1_ENABLES_0;
  wire                DispatchPlugin_logic_candidates_1_ctx_hm_DispatchPlugin_logic_hcs_1_onRs_0_ENABLES_0;
  wire                DispatchPlugin_logic_candidates_1_ctx_hm_DispatchPlugin_logic_hcs_1_onRs_1_ENABLES_0;
  wire                DispatchPlugin_logic_candidates_1_ctx_hm_DispatchPlugin_logic_hcs_1_onRs_1_ENABLES_1;
  wire                DispatchPlugin_logic_candidates_1_ctx_hm_DispatchPlugin_logic_hcs_2_onRs_0_ENABLES_0;
  wire                DispatchPlugin_logic_candidates_1_ctx_hm_DispatchPlugin_logic_hcs_2_onRs_1_ENABLES_0;
  wire                DispatchPlugin_logic_candidates_1_ctx_hm_DispatchPlugin_logic_hcs_3_onRs_0_ENABLES_0;
  wire                DispatchPlugin_logic_candidates_1_ctx_hm_DispatchPlugin_logic_hcs_3_onRs_1_ENABLES_0;
  wire                DispatchPlugin_logic_candidates_1_fire;
  wire                DispatchPlugin_logic_candidates_1_cancel;
  reg        [3:0]    DispatchPlugin_logic_candidates_1_rsHazards;
  reg        [3:0]    DispatchPlugin_logic_candidates_1_reservationHazards;
  wire                DispatchPlugin_logic_candidates_1_flushHazards;
  wire                DispatchPlugin_logic_candidates_1_fenceOlderHazards;
  wire       [0:0]    DispatchPlugin_logic_candidates_1_age;
  wire                DispatchPlugin_logic_candidates_1_moving;
  wire                DispatchPlugin_logic_candidates_2_ctx_valid;
  reg        [3:0]    DispatchPlugin_logic_candidates_2_ctx_laneLayerHits;
  wire       [31:0]   DispatchPlugin_logic_candidates_2_ctx_uop;
  wire                DispatchPlugin_logic_candidates_2_ctx_hm_Prediction_ALIGNED_JUMPED;
  wire       [31:0]   DispatchPlugin_logic_candidates_2_ctx_hm_Prediction_ALIGNED_JUMPED_PC;
  wire       [3:0]    DispatchPlugin_logic_candidates_2_ctx_hm_Prediction_ALIGNED_SLICES_TAKEN;
  wire       [3:0]    DispatchPlugin_logic_candidates_2_ctx_hm_Prediction_ALIGNED_SLICES_BRANCH;
  wire       [1:0]    DispatchPlugin_logic_candidates_2_ctx_hm_GSharePlugin_GSHARE_COUNTER_0;
  wire       [1:0]    DispatchPlugin_logic_candidates_2_ctx_hm_GSharePlugin_GSHARE_COUNTER_1;
  wire       [1:0]    DispatchPlugin_logic_candidates_2_ctx_hm_GSharePlugin_GSHARE_COUNTER_2;
  wire       [1:0]    DispatchPlugin_logic_candidates_2_ctx_hm_GSharePlugin_GSHARE_COUNTER_3;
  wire       [11:0]   DispatchPlugin_logic_candidates_2_ctx_hm_Prediction_BRANCH_HISTORY;
  wire                DispatchPlugin_logic_candidates_2_ctx_hm_DispatchPlugin_FENCE_OLDER;
  wire                DispatchPlugin_logic_candidates_2_ctx_hm_DispatchPlugin_MAY_FLUSH;
  wire                DispatchPlugin_logic_candidates_2_ctx_hm_DispatchPlugin_DONT_FLUSH;
  wire                DispatchPlugin_logic_candidates_2_ctx_hm_DispatchPlugin_DONT_FLUSH_FROM_LANES;
  wire       [0:0]    DispatchPlugin_logic_candidates_2_ctx_hm_Decode_INSTRUCTION_SLICE_COUNT;
  wire                DispatchPlugin_logic_candidates_2_ctx_hm_DONT_FLUSH_PRECISE_3;
  wire                DispatchPlugin_logic_candidates_2_ctx_hm_DONT_FLUSH_PRECISE_4;
  wire       [31:0]   DispatchPlugin_logic_candidates_2_ctx_hm_PC;
  wire                DispatchPlugin_logic_candidates_2_ctx_hm_TRAP;
  wire       [15:0]   DispatchPlugin_logic_candidates_2_ctx_hm_Decode_UOP_ID;
  wire                DispatchPlugin_logic_candidates_2_ctx_hm_RS1_ENABLE;
  wire       [4:0]    DispatchPlugin_logic_candidates_2_ctx_hm_RS1_PHYS;
  wire                DispatchPlugin_logic_candidates_2_ctx_hm_RS2_ENABLE;
  wire       [4:0]    DispatchPlugin_logic_candidates_2_ctx_hm_RS2_PHYS;
  wire                DispatchPlugin_logic_candidates_2_ctx_hm_RD_ENABLE;
  wire       [4:0]    DispatchPlugin_logic_candidates_2_ctx_hm_RD_PHYS;
  wire                DispatchPlugin_logic_candidates_2_ctx_hm_DispatchPlugin_logic_hcs_0_onRs_0_ENABLES_0;
  wire                DispatchPlugin_logic_candidates_2_ctx_hm_DispatchPlugin_logic_hcs_0_onRs_1_ENABLES_0;
  wire                DispatchPlugin_logic_candidates_2_ctx_hm_DispatchPlugin_logic_hcs_1_onRs_0_ENABLES_0;
  wire                DispatchPlugin_logic_candidates_2_ctx_hm_DispatchPlugin_logic_hcs_1_onRs_1_ENABLES_0;
  wire                DispatchPlugin_logic_candidates_2_ctx_hm_DispatchPlugin_logic_hcs_1_onRs_1_ENABLES_1;
  wire                DispatchPlugin_logic_candidates_2_ctx_hm_DispatchPlugin_logic_hcs_2_onRs_0_ENABLES_0;
  wire                DispatchPlugin_logic_candidates_2_ctx_hm_DispatchPlugin_logic_hcs_2_onRs_1_ENABLES_0;
  wire                DispatchPlugin_logic_candidates_2_ctx_hm_DispatchPlugin_logic_hcs_3_onRs_0_ENABLES_0;
  wire                DispatchPlugin_logic_candidates_2_ctx_hm_DispatchPlugin_logic_hcs_3_onRs_1_ENABLES_0;
  wire                DispatchPlugin_logic_candidates_2_fire;
  wire                DispatchPlugin_logic_candidates_2_cancel;
  reg        [3:0]    DispatchPlugin_logic_candidates_2_rsHazards;
  reg        [3:0]    DispatchPlugin_logic_candidates_2_reservationHazards;
  wire                DispatchPlugin_logic_candidates_2_flushHazards;
  wire                DispatchPlugin_logic_candidates_2_fenceOlderHazards;
  wire       [0:0]    DispatchPlugin_logic_candidates_2_age;
  wire                DispatchPlugin_logic_candidates_2_moving;
  wire                DispatchPlugin_logic_rsHazardChecker_0_onLl_0_onRs_0_hazard;
  wire                DispatchPlugin_logic_rsHazardChecker_0_onLl_0_onRs_1_hazard;
  wire                DispatchPlugin_logic_rsHazardChecker_0_onLl_1_onRs_0_hazard;
  wire                DispatchPlugin_logic_rsHazardChecker_0_onLl_1_onRs_1_hazard;
  wire                DispatchPlugin_logic_rsHazardChecker_0_onLl_2_onRs_0_hazard;
  wire                DispatchPlugin_logic_rsHazardChecker_0_onLl_2_onRs_1_hazard;
  wire                DispatchPlugin_logic_rsHazardChecker_0_onLl_3_onRs_0_hazard;
  wire                DispatchPlugin_logic_rsHazardChecker_0_onLl_3_onRs_1_hazard;
  wire                DispatchPlugin_logic_rsHazardChecker_1_onLl_0_onRs_0_hazard;
  wire                DispatchPlugin_logic_rsHazardChecker_1_onLl_0_onRs_1_hazard;
  wire                DispatchPlugin_logic_rsHazardChecker_1_onLl_1_onRs_0_hazard;
  wire                DispatchPlugin_logic_rsHazardChecker_1_onLl_1_onRs_1_hazard;
  wire                DispatchPlugin_logic_rsHazardChecker_1_onLl_2_onRs_0_hazard;
  wire                DispatchPlugin_logic_rsHazardChecker_1_onLl_2_onRs_1_hazard;
  wire                DispatchPlugin_logic_rsHazardChecker_1_onLl_3_onRs_0_hazard;
  wire                DispatchPlugin_logic_rsHazardChecker_1_onLl_3_onRs_1_hazard;
  wire                DispatchPlugin_logic_rsHazardChecker_2_onLl_0_onRs_0_hazard;
  wire                DispatchPlugin_logic_rsHazardChecker_2_onLl_0_onRs_1_hazard;
  wire                DispatchPlugin_logic_rsHazardChecker_2_onLl_1_onRs_0_hazard;
  wire                DispatchPlugin_logic_rsHazardChecker_2_onLl_1_onRs_1_hazard;
  wire                DispatchPlugin_logic_rsHazardChecker_2_onLl_2_onRs_0_hazard;
  wire                DispatchPlugin_logic_rsHazardChecker_2_onLl_2_onRs_1_hazard;
  wire                DispatchPlugin_logic_rsHazardChecker_2_onLl_3_onRs_0_hazard;
  wire                DispatchPlugin_logic_rsHazardChecker_2_onLl_3_onRs_1_hazard;
  wire                DispatchPlugin_logic_reservationChecker_0_onLl_0_hit;
  wire                DispatchPlugin_logic_reservationChecker_0_onLl_1_hit;
  wire                DispatchPlugin_logic_reservationChecker_0_onLl_2_hit;
  wire                DispatchPlugin_logic_reservationChecker_0_onLl_3_hit;
  wire                DispatchPlugin_logic_reservationChecker_1_onLl_0_hit;
  wire                DispatchPlugin_logic_reservationChecker_1_onLl_1_hit;
  wire                DispatchPlugin_logic_reservationChecker_1_onLl_2_hit;
  wire                DispatchPlugin_logic_reservationChecker_1_onLl_3_hit;
  wire                DispatchPlugin_logic_reservationChecker_2_onLl_0_hit;
  wire                DispatchPlugin_logic_reservationChecker_2_onLl_1_hit;
  wire                DispatchPlugin_logic_reservationChecker_2_onLl_2_hit;
  wire                DispatchPlugin_logic_reservationChecker_2_onLl_3_hit;
  wire                DispatchPlugin_logic_flushChecker_0_executeCheck_0_hits_0;
  wire                DispatchPlugin_logic_flushChecker_0_executeCheck_0_hits_1;
  wire                DispatchPlugin_logic_flushChecker_0_executeCheck_1_hits_0;
  wire                DispatchPlugin_logic_flushChecker_0_executeCheck_1_hits_1;
  wire                DispatchPlugin_logic_flushChecker_0_oldersHazard;
  wire                DispatchPlugin_logic_flushChecker_1_executeCheck_0_hits_0;
  wire                DispatchPlugin_logic_flushChecker_1_executeCheck_0_hits_1;
  wire                DispatchPlugin_logic_flushChecker_1_executeCheck_1_hits_0;
  wire                DispatchPlugin_logic_flushChecker_1_executeCheck_1_hits_1;
  wire                DispatchPlugin_logic_flushChecker_1_oldersHazard;
  wire                DispatchPlugin_logic_flushChecker_2_executeCheck_0_hits_0;
  wire                DispatchPlugin_logic_flushChecker_2_executeCheck_0_hits_1;
  wire                DispatchPlugin_logic_flushChecker_2_executeCheck_1_hits_0;
  wire                DispatchPlugin_logic_flushChecker_2_executeCheck_1_hits_1;
  wire                DispatchPlugin_logic_flushChecker_2_oldersHazard;
  wire       [0:0]    DispatchPlugin_logic_fenceChecker_olderInflights;
  wire                DispatchPlugin_logic_feeds_0_sending;
  reg                 DispatchPlugin_logic_feeds_0_sent;
  wire                when_DispatchPlugin_l358;
  wire                DispatchPlugin_logic_feeds_1_sending;
  reg                 DispatchPlugin_logic_feeds_1_sent;
  wire                when_DispatchPlugin_l358_1;
  wire                when_DispatchPlugin_l368;
  wire                _zz_toplevel_decode_ctrls_1_down_DispatchPlugin_logic_LANES_LAYER_HIT_3_0_1;
  wire                _zz_toplevel_decode_ctrls_1_down_DispatchPlugin_logic_LANES_LAYER_HIT_3_0_2;
  wire                _zz_toplevel_decode_ctrls_1_down_DispatchPlugin_logic_hcs_3_onRs_1_ENABLES_0_0;
  wire                _zz_toplevel_decode_ctrls_1_down_DispatchPlugin_logic_LANES_LAYER_HIT_3_0_3;
  wire                _zz_toplevel_decode_ctrls_1_down_DispatchPlugin_logic_LANES_LAYER_HIT_3_0_4;
  wire                _zz_toplevel_decode_ctrls_1_down_DispatchPlugin_logic_hcs_1_onRs_1_ENABLES_0_0;
  wire                _zz_toplevel_decode_ctrls_1_down_DONT_FLUSH_PRECISE_4_0;
  wire                _zz_toplevel_decode_ctrls_1_down_DONT_FLUSH_PRECISE_4_0_1;
  wire                _zz_toplevel_decode_ctrls_1_down_DispatchPlugin_logic_LANES_LAYER_HIT_3_1_1;
  wire                _zz_toplevel_decode_ctrls_1_down_DispatchPlugin_logic_LANES_LAYER_HIT_3_1_2;
  wire                _zz_toplevel_decode_ctrls_1_down_DispatchPlugin_logic_hcs_3_onRs_1_ENABLES_0_1;
  wire                _zz_toplevel_decode_ctrls_1_down_DispatchPlugin_logic_LANES_LAYER_HIT_3_1_3;
  wire                _zz_toplevel_decode_ctrls_1_down_DispatchPlugin_logic_LANES_LAYER_HIT_3_1_4;
  wire                _zz_toplevel_decode_ctrls_1_down_DispatchPlugin_logic_hcs_1_onRs_1_ENABLES_0_1;
  wire                _zz_toplevel_decode_ctrls_1_down_DONT_FLUSH_PRECISE_4_1;
  wire                _zz_toplevel_decode_ctrls_1_down_DONT_FLUSH_PRECISE_4_1_1;
  wire                TrapPlugin_logic_initHold;
  reg                 toplevel_decode_ctrls_1_up_LANE_SEL_0_regNext_1;
  wire                when_CtrlLaneApi_l46_4;
  wire                WhiteboxerPlugin_logic_serializeds_0_fire;
  wire       [9:0]    WhiteboxerPlugin_logic_serializeds_0_decodeId;
  wire       [15:0]   WhiteboxerPlugin_logic_serializeds_0_microOpId;
  wire       [31:0]   WhiteboxerPlugin_logic_serializeds_0_microOp;
  reg                 toplevel_decode_ctrls_1_up_LANE_SEL_1_regNext_1;
  wire                when_CtrlLaneApi_l46_5;
  wire                WhiteboxerPlugin_logic_serializeds_1_fire;
  wire       [9:0]    WhiteboxerPlugin_logic_serializeds_1_decodeId;
  wire       [15:0]   WhiteboxerPlugin_logic_serializeds_1_microOpId;
  wire       [31:0]   WhiteboxerPlugin_logic_serializeds_1_microOp;
  reg                 toplevel_execute_ctrl0_down_LANE_SEL_lane0_regNext;
  wire                when_CtrlLaneApi_l46_6;
  wire                WhiteboxerPlugin_logic_dispatches_0_fire;
  wire       [15:0]   WhiteboxerPlugin_logic_dispatches_0_microOpId;
  wire                toplevel_execute_lane1_ctrls_0_upIsCancel;
  wire                toplevel_execute_lane1_ctrls_0_downIsCancel;
  reg                 toplevel_execute_ctrl0_down_LANE_SEL_lane1_regNext;
  wire                when_CtrlLaneApi_l46_7;
  wire                WhiteboxerPlugin_logic_dispatches_1_fire;
  wire       [15:0]   WhiteboxerPlugin_logic_dispatches_1_microOpId;
  reg                 toplevel_execute_ctrl2_down_LANE_SEL_lane0_regNext;
  wire                when_CtrlLaneApi_l46_8;
  wire                WhiteboxerPlugin_logic_executes_0_fire;
  wire       [15:0]   WhiteboxerPlugin_logic_executes_0_microOpId;
  reg                 toplevel_execute_ctrl2_down_LANE_SEL_lane1_regNext;
  wire                when_CtrlLaneApi_l46_9;
  wire                WhiteboxerPlugin_logic_executes_1_fire;
  wire       [15:0]   WhiteboxerPlugin_logic_executes_1_microOpId;
  wire                WhiteboxerPlugin_logic_csr_access_valid;
  wire       [15:0]   WhiteboxerPlugin_logic_csr_access_payload_uopId;
  wire       [11:0]   WhiteboxerPlugin_logic_csr_access_payload_address;
  wire       [31:0]   WhiteboxerPlugin_logic_csr_access_payload_write;
  wire       [31:0]   WhiteboxerPlugin_logic_csr_access_payload_read;
  wire                WhiteboxerPlugin_logic_csr_access_payload_writeDone;
  wire                WhiteboxerPlugin_logic_csr_access_payload_readDone;
  wire       [15:0]   BtbPlugin_logic_onForget_hash;
  wire                BtbPlugin_logic_readPort_cmd_valid;
  wire       [7:0]    BtbPlugin_logic_readPort_cmd_payload;
  wire       [15:0]   BtbPlugin_logic_readPort_rsp_0_hash;
  wire       [0:0]    BtbPlugin_logic_readPort_rsp_0_sliceLow;
  wire       [30:0]   BtbPlugin_logic_readPort_rsp_0_pcTarget;
  wire                BtbPlugin_logic_readPort_rsp_0_isBranch;
  wire                BtbPlugin_logic_readPort_rsp_0_isPush;
  wire                BtbPlugin_logic_readPort_rsp_0_isPop;
  wire       [15:0]   BtbPlugin_logic_readPort_rsp_1_hash;
  wire       [0:0]    BtbPlugin_logic_readPort_rsp_1_sliceLow;
  wire       [30:0]   BtbPlugin_logic_readPort_rsp_1_pcTarget;
  wire                BtbPlugin_logic_readPort_rsp_1_isBranch;
  wire                BtbPlugin_logic_readPort_rsp_1_isPush;
  wire                BtbPlugin_logic_readPort_rsp_1_isPop;
  wire       [101:0]  _zz_BtbPlugin_logic_readPort_rsp_0_hash;
  wire       [50:0]   _zz_BtbPlugin_logic_readPort_rsp_0_hash_1;
  wire       [50:0]   _zz_BtbPlugin_logic_readPort_rsp_1_hash;
  wire                fetch_logic_ctrls_0_haltRequest_BtbPlugin_l171;
  wire       [3:0]    BtbPlugin_logic_predictions;
  wire       [1:0]    BtbPlugin_logic_applyIt_chunksMask;
  wire       [1:0]    BtbPlugin_logic_applyIt_chunksTakenOh;
  wire                BtbPlugin_logic_applyIt_needIt;
  reg                 BtbPlugin_logic_applyIt_correctionSent;
  wire                when_BtbPlugin_l205;
  wire                BtbPlugin_logic_applyIt_doIt;
  wire                _zz_BtbPlugin_logic_applyIt_doItSlice;
  wire       [15:0]   BtbPlugin_logic_applyIt_entry_hash;
  wire       [0:0]    BtbPlugin_logic_applyIt_entry_sliceLow;
  wire       [30:0]   BtbPlugin_logic_applyIt_entry_pcTarget;
  wire                BtbPlugin_logic_applyIt_entry_isBranch;
  wire                BtbPlugin_logic_applyIt_entry_isPush;
  wire                BtbPlugin_logic_applyIt_entry_isPop;
  wire       [50:0]   _zz_BtbPlugin_logic_applyIt_entry_hash;
  reg        [30:0]   BtbPlugin_logic_applyIt_pcTarget;
  wire       [1:0]    BtbPlugin_logic_applyIt_doItSlice;
  wire                BtbPlugin_logic_applyIt_rasLogic_pushValid;
  reg        [31:0]   BtbPlugin_logic_applyIt_rasLogic_pushPc;
  wire                when_BtbPlugin_l218;
  wire       [11:0]   BtbPlugin_logic_applyIt_history_layers_0_history;
  wire                BtbPlugin_logic_applyIt_history_layers_0_valid;
  wire       [11:0]   BtbPlugin_logic_applyIt_history_layers_1_history;
  wire                BtbPlugin_logic_applyIt_history_layers_1_valid;
  wire       [11:0]   BtbPlugin_logic_applyIt_history_layers_2_history;
  wire                BtbPlugin_logic_applyIt_history_layers_2_valid;
  wire                BtbPlugin_logic_applyIt_history_layersLogic_0_doIt;
  wire       [11:0]   BtbPlugin_logic_applyIt_history_layersLogic_0_shifted;
  wire                BtbPlugin_logic_applyIt_history_layersLogic_1_doIt;
  wire       [11:0]   BtbPlugin_logic_applyIt_history_layersLogic_1_shifted;
  reg        [8:0]    BtbPlugin_logic_initializer_counter;
  wire                BtbPlugin_logic_initializer_busy;
  reg                 TrapPlugin_logic_harts_0_crsPorts_read_valid;
  wire                TrapPlugin_logic_harts_0_crsPorts_read_ready;
  reg        [2:0]    TrapPlugin_logic_harts_0_crsPorts_read_address;
  wire       [31:0]   TrapPlugin_logic_harts_0_crsPorts_read_data;
  wire                AlignerPlugin_logic_buffer_flushIt;
  wire                AlignerPlugin_logic_buffer_readers_0_firstFromBuffer;
  wire                AlignerPlugin_logic_buffer_readers_0_lastFromBuffer;
  wire       [7:0]    _zz_AlignerPlugin_logic_extractors_0_ctx_instruction;
  wire                _zz_AlignerPlugin_logic_extractors_0_ctx_pc;
  wire                _zz_AlignerPlugin_logic_extractors_0_ctx_pc_1;
  wire                _zz_AlignerPlugin_logic_extractors_0_ctx_pc_2;
  wire                AlignerPlugin_logic_buffer_readers_1_firstFromBuffer;
  wire                AlignerPlugin_logic_buffer_readers_1_lastFromBuffer;
  wire       [6:0]    _zz_AlignerPlugin_logic_extractors_1_ctx_instruction;
  wire                _zz_AlignerPlugin_logic_extractors_1_ctx_pc;
  wire                _zz_AlignerPlugin_logic_extractors_1_ctx_pc_1;
  wire                _zz_AlignerPlugin_logic_extractors_1_ctx_pc_2;
  wire                DispatchPlugin_logic_slotsFeeds_free;
  wire                DispatchPlugin_logic_slotsFeeds_fit;
  wire                DispatchPlugin_logic_slotsFeeds_doIt;
  wire       [1:0]    _zz_DispatchPlugin_logic_slots_0_ctx_valid;
  wire                _zz_DispatchPlugin_logic_slots_0_ctx_valid_1;
  reg        [1:0]    _zz_DispatchPlugin_logic_slots_0_ctx_valid_2;
  wire       [1:0]    _zz_DispatchPlugin_logic_slots_0_ctx_valid_3;
  wire       [180:0]  _zz_DispatchPlugin_logic_slots_0_ctx_valid_4;
  wire       [143:0]  _zz_DispatchPlugin_logic_slots_0_ctx_hm_Prediction_ALIGNED_JUMPED;
  wire       [7:0]    _zz_DispatchPlugin_logic_slots_0_ctx_hm_GSharePlugin_GSHARE_COUNTER_0;
  wire       [1:0]    DispatchPlugin_logic_scheduler_eusFree_0;
  wire       [1:0]    DispatchPlugin_logic_scheduler_eusFree_1;
  wire       [1:0]    DispatchPlugin_logic_scheduler_eusFree_2;
  wire       [1:0]    DispatchPlugin_logic_scheduler_eusFree_3;
  wire       [0:0]    DispatchPlugin_logic_scheduler_hartFree_0;
  wire       [0:0]    DispatchPlugin_logic_scheduler_hartFree_1;
  wire       [0:0]    DispatchPlugin_logic_scheduler_hartFree_2;
  wire       [0:0]    DispatchPlugin_logic_scheduler_hartFree_3;
  wire                DispatchPlugin_logic_scheduler_arbiters_0_candHazard;
  wire       [3:0]    DispatchPlugin_logic_scheduler_arbiters_0_layersHits;
  wire       [3:0]    _zz_DispatchPlugin_logic_scheduler_arbiters_0_layersHits_bools_0;
  wire                DispatchPlugin_logic_scheduler_arbiters_0_layersHits_bools_0;
  wire                DispatchPlugin_logic_scheduler_arbiters_0_layersHits_bools_1;
  wire                DispatchPlugin_logic_scheduler_arbiters_0_layersHits_bools_2;
  wire                DispatchPlugin_logic_scheduler_arbiters_0_layersHits_bools_3;
  reg        [3:0]    _zz_DispatchPlugin_logic_scheduler_arbiters_0_layerOh;
  wire                DispatchPlugin_logic_scheduler_arbiters_0_layersHits_range_0_to_1;
  wire                DispatchPlugin_logic_scheduler_arbiters_0_layersHits_range_0_to_2;
  wire       [3:0]    DispatchPlugin_logic_scheduler_arbiters_0_layerOh;
  wire       [1:0]    DispatchPlugin_logic_scheduler_arbiters_0_eusOh;
  wire                DispatchPlugin_logic_scheduler_arbiters_0_doIt;
  wire                DispatchPlugin_logic_scheduler_arbiters_1_candHazards_0_doWrite;
  wire                DispatchPlugin_logic_scheduler_arbiters_1_candHazards_0_rfas_0;
  wire                DispatchPlugin_logic_scheduler_arbiters_1_candHazards_0_rfas_1;
  wire                DispatchPlugin_logic_scheduler_arbiters_1_candHazards_0_rfas_2;
  wire                DispatchPlugin_logic_scheduler_arbiters_1_candHazards_0_hit;
  wire                DispatchPlugin_logic_scheduler_arbiters_1_candHazard;
  wire       [3:0]    DispatchPlugin_logic_scheduler_arbiters_1_layersHits;
  wire       [3:0]    _zz_DispatchPlugin_logic_scheduler_arbiters_1_layersHits_bools_0;
  wire                DispatchPlugin_logic_scheduler_arbiters_1_layersHits_bools_0;
  wire                DispatchPlugin_logic_scheduler_arbiters_1_layersHits_bools_1;
  wire                DispatchPlugin_logic_scheduler_arbiters_1_layersHits_bools_2;
  wire                DispatchPlugin_logic_scheduler_arbiters_1_layersHits_bools_3;
  reg        [3:0]    _zz_DispatchPlugin_logic_scheduler_arbiters_1_layerOh;
  wire                DispatchPlugin_logic_scheduler_arbiters_1_layersHits_range_0_to_1;
  wire                DispatchPlugin_logic_scheduler_arbiters_1_layersHits_range_0_to_2;
  wire       [3:0]    DispatchPlugin_logic_scheduler_arbiters_1_layerOh;
  wire       [1:0]    DispatchPlugin_logic_scheduler_arbiters_1_eusOh;
  wire                DispatchPlugin_logic_scheduler_arbiters_1_doIt;
  wire                DispatchPlugin_logic_scheduler_arbiters_2_candHazards_0_doWrite;
  wire                DispatchPlugin_logic_scheduler_arbiters_2_candHazards_0_rfas_0;
  wire                DispatchPlugin_logic_scheduler_arbiters_2_candHazards_0_rfas_1;
  wire                DispatchPlugin_logic_scheduler_arbiters_2_candHazards_0_rfas_2;
  wire                DispatchPlugin_logic_scheduler_arbiters_2_candHazards_0_hit;
  wire                DispatchPlugin_logic_scheduler_arbiters_2_candHazards_1_doWrite;
  wire                DispatchPlugin_logic_scheduler_arbiters_2_candHazards_1_rfas_0;
  wire                DispatchPlugin_logic_scheduler_arbiters_2_candHazards_1_rfas_1;
  wire                DispatchPlugin_logic_scheduler_arbiters_2_candHazards_1_rfas_2;
  wire                DispatchPlugin_logic_scheduler_arbiters_2_candHazards_1_hit;
  wire                DispatchPlugin_logic_scheduler_arbiters_2_candHazard;
  wire       [3:0]    DispatchPlugin_logic_scheduler_arbiters_2_layersHits;
  wire       [3:0]    _zz_DispatchPlugin_logic_scheduler_arbiters_2_layersHits_bools_0;
  wire                DispatchPlugin_logic_scheduler_arbiters_2_layersHits_bools_0;
  wire                DispatchPlugin_logic_scheduler_arbiters_2_layersHits_bools_1;
  wire                DispatchPlugin_logic_scheduler_arbiters_2_layersHits_bools_2;
  wire                DispatchPlugin_logic_scheduler_arbiters_2_layersHits_bools_3;
  reg        [3:0]    _zz_DispatchPlugin_logic_scheduler_arbiters_2_layerOh;
  wire                DispatchPlugin_logic_scheduler_arbiters_2_layersHits_range_0_to_1;
  wire                DispatchPlugin_logic_scheduler_arbiters_2_layersHits_range_0_to_2;
  wire       [3:0]    DispatchPlugin_logic_scheduler_arbiters_2_layerOh;
  wire       [1:0]    DispatchPlugin_logic_scheduler_arbiters_2_eusOh;
  wire                DispatchPlugin_logic_scheduler_arbiters_2_doIt;
  wire       [2:0]    DispatchPlugin_logic_inserter_0_oh;
  wire                _zz_toplevel_execute_ctrl0_up_LANE_AGE_lane0;
  wire                _zz_toplevel_execute_ctrl0_up_LANE_AGE_lane0_1;
  wire                _zz_toplevel_execute_ctrl0_up_LANE_AGE_lane0_2;
  wire                DispatchPlugin_logic_inserter_0_trap;
  wire       [7:0]    _zz_toplevel_execute_ctrl0_up_GSharePlugin_GSHARE_COUNTER_lane0_0;
  wire                when_DispatchPlugin_l427;
  wire       [3:0]    DispatchPlugin_logic_inserter_0_layerOhUnfiltred;
  wire       [0:0]    DispatchPlugin_logic_inserter_0_layer_0_0;
  wire                DispatchPlugin_logic_inserter_0_layer_0_1;
  wire       [0:0]    DispatchPlugin_logic_inserter_0_layer_1_0;
  wire                DispatchPlugin_logic_inserter_0_layer_1_1;
  wire       [1:0]    _zz_toplevel_execute_ctrl0_up_execute_lane0_LAYER_SEL_lane0;
  wire       [2:0]    DispatchPlugin_logic_inserter_1_oh;
  wire                _zz_toplevel_execute_ctrl0_up_LANE_AGE_lane1;
  wire                _zz_toplevel_execute_ctrl0_up_LANE_AGE_lane1_1;
  wire                _zz_toplevel_execute_ctrl0_up_LANE_AGE_lane1_2;
  wire                DispatchPlugin_logic_inserter_1_trap;
  wire       [7:0]    _zz_toplevel_execute_ctrl0_up_GSharePlugin_GSHARE_COUNTER_lane1_0;
  wire                when_DispatchPlugin_l427_1;
  wire       [3:0]    DispatchPlugin_logic_inserter_1_layerOhUnfiltred;
  wire       [0:0]    DispatchPlugin_logic_inserter_1_layer_0_0;
  wire                DispatchPlugin_logic_inserter_1_layer_0_1;
  wire       [0:0]    DispatchPlugin_logic_inserter_1_layer_1_0;
  wire                DispatchPlugin_logic_inserter_1_layer_1_1;
  wire       [1:0]    _zz_toplevel_execute_ctrl0_up_execute_lane1_LAYER_SEL_lane1;
  wire                decode_logic_flushes_0_onLanes_0_doIt;
  wire                decode_logic_flushes_0_onLanes_1_doIt;
  wire                decode_logic_flushes_1_onLanes_0_doIt;
  wire       [0:0]    _zz_decode_logic_flushes_1_onLanes_1_doIt;
  wire                decode_logic_flushes_1_onLanes_1_doIt;
  wire                toplevel_execute_lane1_bypasser_integer_RS1_port_valid;
  wire       [4:0]    toplevel_execute_lane1_bypasser_integer_RS1_port_address;
  wire       [31:0]   toplevel_execute_lane1_bypasser_integer_RS1_port_data;
  wire                LsuL1Plugin_logic_bus_read_cmd_valid;
  wire                LsuL1Plugin_logic_bus_read_cmd_ready;
  wire       [31:0]   LsuL1Plugin_logic_bus_read_cmd_payload_address;
  wire                LsuL1Plugin_logic_bus_read_rsp_valid;
  wire                LsuL1Plugin_logic_bus_read_rsp_ready;
  wire       [63:0]   LsuL1Plugin_logic_bus_read_rsp_payload_data;
  wire                LsuL1Plugin_logic_bus_read_rsp_payload_error;
  wire                LsuL1Plugin_logic_bus_write_cmd_valid;
  wire                LsuL1Plugin_logic_bus_write_cmd_ready;
  wire                LsuL1Plugin_logic_bus_write_cmd_payload_last;
  wire       [31:0]   LsuL1Plugin_logic_bus_write_cmd_payload_fragment_address;
  wire       [63:0]   LsuL1Plugin_logic_bus_write_cmd_payload_fragment_data;
  wire                LsuL1Plugin_logic_bus_write_rsp_valid;
  wire                LsuL1Plugin_logic_bus_write_rsp_payload_error;
  reg        [0:0]    LsuL1Plugin_logic_refillCompletions;
  wire                LsuL1Plugin_logic_writebackBusy;
  reg        [1:0]    LsuL1Plugin_logic_banksWrite_mask;
  reg        [8:0]    LsuL1Plugin_logic_banksWrite_address;
  reg        [63:0]   LsuL1Plugin_logic_banksWrite_writeData;
  reg        [7:0]    LsuL1Plugin_logic_banksWrite_writeMask;
  reg        [1:0]    LsuL1Plugin_logic_waysWrite_mask;
  reg        [5:0]    LsuL1Plugin_logic_waysWrite_address;
  reg                 LsuL1Plugin_logic_waysWrite_tag_loaded;
  reg        [19:0]   LsuL1Plugin_logic_waysWrite_tag_address;
  reg                 LsuL1Plugin_logic_waysWrite_tag_fault;
  wire                LsuL1Plugin_logic_waysWrite_valid;
  wire                LsuL1Plugin_logic_banks_0_usedByWriteback;
  wire                LsuL1Plugin_logic_banks_0_write_valid;
  wire       [8:0]    LsuL1Plugin_logic_banks_0_write_payload_address;
  wire       [63:0]   LsuL1Plugin_logic_banks_0_write_payload_data;
  wire       [7:0]    LsuL1Plugin_logic_banks_0_write_payload_mask;
  reg                 LsuL1Plugin_logic_banks_0_read_cmd_valid;
  reg        [8:0]    LsuL1Plugin_logic_banks_0_read_cmd_payload;
  (* keep , syn_keep *) wire       [63:0]   LsuL1Plugin_logic_banks_0_read_rsp /* synthesis syn_keep = 1 */ ;
  wire                LsuL1Plugin_logic_banks_1_usedByWriteback;
  wire                LsuL1Plugin_logic_banks_1_write_valid;
  wire       [8:0]    LsuL1Plugin_logic_banks_1_write_payload_address;
  wire       [63:0]   LsuL1Plugin_logic_banks_1_write_payload_data;
  wire       [7:0]    LsuL1Plugin_logic_banks_1_write_payload_mask;
  reg                 LsuL1Plugin_logic_banks_1_read_cmd_valid;
  reg        [8:0]    LsuL1Plugin_logic_banks_1_read_cmd_payload;
  (* keep , syn_keep *) wire       [63:0]   LsuL1Plugin_logic_banks_1_read_rsp /* synthesis syn_keep = 1 */ ;
  wire                LsuL1Plugin_logic_ways_0_lsuRead_cmd_valid;
  wire       [5:0]    LsuL1Plugin_logic_ways_0_lsuRead_cmd_payload;
  (* keep , syn_keep *) wire                LsuL1Plugin_logic_ways_0_lsuRead_rsp_loaded /* synthesis syn_keep = 1 */ ;
  (* keep , syn_keep *) wire       [19:0]   LsuL1Plugin_logic_ways_0_lsuRead_rsp_address /* synthesis syn_keep = 1 */ ;
  (* keep , syn_keep *) wire                LsuL1Plugin_logic_ways_0_lsuRead_rsp_fault /* synthesis syn_keep = 1 */ ;
  wire       [21:0]   _zz_LsuL1Plugin_logic_ways_0_lsuRead_rsp_loaded;
  wire                LsuL1Plugin_logic_ways_1_lsuRead_cmd_valid;
  wire       [5:0]    LsuL1Plugin_logic_ways_1_lsuRead_cmd_payload;
  (* keep , syn_keep *) wire                LsuL1Plugin_logic_ways_1_lsuRead_rsp_loaded /* synthesis syn_keep = 1 */ ;
  (* keep , syn_keep *) wire       [19:0]   LsuL1Plugin_logic_ways_1_lsuRead_rsp_address /* synthesis syn_keep = 1 */ ;
  (* keep , syn_keep *) wire                LsuL1Plugin_logic_ways_1_lsuRead_rsp_fault /* synthesis syn_keep = 1 */ ;
  wire       [21:0]   _zz_LsuL1Plugin_logic_ways_1_lsuRead_rsp_loaded;
  reg                 LsuL1Plugin_logic_shared_write_valid;
  reg        [5:0]    LsuL1Plugin_logic_shared_write_payload_address;
  reg        [0:0]    LsuL1Plugin_logic_shared_write_payload_data_plru_0;
  reg        [1:0]    LsuL1Plugin_logic_shared_write_payload_data_dirty;
  wire                LsuL1Plugin_logic_shared_lsuRead_cmd_valid;
  wire       [5:0]    LsuL1Plugin_logic_shared_lsuRead_cmd_payload;
  (* keep , syn_keep *) wire       [0:0]    LsuL1Plugin_logic_shared_lsuRead_rsp_plru_0 /* synthesis syn_keep = 1 */ ;
  (* keep , syn_keep *) wire       [1:0]    LsuL1Plugin_logic_shared_lsuRead_rsp_dirty /* synthesis syn_keep = 1 */ ;
  wire       [2:0]    _zz_LsuL1Plugin_logic_shared_lsuRead_rsp_plru_0;
  reg                 LsuL1Plugin_logic_refill_slots_0_valid;
  reg                 LsuL1Plugin_logic_refill_slots_0_dirty;
  reg        [31:0]   LsuL1Plugin_logic_refill_slots_0_address;
  reg        [0:0]    LsuL1Plugin_logic_refill_slots_0_way;
  reg                 LsuL1Plugin_logic_refill_slots_0_cmdSent;
  reg                 LsuL1Plugin_logic_refill_slots_0_loadedSet;
  reg                 LsuL1Plugin_logic_refill_slots_0_loaded;
  reg        [0:0]    LsuL1Plugin_logic_refill_slots_0_loadedCounter;
  wire                LsuL1Plugin_logic_refill_slots_0_loadedDone;
  wire                LsuL1Plugin_logic_refill_slots_0_fire;
  wire                LsuL1Plugin_logic_refill_slots_0_free;
  reg        [0:0]    LsuL1Plugin_logic_refill_slots_0_victim;
  reg        [0:0]    LsuL1Plugin_logic_refill_slots_0_writebackHazards;
  wire       [0:0]    LsuL1Plugin_logic_refill_free;
  wire                LsuL1Plugin_logic_refill_full;
  reg                 LsuL1Plugin_logic_refill_push_valid;
  wire       [31:0]   LsuL1Plugin_logic_refill_push_payload_address;
  reg        [0:0]    LsuL1Plugin_logic_refill_push_payload_way;
  reg        [0:0]    LsuL1Plugin_logic_refill_push_payload_victim;
  wire                LsuL1Plugin_logic_refill_push_payload_dirty;
  wire                LsuL1Plugin_logic_refill_push_payload_unique;
  wire                LsuL1Plugin_logic_refill_push_payload_data;
  reg        [31:0]   LsuL1Plugin_logic_refill_pushCounter;
  wire                when_LsuL1Plugin_l358;
  wire                LsuL1Plugin_logic_refill_read_arbiter_slotsWithId_0_0;
  wire       [0:0]    LsuL1Plugin_logic_refill_read_arbiter_hits;
  wire                LsuL1Plugin_logic_refill_read_arbiter_hit;
  reg        [0:0]    LsuL1Plugin_logic_refill_read_arbiter_oh;
  reg        [0:0]    LsuL1Plugin_logic_refill_read_arbiter_lock;
  wire                when_LsuL1Plugin_l288;
  wire                LsuL1Plugin_logic_bus_read_cmd_fire;
  wire       [31:0]   LsuL1Plugin_logic_refill_read_cmdAddress;
  wire       [31:0]   LsuL1Plugin_logic_refill_read_rspAddress;
  wire                LsuL1Plugin_logic_refill_read_dirty;
  wire       [0:0]    LsuL1Plugin_logic_refill_read_way;
  (* keep , syn_keep *) reg        [2:0]    LsuL1Plugin_logic_refill_read_wordIndex /* synthesis syn_keep = 1 */ ;
  wire                LsuL1Plugin_logic_refill_read_rspWithData;
  reg        [1:0]    LsuL1Plugin_logic_refill_read_bankWriteNotif;
  wire                LsuL1Plugin_logic_refill_read_writeReservation_win;
  reg                 LsuL1Plugin_logic_refill_read_writeReservation_take;
  reg                 LsuL1Plugin_logic_refill_read_hadError;
  wire                when_LsuL1Plugin_l434;
  reg                 LsuL1Plugin_logic_refill_read_fire;
  wire                LsuL1Plugin_logic_refill_read_reservation_win;
  reg                 LsuL1Plugin_logic_refill_read_reservation_take;
  wire                LsuL1Plugin_logic_refill_read_faulty;
  wire                when_LsuL1Plugin_l446;
  wire       [0:0]    LsuL1_REFILL_BUSY;
  reg                 LsuL1Plugin_logic_writeback_slots_0_fire;
  reg                 LsuL1Plugin_logic_writeback_slots_0_valid;
  reg                 LsuL1Plugin_logic_writeback_slots_0_busy;
  reg        [31:0]   LsuL1Plugin_logic_writeback_slots_0_address;
  reg        [0:0]    LsuL1Plugin_logic_writeback_slots_0_way;
  reg                 LsuL1Plugin_logic_writeback_slots_0_readCmdDone;
  reg                 LsuL1Plugin_logic_writeback_slots_0_victimBufferReady;
  reg                 LsuL1Plugin_logic_writeback_slots_0_readRspDone;
  reg                 LsuL1Plugin_logic_writeback_slots_0_writeCmdDone;
  reg        [0:0]    LsuL1Plugin_logic_writeback_slots_0_timer_counter;
  wire                LsuL1Plugin_logic_writeback_slots_0_timer_done;
  wire                when_LsuL1Plugin_l509;
  wire                LsuL1Plugin_logic_writeback_slots_0_free;
  wire       [0:0]    LsuL1_WRITEBACK_BUSY;
  wire       [0:0]    LsuL1Plugin_logic_writeback_free;
  wire                LsuL1Plugin_logic_writeback_full;
  reg                 LsuL1Plugin_logic_writeback_push_valid;
  reg        [31:0]   LsuL1Plugin_logic_writeback_push_payload_address;
  reg        [0:0]    LsuL1Plugin_logic_writeback_push_payload_way;
  wire                when_LsuL1Plugin_l532;
  wire                LsuL1Plugin_logic_writeback_read_arbiter_slotsWithId_0_0;
  wire       [0:0]    LsuL1Plugin_logic_writeback_read_arbiter_hits;
  wire                LsuL1Plugin_logic_writeback_read_arbiter_hit;
  reg        [0:0]    LsuL1Plugin_logic_writeback_read_arbiter_oh;
  reg        [0:0]    LsuL1Plugin_logic_writeback_read_arbiter_lock;
  wire                when_LsuL1Plugin_l288_1;
  wire       [31:0]   LsuL1Plugin_logic_writeback_read_address;
  wire       [0:0]    LsuL1Plugin_logic_writeback_read_way;
  (* keep , syn_keep *) reg        [2:0]    LsuL1Plugin_logic_writeback_read_wordIndex /* synthesis syn_keep = 1 */ ;
  wire                LsuL1Plugin_logic_writeback_read_slotRead_valid;
  wire                LsuL1Plugin_logic_writeback_read_slotRead_payload_last;
  wire       [2:0]    LsuL1Plugin_logic_writeback_read_slotRead_payload_wordIndex;
  wire       [0:0]    LsuL1Plugin_logic_writeback_read_slotRead_payload_way;
  wire                when_LsuL1Plugin_l577;
  reg                 LsuL1Plugin_logic_writeback_read_slotReadLast_valid;
  reg                 LsuL1Plugin_logic_writeback_read_slotReadLast_payload_last;
  reg        [2:0]    LsuL1Plugin_logic_writeback_read_slotReadLast_payload_wordIndex;
  reg        [0:0]    LsuL1Plugin_logic_writeback_read_slotReadLast_payload_way;
  wire       [63:0]   LsuL1Plugin_logic_writeback_read_readedData;
  wire                LsuL1Plugin_logic_writeback_write_arbiter_slotsWithId_0_0;
  wire       [0:0]    LsuL1Plugin_logic_writeback_write_arbiter_hits;
  wire                LsuL1Plugin_logic_writeback_write_arbiter_hit;
  reg        [0:0]    LsuL1Plugin_logic_writeback_write_arbiter_oh;
  reg        [0:0]    LsuL1Plugin_logic_writeback_write_arbiter_lock;
  wire                when_LsuL1Plugin_l288_2;
  (* keep , syn_keep *) reg        [2:0]    LsuL1Plugin_logic_writeback_write_wordIndex /* synthesis syn_keep = 1 */ ;
  wire                LsuL1Plugin_logic_writeback_write_last;
  wire                LsuL1Plugin_logic_writeback_write_bufferRead_valid;
  reg                 LsuL1Plugin_logic_writeback_write_bufferRead_ready;
  wire       [31:0]   LsuL1Plugin_logic_writeback_write_bufferRead_payload_address;
  wire                LsuL1Plugin_logic_writeback_write_bufferRead_payload_last;
  wire                LsuL1Plugin_logic_writeback_write_bufferRead_fire;
  wire                when_LsuL1Plugin_l651;
  wire                LsuL1Plugin_logic_writeback_write_cmd_valid;
  wire                LsuL1Plugin_logic_writeback_write_cmd_ready;
  wire       [31:0]   LsuL1Plugin_logic_writeback_write_cmd_payload_address;
  wire                LsuL1Plugin_logic_writeback_write_cmd_payload_last;
  reg                 LsuL1Plugin_logic_writeback_write_bufferRead_rValid;
  reg        [31:0]   LsuL1Plugin_logic_writeback_write_bufferRead_rData_address;
  reg                 LsuL1Plugin_logic_writeback_write_bufferRead_rData_last;
  wire                when_Stream_l393_2;
  wire       [2:0]    _zz_LsuL1Plugin_logic_writeback_write_word;
  wire       [63:0]   LsuL1Plugin_logic_writeback_write_word;
  wire       [8:0]    LsuL1Plugin_logic_ls_rb0_readAddress;
  wire                when_LsuL1Plugin_l690;
  wire                when_LsuL1Plugin_l691;
  wire                when_LsuL1Plugin_l690_1;
  wire                when_LsuL1Plugin_l691_1;
  reg                 LsuL1Plugin_logic_ls_rb1_onBanks_0_busyReg;
  wire                when_LsuL1Plugin_l706;
  reg                 LsuL1Plugin_logic_ls_rb1_onBanks_1_busyReg;
  wire                when_LsuL1Plugin_l706_1;
  wire                _zz_toplevel_execute_ctrl4_down_LsuL1Plugin_logic_MUXED_DATA_lane0;
  wire                _zz_toplevel_execute_ctrl4_down_LsuL1Plugin_logic_MUXED_DATA_lane0_1;
  wire                LsuL1Plugin_logic_ls_sharedBypassers_0_hit;
  wire       [0:0]    LsuL1Plugin_logic_ls_ctrl_plruLogic_core_io_context_state_0;
  wire       [0:0]    LsuL1Plugin_logic_ls_ctrl_plruLogic_core_io_evict_id;
  reg        [0:0]    LsuL1Plugin_logic_ls_ctrl_plruLogic_core_io_update_id;
  wire       [0:0]    LsuL1Plugin_logic_ls_ctrl_plruLogic_core_io_update_state_0;
  wire                LsuL1Plugin_logic_ls_ctrl_plruLogic_core_evict_sel_0;
  wire                LsuL1Plugin_logic_ls_ctrl_plruLogic_core_evict_logic_0_state;
  wire                LsuL1Plugin_logic_ls_ctrl_wayWriteReservation_win;
  reg                 LsuL1Plugin_logic_ls_ctrl_wayWriteReservation_take;
  wire                LsuL1Plugin_logic_ls_ctrl_bankWriteReservation_win;
  wire                LsuL1Plugin_logic_ls_ctrl_bankWriteReservation_take;
  wire       [0:0]    LsuL1Plugin_logic_ls_ctrl_refillWayWithoutUpdate;
  wire                LsuL1Plugin_logic_ls_ctrl_refillWayNeedWriteback;
  wire       [0:0]    LsuL1Plugin_logic_ls_ctrl_refillHazards;
  wire       [0:0]    LsuL1Plugin_logic_ls_ctrl_writebackHazards;
  wire                LsuL1Plugin_logic_ls_ctrl_refillHazard;
  wire                LsuL1Plugin_logic_ls_ctrl_writebackHazard;
  wire                LsuL1Plugin_logic_ls_ctrl_wasDirty;
  wire       [1:0]    LsuL1Plugin_logic_ls_ctrl_loadedDirties;
  wire                LsuL1Plugin_logic_ls_ctrl_refillWayWasDirty;
  wire                LsuL1Plugin_logic_ls_ctrl_writeToReadHazard;
  wire                LsuL1Plugin_logic_ls_ctrl_bankNotRead;
  wire                LsuL1Plugin_logic_ls_ctrl_loadHazard;
  wire                LsuL1Plugin_logic_ls_ctrl_storeHazard;
  wire                LsuL1Plugin_logic_ls_ctrl_flushHazard;
  wire                LsuL1Plugin_logic_ls_ctrl_coherencyHazard;
  reg                 LsuL1Plugin_logic_ls_ctrl_hazardReg;
  reg                 LsuL1Plugin_logic_ls_ctrl_flushHazardReg;
  wire                LsuL1Plugin_logic_ls_ctrl_canRefill;
  wire                LsuL1Plugin_logic_ls_ctrl_canFlush;
  wire       [1:0]    LsuL1Plugin_logic_ls_ctrl_needFlushs;
  wire       [1:0]    _zz_LsuL1Plugin_logic_ls_ctrl_needFlushs_bools_0;
  wire                LsuL1Plugin_logic_ls_ctrl_needFlushs_bools_0;
  wire                LsuL1Plugin_logic_ls_ctrl_needFlushs_bools_1;
  reg        [1:0]    _zz_LsuL1Plugin_logic_ls_ctrl_needFlushOh;
  wire       [1:0]    LsuL1Plugin_logic_ls_ctrl_needFlushOh;
  wire                _zz_LsuL1Plugin_logic_ls_ctrl_needFlushSel;
  wire       [0:0]    LsuL1Plugin_logic_ls_ctrl_needFlushSel;
  wire                LsuL1Plugin_logic_ls_ctrl_isAccess;
  wire                LsuL1Plugin_logic_ls_ctrl_askRefill;
  wire                LsuL1Plugin_logic_ls_ctrl_askUpgrade;
  wire                LsuL1Plugin_logic_ls_ctrl_askFlush;
  wire                LsuL1Plugin_logic_ls_ctrl_doRefill;
  wire                LsuL1Plugin_logic_ls_ctrl_doUpgrade;
  wire                LsuL1Plugin_logic_ls_ctrl_doFlush;
  wire                LsuL1Plugin_logic_ls_ctrl_doWrite;
  wire       [0:0]    LsuL1Plugin_logic_ls_ctrl_wayId;
  wire       [0:0]    LsuL1Plugin_logic_ls_ctrl_targetWay;
  wire                LsuL1Plugin_logic_ls_ctrl_doRefillPush;
  wire                when_LsuL1Plugin_l876;
  wire       [2:0]    _zz_38;
  wire       [1:0]    _zz_39;
  wire                when_LsuL1Plugin_l890;
  wire                when_LsuL1Plugin_l890_1;
  wire       [19:0]   _zz_LsuL1Plugin_logic_waysWrite_tag_address;
  wire                when_LsuL1Plugin_l956;
  wire                when_LsuL1Plugin_l963;
  wire                when_LsuL1Plugin_l967;
  wire                when_LsuL1Plugin_l967_1;
  wire                when_LsuL1Plugin_l967_2;
  wire                when_LsuL1Plugin_l967_3;
  wire                when_LsuL1Plugin_l963_1;
  wire                when_LsuL1Plugin_l967_4;
  wire                when_LsuL1Plugin_l967_5;
  wire                when_LsuL1Plugin_l967_6;
  wire                when_LsuL1Plugin_l967_7;
  wire                LsuL1Plugin_logic_ls_ctrl_preventSideEffects;
  reg        [6:0]    LsuL1Plugin_logic_initializer_counter;
  wire                LsuL1Plugin_logic_initializer_done;
  wire                when_LsuL1Plugin_l1160;
  wire       [2:0]    _zz_LsuL1Plugin_logic_shared_write_payload_data_plru_0;
  reg        [9:0]    LsuL1Plugin_logic_initializerMem_counter;
  wire                LsuL1Plugin_logic_initializerMem_busy;
  reg                 TrapPlugin_logic_harts_0_crsPorts_write_valid;
  wire                TrapPlugin_logic_harts_0_crsPorts_write_ready;
  reg        [2:0]    TrapPlugin_logic_harts_0_crsPorts_write_address;
  reg        [31:0]   TrapPlugin_logic_harts_0_crsPorts_write_data;
  reg        [0:0]    LsuPlugin_logic_flusher_waiter;
  wire       [4:0]    LsuPlugin_logic_onAddress0_ls_prefetchOp;
  wire                LsuPlugin_logic_onAddress0_ls_port_valid;
  wire                LsuPlugin_logic_onAddress0_ls_port_ready;
  wire       [2:0]    LsuPlugin_logic_onAddress0_ls_port_payload_op;
  wire       [31:0]   LsuPlugin_logic_onAddress0_ls_port_payload_address;
  wire       [1:0]    LsuPlugin_logic_onAddress0_ls_port_payload_size;
  wire                LsuPlugin_logic_onAddress0_ls_port_payload_load;
  wire                LsuPlugin_logic_onAddress0_ls_port_payload_store;
  wire                LsuPlugin_logic_onAddress0_ls_port_payload_atomic;
  wire       [11:0]   LsuPlugin_logic_onAddress0_ls_port_payload_storeId;
  reg        [11:0]   LsuPlugin_logic_onAddress0_ls_storeId;
  wire                LsuPlugin_logic_onAddress0_ls_port_fire;
  reg        [0:0]    LsuPlugin_logic_onAddress0_access_waiter_refill;
  reg                 LsuPlugin_logic_onAddress0_access_waiter_valid;
  wire                when_LsuPlugin_l200;
  wire                LsuPlugin_logic_onAddress0_access_sbWaiter;
  wire                LsuPlugin_logic_onAddress0_access_port_valid;
  wire                LsuPlugin_logic_onAddress0_access_port_ready;
  wire       [2:0]    LsuPlugin_logic_onAddress0_access_port_payload_op;
  wire       [31:0]   LsuPlugin_logic_onAddress0_access_port_payload_address;
  wire       [1:0]    LsuPlugin_logic_onAddress0_access_port_payload_size;
  wire                LsuPlugin_logic_onAddress0_access_port_payload_load;
  wire                LsuPlugin_logic_onAddress0_access_port_payload_store;
  wire                LsuPlugin_logic_onAddress0_access_port_payload_atomic;
  wire       [11:0]   LsuPlugin_logic_onAddress0_access_port_payload_storeId;
  wire                _zz_MmuPlugin_logic_accessBus_cmd_ready;
  wire                LsuPlugin_logic_onAddress0_flush_port_valid;
  wire                LsuPlugin_logic_onAddress0_flush_port_ready;
  wire       [2:0]    LsuPlugin_logic_onAddress0_flush_port_payload_op;
  wire       [31:0]   LsuPlugin_logic_onAddress0_flush_port_payload_address;
  wire       [1:0]    LsuPlugin_logic_onAddress0_flush_port_payload_size;
  wire                LsuPlugin_logic_onAddress0_flush_port_payload_load;
  wire                LsuPlugin_logic_onAddress0_flush_port_payload_store;
  wire                LsuPlugin_logic_onAddress0_flush_port_payload_atomic;
  wire       [11:0]   LsuPlugin_logic_onAddress0_flush_port_payload_storeId;
  wire                LsuPlugin_logic_onAddress0_flush_port_fire;
  reg        [3:0]    _zz_toplevel_execute_ctrl2_down_LsuL1_MASK_lane0;
  wire                when_LsuPlugin_l449;
  wire                when_LsuPlugin_l449_1;
  wire       [31:0]   LsuPlugin_logic_onPma_cached_cmd_address;
  wire       [0:0]    LsuPlugin_logic_onPma_cached_cmd_op;
  wire                LsuPlugin_logic_onPma_cached_rsp_fault;
  wire                LsuPlugin_logic_onPma_cached_rsp_io;
  wire       [31:0]   LsuPlugin_logic_onPma_io_cmd_address;
  wire       [1:0]    LsuPlugin_logic_onPma_io_cmd_size;
  wire       [0:0]    LsuPlugin_logic_onPma_io_cmd_op;
  wire                LsuPlugin_logic_onPma_io_rsp_fault;
  wire                LsuPlugin_logic_onPma_io_rsp_io;
  wire                LsuPlugin_logic_onPma_addressExtension;
  reg                 LsuPlugin_logic_onCtrl_lsuTrap;
  reg        [31:0]   LsuPlugin_logic_onCtrl_writeData;
  wire                LsuPlugin_logic_onCtrl_scMiss;
  reg                 LsuPlugin_logic_onCtrl_io_tooEarly;
  reg                 LsuPlugin_logic_onCtrl_io_allowIt;
  wire                when_LsuPlugin_l491;
  wire                LsuPlugin_logic_onCtrl_io_doIt;
  reg                 LsuPlugin_logic_onCtrl_io_doItReg;
  reg                 LsuPlugin_logic_onCtrl_io_cmdSent;
  wire                LsuPlugin_logic_bus_cmd_fire;
  wire                when_LsuPlugin_l495;
  wire                LsuPlugin_logic_bus_rsp_toStream_valid;
  wire                LsuPlugin_logic_bus_rsp_toStream_ready;
  wire                LsuPlugin_logic_bus_rsp_toStream_payload_error;
  wire       [31:0]   LsuPlugin_logic_bus_rsp_toStream_payload_data;
  wire                LsuPlugin_logic_onCtrl_io_rsp_valid;
  wire                LsuPlugin_logic_onCtrl_io_rsp_ready;
  wire                LsuPlugin_logic_onCtrl_io_rsp_payload_error;
  wire       [31:0]   LsuPlugin_logic_onCtrl_io_rsp_payload_data;
  reg                 LsuPlugin_logic_bus_rsp_toStream_rValid;
  wire                LsuPlugin_logic_onCtrl_io_rsp_fire;
  reg                 LsuPlugin_logic_bus_rsp_toStream_rData_error;
  reg        [31:0]   LsuPlugin_logic_bus_rsp_toStream_rData_data;
  wire                LsuPlugin_logic_onCtrl_io_freezeIt;
  wire       [31:0]   LsuPlugin_logic_onCtrl_loadData_input;
  wire       [7:0]    LsuPlugin_logic_onCtrl_loadData_splited_0;
  wire       [7:0]    LsuPlugin_logic_onCtrl_loadData_splited_1;
  wire       [7:0]    LsuPlugin_logic_onCtrl_loadData_splited_2;
  wire       [7:0]    LsuPlugin_logic_onCtrl_loadData_splited_3;
  reg        [31:0]   LsuPlugin_logic_onCtrl_loadData_shited;
  wire       [31:0]   LsuPlugin_logic_onCtrl_storeData_mapping_0_1;
  wire       [31:0]   LsuPlugin_logic_onCtrl_storeData_mapping_1_1;
  wire       [31:0]   LsuPlugin_logic_onCtrl_storeData_mapping_2_1;
  reg        [31:0]   _zz_toplevel_execute_ctrl4_down_LsuL1_WRITE_DATA_lane0;
  reg        [31:0]   LsuPlugin_logic_onCtrl_rva_srcBuffer;
  wire       [2:0]    _zz_LsuPlugin_logic_onCtrl_rva_alu_compare;
  wire                _zz_LsuPlugin_logic_onCtrl_rva_alu_selectRf;
  wire                LsuPlugin_logic_onCtrl_rva_alu_compare;
  wire                LsuPlugin_logic_onCtrl_rva_alu_unsigned;
  wire       [31:0]   LsuPlugin_logic_onCtrl_rva_alu_addSub;
  wire                LsuPlugin_logic_onCtrl_rva_alu_less;
  wire                LsuPlugin_logic_onCtrl_rva_alu_selectRf;
  wire       [2:0]    switch_Misc_l241_4;
  reg        [31:0]   LsuPlugin_logic_onCtrl_rva_alu_raw;
  wire       [31:0]   LsuPlugin_logic_onCtrl_rva_alu_result;
  reg        [31:0]   LsuPlugin_logic_onCtrl_rva_aluBuffer;
  wire                LsuPlugin_logic_onCtrl_rva_delay_0;
  wire                LsuPlugin_logic_onCtrl_rva_delay_1;
  reg                 _zz_LsuPlugin_logic_onCtrl_rva_delay_0;
  reg                 _zz_LsuPlugin_logic_onCtrl_rva_delay_1;
  wire                LsuPlugin_logic_onCtrl_rva_freezeIt;
  reg                 LsuPlugin_logic_onCtrl_rva_nc_capture;
  reg                 LsuPlugin_logic_onCtrl_rva_nc_reserved;
  reg        [31:0]   LsuPlugin_logic_onCtrl_rva_nc_address;
  wire                when_LsuPlugin_l573;
  reg        [5:0]    LsuPlugin_logic_onCtrl_rva_nc_age;
  wire                when_LsuPlugin_l585;
  wire                LsuPlugin_logic_onCtrl_traps_accessFault;
  wire                LsuPlugin_logic_onCtrl_traps_l1Failed;
  wire                LsuPlugin_logic_onCtrl_traps_pmaFault;
  wire                when_LsuPlugin_l683;
  wire                when_LsuPlugin_l710;
  wire                when_LsuPlugin_l723;
  wire                LsuPlugin_logic_onCtrl_mmuNeeded;
  wire                when_LsuPlugin_l761;
  wire                when_LsuPlugin_l796;
  wire                when_LsuPlugin_l204;
  reg        [0:0]    LsuPlugin_logic_onCtrl_hartRegulation_refill;
  reg                 LsuPlugin_logic_onCtrl_hartRegulation_valid;
  wire                when_LsuPlugin_l200_1;
  wire                when_LsuPlugin_l803;
  wire                when_LsuPlugin_l204_1;
  wire                when_LsuPlugin_l824;
  wire                LsuPlugin_logic_onWb_storeFire;
  wire                LsuPlugin_logic_onWb_storeBroadcast;
  reg                 LsuL1Plugin_logic_bus_toTilelink_nonCoherent_onA_lock;
  wire                LsuL1TileLinkPlugin_logic_down_a_fire;
  reg        [2:0]    LsuL1Plugin_logic_bus_toTilelink_nonCoherent_onA_beat;
  wire                LsuL1TileLinkPlugin_logic_down_a_tracker_last;
  wire                when_LsuL1Bus_l402;
  reg                 LsuL1Plugin_logic_bus_toTilelink_nonCoherent_onA_selReg;
  wire                LsuL1Plugin_logic_bus_toTilelink_nonCoherent_onA_sel;
  wire                LsuL1Plugin_logic_bus_toTilelink_nonCoherent_onD_sel;
  reg                 TrapPlugin_logic_harts_0_interrupt_valid;
  reg        [3:0]    TrapPlugin_logic_harts_0_interrupt_code;
  reg        [1:0]    TrapPlugin_logic_harts_0_interrupt_targetPrivilege;
  wire                when_TrapPlugin_l189;
  wire                when_TrapPlugin_l189_1;
  wire                when_TrapPlugin_l195;
  wire                when_TrapPlugin_l195_1;
  wire                when_TrapPlugin_l195_2;
  wire                when_TrapPlugin_l195_3;
  wire                when_TrapPlugin_l195_4;
  wire                when_TrapPlugin_l195_5;
  wire                when_TrapPlugin_l195_6;
  wire                when_TrapPlugin_l195_7;
  wire                when_TrapPlugin_l195_8;
  reg                 TrapPlugin_logic_harts_0_interrupt_validBuffer;
  wire                TrapPlugin_logic_harts_0_interrupt_pendingInterrupt;
  wire                when_TrapPlugin_l214;
  wire                _zz_TrapPlugin_logic_harts_0_trap_pending_arbiter_ports_1_valid;
  wire                _zz_TrapPlugin_logic_harts_0_trap_pending_arbiter_ports_3_valid;
  wire                _zz_TrapPlugin_logic_harts_0_trap_pending_arbiter_ports_0_valid;
  wire                _zz_TrapPlugin_logic_harts_0_trap_pending_arbiter_ports_1_valid_1;
  wire                _zz_TrapPlugin_logic_harts_0_trap_pending_arbiter_ports_2_valid;
  wire                _zz_TrapPlugin_logic_harts_0_trap_pending_arbiter_ports_2_valid_1;
  wire                TrapPlugin_logic_harts_0_trap_pending_arbiter_ports_0_valid;
  wire                TrapPlugin_logic_harts_0_trap_pending_arbiter_ports_0_payload_exception;
  wire       [31:0]   TrapPlugin_logic_harts_0_trap_pending_arbiter_ports_0_payload_tval;
  wire       [3:0]    TrapPlugin_logic_harts_0_trap_pending_arbiter_ports_0_payload_code;
  wire       [2:0]    TrapPlugin_logic_harts_0_trap_pending_arbiter_ports_0_payload_arg;
  wire                TrapPlugin_logic_harts_0_trap_pending_arbiter_ports_1_valid;
  wire                TrapPlugin_logic_harts_0_trap_pending_arbiter_ports_1_payload_exception;
  wire       [31:0]   TrapPlugin_logic_harts_0_trap_pending_arbiter_ports_1_payload_tval;
  wire       [3:0]    TrapPlugin_logic_harts_0_trap_pending_arbiter_ports_1_payload_code;
  wire       [2:0]    TrapPlugin_logic_harts_0_trap_pending_arbiter_ports_1_payload_arg;
  wire       [1:0]    _zz_TrapPlugin_logic_harts_0_trap_pending_arbiter_ports_1_payload_exception;
  wire       [39:0]   _zz_TrapPlugin_logic_harts_0_trap_pending_arbiter_ports_1_payload_exception_1;
  wire                TrapPlugin_logic_harts_0_trap_pending_arbiter_ports_2_valid;
  wire                TrapPlugin_logic_harts_0_trap_pending_arbiter_ports_2_payload_exception;
  wire       [31:0]   TrapPlugin_logic_harts_0_trap_pending_arbiter_ports_2_payload_tval;
  wire       [3:0]    TrapPlugin_logic_harts_0_trap_pending_arbiter_ports_2_payload_code;
  wire       [2:0]    TrapPlugin_logic_harts_0_trap_pending_arbiter_ports_2_payload_arg;
  wire       [1:0]    _zz_TrapPlugin_logic_harts_0_trap_pending_arbiter_ports_2_payload_exception;
  wire       [39:0]   _zz_TrapPlugin_logic_harts_0_trap_pending_arbiter_ports_2_payload_exception_1;
  wire                TrapPlugin_logic_harts_0_trap_pending_arbiter_ports_3_valid;
  wire                TrapPlugin_logic_harts_0_trap_pending_arbiter_ports_3_payload_exception;
  wire       [31:0]   TrapPlugin_logic_harts_0_trap_pending_arbiter_ports_3_payload_tval;
  wire       [3:0]    TrapPlugin_logic_harts_0_trap_pending_arbiter_ports_3_payload_code;
  wire       [2:0]    TrapPlugin_logic_harts_0_trap_pending_arbiter_ports_3_payload_arg;
  wire       [3:0]    _zz_TrapPlugin_logic_harts_0_trap_pending_arbiter_oh;
  wire                _zz_TrapPlugin_logic_harts_0_trap_pending_arbiter_oh_1;
  wire                _zz_TrapPlugin_logic_harts_0_trap_pending_arbiter_oh_2;
  wire                _zz_TrapPlugin_logic_harts_0_trap_pending_arbiter_oh_3;
  reg        [3:0]    _zz_TrapPlugin_logic_harts_0_trap_pending_arbiter_oh_4;
  wire       [3:0]    TrapPlugin_logic_harts_0_trap_pending_arbiter_oh;
  wire                TrapPlugin_logic_harts_0_trap_pending_arbiter_down_valid;
  wire                TrapPlugin_logic_harts_0_trap_pending_arbiter_down_payload_exception;
  wire       [31:0]   TrapPlugin_logic_harts_0_trap_pending_arbiter_down_payload_tval;
  wire       [3:0]    TrapPlugin_logic_harts_0_trap_pending_arbiter_down_payload_code;
  wire       [2:0]    TrapPlugin_logic_harts_0_trap_pending_arbiter_down_payload_arg;
  wire       [39:0]   _zz_TrapPlugin_logic_harts_0_trap_pending_arbiter_down_payload_exception;
  reg                 TrapPlugin_logic_harts_0_trap_pending_state_exception;
  reg        [31:0]   TrapPlugin_logic_harts_0_trap_pending_state_tval;
  reg        [3:0]    TrapPlugin_logic_harts_0_trap_pending_state_code;
  reg        [2:0]    TrapPlugin_logic_harts_0_trap_pending_state_arg;
  reg        [31:0]   TrapPlugin_logic_harts_0_trap_pending_pc;
  reg        [11:0]   TrapPlugin_logic_harts_0_trap_pending_history;
  reg        [1:0]    TrapPlugin_logic_harts_0_trap_pending_slices;
  wire       [1:0]    TrapPlugin_logic_harts_0_trap_pending_xret_sourcePrivilege;
  reg        [1:0]    TrapPlugin_logic_harts_0_trap_pending_xret_targetPrivilege;
  reg        [1:0]    TrapPlugin_logic_harts_0_trap_exception_exceptionTargetPrivilegeUncapped;
  wire       [3:0]    TrapPlugin_logic_harts_0_trap_exception_code;
  wire                when_TrapPlugin_l251;
  wire                when_TrapPlugin_l251_1;
  wire                when_TrapPlugin_l251_2;
  wire                when_TrapPlugin_l251_3;
  wire                when_TrapPlugin_l251_4;
  wire                when_TrapPlugin_l251_5;
  wire                when_TrapPlugin_l251_6;
  wire       [1:0]    TrapPlugin_logic_harts_0_trap_exception_targetPrivilege;
  wire                toplevel_execute_lane0_ctrls_5_upIsCancel;
  wire                toplevel_execute_lane0_ctrls_5_downIsCancel;
  wire                toplevel_execute_lane1_ctrls_5_upIsCancel;
  wire                toplevel_execute_lane1_ctrls_5_downIsCancel;
  wire       [1:0]    TrapPlugin_logic_harts_0_trap_trigger_oh;
  wire                TrapPlugin_logic_harts_0_trap_trigger_valid;
  wire                _zz_TrapPlugin_logic_harts_0_trap_pending_pc;
  wire                _zz_TrapPlugin_logic_harts_0_trap_pending_pc_1;
  reg                 TrapPlugin_logic_harts_0_trap_whitebox_trap;
  reg                 TrapPlugin_logic_harts_0_trap_whitebox_interrupt;
  reg        [3:0]    TrapPlugin_logic_harts_0_trap_whitebox_code;
  reg                 TrapPlugin_logic_harts_0_trap_historyPort_valid;
  wire       [11:0]   TrapPlugin_logic_harts_0_trap_historyPort_payload_history;
  reg                 TrapPlugin_logic_harts_0_trap_pcPort_valid;
  wire                TrapPlugin_logic_harts_0_trap_pcPort_payload_fault;
  reg        [31:0]   TrapPlugin_logic_harts_0_trap_pcPort_payload_pc;
  wire                PcPlugin_logic_harts_0_aggregator_sortedByPriority_0_laneValid;
  wire                TrapPlugin_logic_harts_0_trap_fsm_wantExit;
  reg                 TrapPlugin_logic_harts_0_trap_fsm_wantStart;
  wire                TrapPlugin_logic_harts_0_trap_fsm_wantKill;
  wire                TrapPlugin_logic_harts_0_trap_fsm_inflightTrap;
  wire                TrapPlugin_logic_harts_0_trap_fsm_holdPort;
  reg                 TrapPlugin_logic_harts_0_trap_fsm_wfi;
  reg                 TrapPlugin_logic_harts_0_trap_fsm_buffer_sampleIt;
  reg                 TrapPlugin_logic_harts_0_trap_fsm_buffer_i_valid;
  reg        [3:0]    TrapPlugin_logic_harts_0_trap_fsm_buffer_i_code;
  reg        [1:0]    TrapPlugin_logic_harts_0_trap_fsm_buffer_i_targetPrivilege;
  wire                TrapPlugin_logic_harts_0_trap_fsm_buffer_trap_interrupt;
  wire       [1:0]    TrapPlugin_logic_harts_0_trap_fsm_buffer_trap_targetPrivilege;
  wire       [31:0]   TrapPlugin_logic_harts_0_trap_fsm_buffer_trap_tval;
  wire       [3:0]    TrapPlugin_logic_harts_0_trap_fsm_buffer_trap_code;
  wire                TrapPlugin_logic_harts_0_trap_fsm_resetToRunConditions_0;
  reg                 TrapPlugin_logic_harts_0_trap_fsm_atsPorts_refill_cmd_valid;
  wire                TrapPlugin_logic_harts_0_trap_fsm_atsPorts_refill_cmd_ready;
  wire       [31:0]   TrapPlugin_logic_harts_0_trap_fsm_atsPorts_refill_cmd_payload_address;
  wire       [0:0]    TrapPlugin_logic_harts_0_trap_fsm_atsPorts_refill_cmd_payload_storageId;
  reg                 TrapPlugin_logic_harts_0_trap_fsm_atsPorts_refill_rsp_valid;
  reg                 TrapPlugin_logic_harts_0_trap_fsm_atsPorts_refill_rsp_payload_pageFault;
  reg                 TrapPlugin_logic_harts_0_trap_fsm_atsPorts_refill_rsp_payload_accessFault;
  reg                 TrapPlugin_logic_harts_0_trap_fsm_atsPorts_invalidate_cmd_valid;
  wire                TrapPlugin_logic_harts_0_trap_fsm_atsPorts_invalidate_cmd_ready;
  reg                 TrapPlugin_logic_harts_0_trap_fsm_atsPorts_invalidated;
  wire                TrapPlugin_logic_harts_0_trap_fsm_atsPorts_invalidate_cmd_fire;
  wire                when_TrapPlugin_l340;
  reg        [31:0]   TrapPlugin_logic_harts_0_trap_fsm_jumpTarget;
  wire       [1:0]    TrapPlugin_logic_harts_0_trap_fsm_jumpOffset;
  reg                 TrapPlugin_logic_harts_0_trap_fsm_trapEnterDebug;
  wire                TrapPlugin_logic_harts_0_trap_fsm_triggerEbreak;
  reg                 TrapPlugin_logic_harts_0_trap_fsm_triggerEbreakReg;
  wire                when_TrapPlugin_l539;
  reg        [31:0]   TrapPlugin_logic_harts_0_trap_fsm_readed;
  wire       [1:0]    TrapPlugin_logic_harts_0_trap_fsm_xretPrivilege;
  reg        [1:0]    FetchL1Plugin_logic_translationStorage_logic_sl_0_write_mask;
  reg        [5:0]    FetchL1Plugin_logic_translationStorage_logic_sl_0_write_address;
  reg                 FetchL1Plugin_logic_translationStorage_logic_sl_0_write_data_valid;
  reg        [13:0]   FetchL1Plugin_logic_translationStorage_logic_sl_0_write_data_virtualAddress;
  reg        [19:0]   FetchL1Plugin_logic_translationStorage_logic_sl_0_write_data_physicalAddress;
  reg                 FetchL1Plugin_logic_translationStorage_logic_sl_0_write_data_allowRead;
  reg                 FetchL1Plugin_logic_translationStorage_logic_sl_0_write_data_allowWrite;
  reg                 FetchL1Plugin_logic_translationStorage_logic_sl_0_write_data_allowExecute;
  reg                 FetchL1Plugin_logic_translationStorage_logic_sl_0_write_data_allowUser;
  reg                 FetchL1Plugin_logic_translationStorage_logic_sl_0_allocId_willIncrement;
  wire                FetchL1Plugin_logic_translationStorage_logic_sl_0_allocId_willClear;
  reg        [0:0]    FetchL1Plugin_logic_translationStorage_logic_sl_0_allocId_valueNext;
  reg        [0:0]    FetchL1Plugin_logic_translationStorage_logic_sl_0_allocId_value;
  wire                FetchL1Plugin_logic_translationStorage_logic_sl_0_allocId_willOverflowIfInc;
  wire                FetchL1Plugin_logic_translationStorage_logic_sl_0_allocId_willOverflow;
  reg        [0:0]    FetchL1Plugin_logic_translationStorage_logic_sl_1_write_mask;
  reg        [5:0]    FetchL1Plugin_logic_translationStorage_logic_sl_1_write_address;
  reg                 FetchL1Plugin_logic_translationStorage_logic_sl_1_write_data_valid;
  reg        [3:0]    FetchL1Plugin_logic_translationStorage_logic_sl_1_write_data_virtualAddress;
  reg        [9:0]    FetchL1Plugin_logic_translationStorage_logic_sl_1_write_data_physicalAddress;
  reg                 FetchL1Plugin_logic_translationStorage_logic_sl_1_write_data_allowRead;
  reg                 FetchL1Plugin_logic_translationStorage_logic_sl_1_write_data_allowWrite;
  reg                 FetchL1Plugin_logic_translationStorage_logic_sl_1_write_data_allowExecute;
  reg                 FetchL1Plugin_logic_translationStorage_logic_sl_1_write_data_allowUser;
  reg                 FetchL1Plugin_logic_translationStorage_logic_sl_1_allocId_willIncrement;
  wire                FetchL1Plugin_logic_translationStorage_logic_sl_1_allocId_willClear;
  wire                FetchL1Plugin_logic_translationStorage_logic_sl_1_allocId_willOverflowIfInc;
  wire                FetchL1Plugin_logic_translationStorage_logic_sl_1_allocId_willOverflow;
  reg        [1:0]    LsuPlugin_logic_translationStorage_logic_sl_0_write_mask;
  reg        [5:0]    LsuPlugin_logic_translationStorage_logic_sl_0_write_address;
  reg                 LsuPlugin_logic_translationStorage_logic_sl_0_write_data_valid;
  reg        [13:0]   LsuPlugin_logic_translationStorage_logic_sl_0_write_data_virtualAddress;
  reg        [19:0]   LsuPlugin_logic_translationStorage_logic_sl_0_write_data_physicalAddress;
  reg                 LsuPlugin_logic_translationStorage_logic_sl_0_write_data_allowRead;
  reg                 LsuPlugin_logic_translationStorage_logic_sl_0_write_data_allowWrite;
  reg                 LsuPlugin_logic_translationStorage_logic_sl_0_write_data_allowExecute;
  reg                 LsuPlugin_logic_translationStorage_logic_sl_0_write_data_allowUser;
  reg                 LsuPlugin_logic_translationStorage_logic_sl_0_allocId_willIncrement;
  wire                LsuPlugin_logic_translationStorage_logic_sl_0_allocId_willClear;
  reg        [0:0]    LsuPlugin_logic_translationStorage_logic_sl_0_allocId_valueNext;
  reg        [0:0]    LsuPlugin_logic_translationStorage_logic_sl_0_allocId_value;
  wire                LsuPlugin_logic_translationStorage_logic_sl_0_allocId_willOverflowIfInc;
  wire                LsuPlugin_logic_translationStorage_logic_sl_0_allocId_willOverflow;
  reg        [0:0]    LsuPlugin_logic_translationStorage_logic_sl_1_write_mask;
  reg        [5:0]    LsuPlugin_logic_translationStorage_logic_sl_1_write_address;
  reg                 LsuPlugin_logic_translationStorage_logic_sl_1_write_data_valid;
  reg        [3:0]    LsuPlugin_logic_translationStorage_logic_sl_1_write_data_virtualAddress;
  reg        [9:0]    LsuPlugin_logic_translationStorage_logic_sl_1_write_data_physicalAddress;
  reg                 LsuPlugin_logic_translationStorage_logic_sl_1_write_data_allowRead;
  reg                 LsuPlugin_logic_translationStorage_logic_sl_1_write_data_allowWrite;
  reg                 LsuPlugin_logic_translationStorage_logic_sl_1_write_data_allowExecute;
  reg                 LsuPlugin_logic_translationStorage_logic_sl_1_write_data_allowUser;
  reg                 LsuPlugin_logic_translationStorage_logic_sl_1_allocId_willIncrement;
  wire                LsuPlugin_logic_translationStorage_logic_sl_1_allocId_willClear;
  wire                LsuPlugin_logic_translationStorage_logic_sl_1_allocId_willOverflowIfInc;
  wire                LsuPlugin_logic_translationStorage_logic_sl_1_allocId_willOverflow;
  wire                MmuPlugin_logic_isMachine;
  wire                MmuPlugin_logic_isSupervisor;
  wire                MmuPlugin_logic_isUser;
  wire                when_MmuPlugin_l264;
  wire                when_MmuPlugin_l266;
  wire       [5:0]    LsuPlugin_logic_onAddress0_translationPort_logic_read_0_readAddress;
  wire       [38:0]   _zz_toplevel_execute_ctrl3_down_MMU_L0_ENTRIES_lane0_0_valid;
  wire       [38:0]   _zz_toplevel_execute_ctrl3_down_MMU_L0_ENTRIES_lane0_1_valid;
  wire       [5:0]    LsuPlugin_logic_onAddress0_translationPort_logic_read_1_readAddress;
  wire       [18:0]   _zz_toplevel_execute_ctrl3_down_MMU_L1_ENTRIES_lane0_0_valid;
  wire       [2:0]    LsuPlugin_logic_onAddress0_translationPort_logic_ctrl_hits;
  wire                LsuPlugin_logic_onAddress0_translationPort_logic_ctrl_hit;
  wire       [2:0]    _zz_LsuPlugin_logic_onAddress0_translationPort_logic_ctrl_hits_bools_0;
  wire                LsuPlugin_logic_onAddress0_translationPort_logic_ctrl_hits_bools_0;
  wire                LsuPlugin_logic_onAddress0_translationPort_logic_ctrl_hits_bools_1;
  wire                LsuPlugin_logic_onAddress0_translationPort_logic_ctrl_hits_bools_2;
  reg        [2:0]    _zz_LsuPlugin_logic_onAddress0_translationPort_logic_ctrl_oh;
  wire                LsuPlugin_logic_onAddress0_translationPort_logic_ctrl_hits_range_0_to_1;
  wire       [2:0]    LsuPlugin_logic_onAddress0_translationPort_logic_ctrl_oh;
  wire                _zz_LsuPlugin_logic_onAddress0_translationPort_logic_ctrl_lineAllowExecute;
  wire                _zz_LsuPlugin_logic_onAddress0_translationPort_logic_ctrl_lineAllowExecute_1;
  wire                _zz_LsuPlugin_logic_onAddress0_translationPort_logic_ctrl_lineAllowExecute_2;
  wire                LsuPlugin_logic_onAddress0_translationPort_logic_ctrl_lineAllowExecute;
  wire                LsuPlugin_logic_onAddress0_translationPort_logic_ctrl_lineAllowRead;
  wire                LsuPlugin_logic_onAddress0_translationPort_logic_ctrl_lineAllowWrite;
  wire                LsuPlugin_logic_onAddress0_translationPort_logic_ctrl_lineAllowUser;
  wire       [31:0]   LsuPlugin_logic_onAddress0_translationPort_logic_ctrl_lineTranslated;
  reg                 LsuPlugin_logic_onAddress0_translationPort_logic_ctrl_requireMmuLockup;
  wire       [5:0]    FetchL1Plugin_logic_translationPort_logic_read_0_readAddress;
  wire       [38:0]   _zz_fetch_logic_ctrls_1_down_MMU_L0_ENTRIES_0_valid;
  wire       [38:0]   _zz_fetch_logic_ctrls_1_down_MMU_L0_ENTRIES_1_valid;
  wire       [5:0]    FetchL1Plugin_logic_translationPort_logic_read_1_readAddress;
  wire       [18:0]   _zz_fetch_logic_ctrls_1_down_MMU_L1_ENTRIES_0_valid;
  wire       [2:0]    FetchL1Plugin_logic_translationPort_logic_ctrl_hits;
  wire                FetchL1Plugin_logic_translationPort_logic_ctrl_hit;
  wire       [2:0]    _zz_FetchL1Plugin_logic_translationPort_logic_ctrl_hits_bools_0;
  wire                FetchL1Plugin_logic_translationPort_logic_ctrl_hits_bools_0;
  wire                FetchL1Plugin_logic_translationPort_logic_ctrl_hits_bools_1;
  wire                FetchL1Plugin_logic_translationPort_logic_ctrl_hits_bools_2;
  reg        [2:0]    _zz_FetchL1Plugin_logic_translationPort_logic_ctrl_oh;
  wire                FetchL1Plugin_logic_translationPort_logic_ctrl_hits_range_0_to_1;
  wire       [2:0]    FetchL1Plugin_logic_translationPort_logic_ctrl_oh;
  wire                _zz_FetchL1Plugin_logic_translationPort_logic_ctrl_lineAllowExecute;
  wire                _zz_FetchL1Plugin_logic_translationPort_logic_ctrl_lineAllowExecute_1;
  wire                _zz_FetchL1Plugin_logic_translationPort_logic_ctrl_lineAllowExecute_2;
  wire                FetchL1Plugin_logic_translationPort_logic_ctrl_lineAllowExecute;
  wire                FetchL1Plugin_logic_translationPort_logic_ctrl_lineAllowRead;
  wire                FetchL1Plugin_logic_translationPort_logic_ctrl_lineAllowWrite;
  wire                FetchL1Plugin_logic_translationPort_logic_ctrl_lineAllowUser;
  wire       [31:0]   FetchL1Plugin_logic_translationPort_logic_ctrl_lineTranslated;
  reg                 FetchL1Plugin_logic_translationPort_logic_ctrl_requireMmuLockup;
  wire                MmuPlugin_logic_refill_wantExit;
  reg                 MmuPlugin_logic_refill_wantStart;
  wire                MmuPlugin_logic_refill_wantKill;
  wire                MmuPlugin_logic_refill_busy;
  reg        [31:0]   MmuPlugin_logic_refill_virtual;
  reg                 MmuPlugin_logic_refill_cacheRefillAny;
  reg                 MmuPlugin_logic_refill_cacheRefillAnySet;
  reg        [0:0]    MmuPlugin_logic_refill_portOhReg;
  reg        [1:0]    MmuPlugin_logic_refill_storageOhReg;
  reg        [31:0]   MmuPlugin_logic_refill_load_address;
  reg                 MmuPlugin_logic_refill_load_rsp_valid;
  reg        [31:0]   MmuPlugin_logic_refill_load_rsp_payload_data;
  reg                 MmuPlugin_logic_refill_load_rsp_payload_error;
  reg                 MmuPlugin_logic_refill_load_rsp_payload_redo;
  reg                 MmuPlugin_logic_refill_load_rsp_payload_waitAny;
  wire       [31:0]   MmuPlugin_logic_refill_load_readed;
  wire                when_MmuPlugin_l383;
  wire                MmuPlugin_logic_refill_load_flags_V;
  wire                MmuPlugin_logic_refill_load_flags_R;
  wire                MmuPlugin_logic_refill_load_flags_W;
  wire                MmuPlugin_logic_refill_load_flags_X;
  wire                MmuPlugin_logic_refill_load_flags_U;
  wire                MmuPlugin_logic_refill_load_flags_G;
  wire                MmuPlugin_logic_refill_load_flags_A;
  wire                MmuPlugin_logic_refill_load_flags_D;
  wire       [31:0]   _zz_MmuPlugin_logic_refill_load_flags_V;
  wire                MmuPlugin_logic_refill_load_leaf;
  reg                 MmuPlugin_logic_refill_load_exception;
  reg        [31:0]   MmuPlugin_logic_refill_load_levelToPhysicalAddress_0;
  reg        [31:0]   MmuPlugin_logic_refill_load_levelToPhysicalAddress_1;
  wire                MmuPlugin_logic_refill_load_levelException_0;
  reg                 MmuPlugin_logic_refill_load_levelException_1;
  reg        [31:0]   MmuPlugin_logic_refill_load_nextLevelBase;
  wire                when_MmuPlugin_l403;
  wire                MmuPlugin_logic_refill_fetch_0_pageFault;
  wire                MmuPlugin_logic_refill_fetch_0_accessFault;
  wire                MmuPlugin_logic_refill_fetch_1_pageFault;
  wire                MmuPlugin_logic_refill_fetch_1_accessFault;
  reg        [5:0]    MmuPlugin_logic_invalidate_counter;
  reg                 MmuPlugin_logic_invalidate_busy;
  wire                when_MmuPlugin_l496;
  wire                when_MmuPlugin_l510;
  wire       [7:0]    LsuTileLinkPlugin_logic_bridge_cmdHash;
  reg                 LsuTileLinkPlugin_logic_bridge_pendings_0_valid;
  reg        [7:0]    LsuTileLinkPlugin_logic_bridge_pendings_0_hash;
  reg        [3:0]    LsuTileLinkPlugin_logic_bridge_pendings_0_mask;
  reg                 LsuTileLinkPlugin_logic_bridge_pendings_0_io;
  wire                LsuTileLinkPlugin_logic_bridge_pendings_0_hazard;
  wire                LsuTileLinkPlugin_logic_bridge_hazard;
  wire                LsuTileLinkPlugin_logic_bridge_down_d_fire;
  wire                LsuTileLinkPlugin_logic_bridge_down_a_fire;
  wire                _zz_LsuPlugin_logic_bus_cmd_ready;
  wire       [2:0]    _zz_LsuTileLinkPlugin_logic_bridge_down_a_payload_opcode;
  wire                PcPlugin_logic_forcedSpawn;
  reg        [9:0]    PcPlugin_logic_harts_0_self_id;
  wire                PcPlugin_logic_harts_0_self_flow_valid;
  wire                PcPlugin_logic_harts_0_self_flow_payload_fault;
  wire       [31:0]   PcPlugin_logic_harts_0_self_flow_payload_pc;
  wire                PcPlugin_logic_harts_0_aggregator_sortedByPriority_6_laneValid;
  reg                 PcPlugin_logic_harts_0_self_increment;
  reg                 PcPlugin_logic_harts_0_self_fault;
  reg        [31:0]   PcPlugin_logic_harts_0_self_state;
  wire       [31:0]   PcPlugin_logic_harts_0_self_pc;
  wire                PcPlugin_logic_harts_0_aggregator_valids_0;
  wire                PcPlugin_logic_harts_0_aggregator_valids_1;
  wire                PcPlugin_logic_harts_0_aggregator_valids_2;
  wire                PcPlugin_logic_harts_0_aggregator_valids_3;
  wire                PcPlugin_logic_harts_0_aggregator_valids_4;
  wire                PcPlugin_logic_harts_0_aggregator_valids_5;
  wire                PcPlugin_logic_harts_0_aggregator_valids_6;
  wire       [6:0]    _zz_PcPlugin_logic_harts_0_aggregator_oh;
  wire                _zz_PcPlugin_logic_harts_0_aggregator_oh_1;
  wire                _zz_PcPlugin_logic_harts_0_aggregator_oh_2;
  wire                _zz_PcPlugin_logic_harts_0_aggregator_oh_3;
  wire                _zz_PcPlugin_logic_harts_0_aggregator_oh_4;
  wire                _zz_PcPlugin_logic_harts_0_aggregator_oh_5;
  wire                _zz_PcPlugin_logic_harts_0_aggregator_oh_6;
  reg        [6:0]    _zz_PcPlugin_logic_harts_0_aggregator_oh_7;
  wire                _zz_PcPlugin_logic_harts_0_aggregator_oh_8;
  wire       [6:0]    PcPlugin_logic_harts_0_aggregator_oh;
  wire       [31:0]   PcPlugin_logic_harts_0_aggregator_target;
  wire                PcPlugin_logic_harts_0_aggregator_fault;
  wire                _zz_PcPlugin_logic_harts_0_aggregator_target;
  wire                _zz_PcPlugin_logic_harts_0_aggregator_target_1;
  wire                _zz_PcPlugin_logic_harts_0_aggregator_target_2;
  wire                _zz_PcPlugin_logic_harts_0_aggregator_target_3;
  wire                _zz_PcPlugin_logic_harts_0_aggregator_target_4;
  wire                _zz_PcPlugin_logic_harts_0_aggregator_target_5;
  wire                _zz_PcPlugin_logic_harts_0_aggregator_target_6;
  wire                PcPlugin_logic_harts_0_holdComb;
  reg                 PcPlugin_logic_harts_0_holdReg;
  wire                PcPlugin_logic_harts_0_output_valid;
  wire                PcPlugin_logic_harts_0_output_ready;
  reg        [31:0]   PcPlugin_logic_harts_0_output_payload_pc;
  wire                PcPlugin_logic_harts_0_output_payload_fault;
  wire                PcPlugin_logic_harts_0_output_fire;
  wire                PcPlugin_logic_holdHalter_doIt;
  wire                fetch_logic_ctrls_0_haltRequest_PcPlugin_l136;
  wire                CsrAccessPlugin_logic_fsm_wantExit;
  reg                 CsrAccessPlugin_logic_fsm_wantStart;
  wire                CsrAccessPlugin_logic_fsm_wantKill;
  reg                 REG_CSR_1952;
  reg                 REG_CSR_1953;
  reg                 REG_CSR_1954;
  reg                 REG_CSR_3857;
  reg                 REG_CSR_3858;
  reg                 REG_CSR_3859;
  reg                 REG_CSR_3860;
  reg                 REG_CSR_769;
  reg                 REG_CSR_768;
  reg                 REG_CSR_834;
  reg                 REG_CSR_836;
  reg                 REG_CSR_772;
  reg                 REG_CSR_770;
  reg                 REG_CSR_771;
  reg                 REG_CSR_322;
  reg                 REG_CSR_256;
  reg                 REG_CSR_260;
  reg                 REG_CSR_324;
  reg                 REG_CSR_3073;
  reg                 REG_CSR_3201;
  reg                 REG_CSR_PrivilegedPlugin_logic_readAnyWriteLegal_tvecFilter;
  reg                 REG_CSR_PrivilegedPlugin_logic_readAnyWriteLegal_epcFilter;
  reg                 REG_CSR_384;
  reg                 REG_CSR_CsrRamPlugin_csrMapper_selFilter;
  reg                 REG_CSR_CsrAccessPlugin_logic_trapNextOnWriteFilter;
  reg                 CsrAccessPlugin_logic_fsm_regs_read;
  reg                 CsrAccessPlugin_logic_fsm_regs_write;
  wire       [31:0]   CsrAccessPlugin_logic_fsm_regs_rs1;
  reg        [31:0]   CsrAccessPlugin_logic_fsm_regs_aluInput;
  reg        [31:0]   CsrAccessPlugin_logic_fsm_regs_csrValue;
  reg        [31:0]   CsrAccessPlugin_logic_fsm_regs_onWriteBits;
  wire       [15:0]   CsrAccessPlugin_logic_fsm_regs_uopId;
  wire       [31:0]   CsrAccessPlugin_logic_fsm_regs_uop;
  wire                CsrAccessPlugin_logic_fsm_regs_doImm;
  wire                CsrAccessPlugin_logic_fsm_regs_doMask;
  wire                CsrAccessPlugin_logic_fsm_regs_doClear;
  wire       [4:0]    CsrAccessPlugin_logic_fsm_regs_rdPhys;
  wire                CsrAccessPlugin_logic_fsm_regs_rdEnable;
  reg                 CsrAccessPlugin_logic_fsm_regs_fire;
  wire       [11:0]   CsrAccessPlugin_logic_fsm_inject_csrAddress;
  wire                CsrAccessPlugin_logic_fsm_inject_immZero;
  wire                CsrAccessPlugin_logic_fsm_inject_srcZero;
  wire                CsrAccessPlugin_logic_fsm_inject_csrWrite;
  wire                CsrAccessPlugin_logic_fsm_inject_csrRead;
  wire                COMB_CSR_1952;
  wire                COMB_CSR_1953;
  wire                COMB_CSR_1954;
  wire                COMB_CSR_3857;
  wire                COMB_CSR_3858;
  wire                COMB_CSR_3859;
  wire                COMB_CSR_3860;
  wire                COMB_CSR_769;
  wire                COMB_CSR_768;
  wire                COMB_CSR_834;
  wire                COMB_CSR_836;
  wire                COMB_CSR_772;
  wire                COMB_CSR_770;
  wire                COMB_CSR_771;
  wire                COMB_CSR_322;
  wire                COMB_CSR_256;
  wire                COMB_CSR_260;
  wire                COMB_CSR_324;
  wire                COMB_CSR_3073;
  wire                COMB_CSR_3201;
  wire                COMB_CSR_PrivilegedPlugin_logic_readAnyWriteLegal_tvecFilter;
  wire                COMB_CSR_PrivilegedPlugin_logic_readAnyWriteLegal_epcFilter;
  wire                COMB_CSR_384;
  wire                COMB_CSR_CsrRamPlugin_csrMapper_selFilter;
  wire                COMB_CSR_CsrAccessPlugin_logic_trapNextOnWriteFilter;
  wire                CsrAccessPlugin_logic_fsm_inject_implemented;
  wire                CsrAccessPlugin_logic_fsm_inject_onDecodeDo;
  wire                when_CsrAccessPlugin_l155;
  wire                when_MmuPlugin_l212;
  wire                when_CsrAccessPlugin_l155_1;
  wire                CsrAccessPlugin_logic_fsm_inject_trap;
  reg                 CsrAccessPlugin_logic_fsm_inject_unfreeze;
  wire                CsrAccessPlugin_logic_fsm_inject_iLogic_freeze;
  reg                 CsrAccessPlugin_logic_fsm_inject_flushReg;
  wire                when_CsrAccessPlugin_l209;
  reg                 CsrAccessPlugin_logic_fsm_inject_sampled;
  reg                 CsrAccessPlugin_logic_fsm_inject_trapReg;
  reg                 CsrAccessPlugin_logic_fsm_inject_busTrapReg;
  reg        [3:0]    CsrAccessPlugin_logic_fsm_inject_busTrapCodeReg;
  reg                 CsrAccessPlugin_logic_fsm_readLogic_onReadsDo;
  reg                 CsrAccessPlugin_logic_fsm_readLogic_onReadsFireDo;
  wire                when_CsrAccessPlugin_l264;
  wire       [31:0]   CsrAccessPlugin_logic_fsm_readLogic_csrValue;
  wire                when_CsrAccessPlugin_l291;
  wire       [31:0]   CsrAccessPlugin_logic_fsm_writeLogic_alu_mask;
  wire       [31:0]   CsrAccessPlugin_logic_fsm_writeLogic_alu_masked;
  wire       [31:0]   CsrAccessPlugin_logic_fsm_writeLogic_alu_result;
  reg                 CsrAccessPlugin_logic_fsm_writeLogic_onWritesDo;
  reg                 CsrAccessPlugin_logic_fsm_writeLogic_onWritesFireDo;
  wire                when_CsrAccessPlugin_l359;
  wire       [1:0]    switch_PrivilegedPlugin_l540;
  wire                when_CsrAccessPlugin_l359_1;
  wire                when_CsrAccessPlugin_l359_2;
  wire                when_CsrAccessPlugin_l359_3;
  wire                when_CsrAccessPlugin_l359_4;
  wire                when_CsrAccessPlugin_l359_5;
  wire                when_CsrAccessPlugin_l359_6;
  wire                when_CsrAccessPlugin_l359_7;
  wire                when_CsrAccessPlugin_l359_8;
  wire                when_CsrAccessPlugin_l359_9;
  wire                when_CsrAccessPlugin_l356;
  wire                when_CsrAccessPlugin_l356_1;
  wire                when_CsrAccessPlugin_l366;
  wire                when_CsrAccessPlugin_l359_10;
  wire                when_CsrAccessPlugin_l356_2;
  reg                 CsrAccessPlugin_logic_fsm_completion_valid;
  wire       [15:0]   CsrAccessPlugin_logic_fsm_completion_payload_uopId;
  wire                CsrAccessPlugin_logic_fsm_completion_payload_trap;
  wire                CsrAccessPlugin_logic_fsm_completion_payload_commit;
  reg        [11:0]   HistoryPlugin_logic_onFetch_value;
  reg        [11:0]   HistoryPlugin_logic_onFetch_valueNext;
  wire                HistoryPlugin_logic_onFetch_ports_0_valid;
  wire       [11:0]   HistoryPlugin_logic_onFetch_ports_0_payload_history;
  wire                HistoryPlugin_logic_onFetch_ports_1_valid;
  wire       [11:0]   HistoryPlugin_logic_onFetch_ports_1_payload_history;
  wire       [0:0]    HistoryPlugin_logic_onFetch_ports_1_payload_age;
  wire       [12:0]   _zz_HistoryPlugin_logic_onFetch_ports_1_payload_history;
  wire                HistoryPlugin_logic_onFetch_ports_2_valid;
  wire       [11:0]   HistoryPlugin_logic_onFetch_ports_2_payload_history;
  wire       [0:0]    HistoryPlugin_logic_onFetch_ports_2_payload_age;
  wire       [12:0]   _zz_HistoryPlugin_logic_onFetch_ports_2_payload_history;
  wire                HistoryPlugin_logic_onFetch_ports_3_valid;
  wire       [11:0]   HistoryPlugin_logic_onFetch_ports_3_payload_history;
  wire       [2:0]    CsrRamPlugin_logic_writeLogic_hits;
  wire                CsrRamPlugin_logic_writeLogic_hit;
  wire       [2:0]    CsrRamPlugin_logic_writeLogic_hits_ohFirst_input;
  wire       [2:0]    CsrRamPlugin_logic_writeLogic_hits_ohFirst_masked;
  wire       [2:0]    CsrRamPlugin_logic_writeLogic_oh;
  wire                CsrRamPlugin_logic_writeLogic_port_valid;
  wire       [2:0]    CsrRamPlugin_logic_writeLogic_port_payload_address;
  wire       [31:0]   CsrRamPlugin_logic_writeLogic_port_payload_data;
  wire                _zz_TrapPlugin_logic_harts_0_crsPorts_write_ready;
  wire                _zz_CsrRamPlugin_csrMapper_write_ready;
  wire                _zz_CsrRamPlugin_setup_initPort_ready;
  wire       [1:0]    CsrRamPlugin_logic_readLogic_hits;
  wire                CsrRamPlugin_logic_readLogic_hit;
  wire       [1:0]    CsrRamPlugin_logic_readLogic_hits_ohFirst_input;
  wire       [1:0]    CsrRamPlugin_logic_readLogic_hits_ohFirst_masked;
  wire       [1:0]    CsrRamPlugin_logic_readLogic_oh;
  wire                _zz_CsrRamPlugin_logic_readLogic_sel;
  wire       [0:0]    CsrRamPlugin_logic_readLogic_sel;
  wire                CsrRamPlugin_logic_readLogic_port_cmd_valid;
  wire       [2:0]    CsrRamPlugin_logic_readLogic_port_cmd_payload;
  wire       [31:0]   CsrRamPlugin_logic_readLogic_port_rsp;
  reg        [1:0]    CsrRamPlugin_logic_readLogic_ohReg;
  reg                 CsrRamPlugin_logic_readLogic_busy;
  reg        [3:0]    CsrRamPlugin_logic_flush_counter;
  wire                CsrRamPlugin_logic_flush_done;
  wire                toplevel_execute_lane0_bypasser_integer_RS1_port_valid;
  wire       [4:0]    toplevel_execute_lane0_bypasser_integer_RS1_port_address;
  wire       [31:0]   toplevel_execute_lane0_bypasser_integer_RS1_port_data;
  reg        [8:0]    toplevel_execute_lane0_bypasser_integer_RS1_bypassEnables;
  wire       [8:0]    _zz_toplevel_execute_lane0_bypasser_integer_RS1_bypassEnables_bools_0;
  wire                toplevel_execute_lane0_bypasser_integer_RS1_bypassEnables_bools_0;
  wire                toplevel_execute_lane0_bypasser_integer_RS1_bypassEnables_bools_1;
  wire                toplevel_execute_lane0_bypasser_integer_RS1_bypassEnables_bools_2;
  wire                toplevel_execute_lane0_bypasser_integer_RS1_bypassEnables_bools_3;
  wire                toplevel_execute_lane0_bypasser_integer_RS1_bypassEnables_bools_4;
  wire                toplevel_execute_lane0_bypasser_integer_RS1_bypassEnables_bools_5;
  wire                toplevel_execute_lane0_bypasser_integer_RS1_bypassEnables_bools_6;
  wire                toplevel_execute_lane0_bypasser_integer_RS1_bypassEnables_bools_7;
  wire                toplevel_execute_lane0_bypasser_integer_RS1_bypassEnables_bools_8;
  reg        [8:0]    _zz_toplevel_execute_lane0_bypasser_integer_RS1_sel;
  wire                toplevel_execute_lane0_bypasser_integer_RS1_bypassEnables_range_0_to_1;
  wire                toplevel_execute_lane0_bypasser_integer_RS1_bypassEnables_range_0_to_2;
  wire                toplevel_execute_lane0_bypasser_integer_RS1_bypassEnables_range_0_to_3;
  wire                toplevel_execute_lane0_bypasser_integer_RS1_bypassEnables_range_4_to_5;
  wire                toplevel_execute_lane0_bypasser_integer_RS1_bypassEnables_range_4_to_6;
  wire                toplevel_execute_lane0_bypasser_integer_RS1_bypassEnables_range_4_to_7;
  wire       [8:0]    toplevel_execute_lane0_bypasser_integer_RS1_sel;
  wire       [7:0]    _zz_toplevel_execute_ctrl1_down_integer_RS1_lane0;
  (* keep , syn_keep *) reg        [31:0]   _zz_toplevel_execute_ctrl1_down_integer_RS1_lane0_1 /* synthesis syn_keep = 1 */ ;
  wire                when_ExecuteLanePlugin_l190;
  wire                toplevel_execute_lane0_bypasser_integer_RS1_along_bypasses_0_checks_0_selfHit;
  wire                toplevel_execute_lane0_bypasser_integer_RS1_along_bypasses_0_checks_0_hit;
  wire                toplevel_execute_lane0_bypasser_integer_RS1_along_bypasses_0_checks_1_selfHit;
  wire                toplevel_execute_lane0_bypasser_integer_RS1_along_bypasses_0_checks_1_youngerHits_0;
  wire                toplevel_execute_lane0_bypasser_integer_RS1_along_bypasses_0_checks_1_youngerHits_1;
  wire                toplevel_execute_lane0_bypasser_integer_RS1_along_bypasses_0_checks_1_hit;
  wire                toplevel_execute_lane0_bypasser_integer_RS1_along_bypasses_0_checks_2_selfHit;
  wire                toplevel_execute_lane0_bypasser_integer_RS1_along_bypasses_0_checks_2_hit;
  wire                toplevel_execute_lane0_bypasser_integer_RS1_along_bypasses_0_checks_3_selfHit;
  wire                toplevel_execute_lane0_bypasser_integer_RS1_along_bypasses_0_checks_3_youngerHits_0;
  wire                toplevel_execute_lane0_bypasser_integer_RS1_along_bypasses_0_checks_3_youngerHits_1;
  wire                toplevel_execute_lane0_bypasser_integer_RS1_along_bypasses_0_checks_3_hit;
  wire       [3:0]    toplevel_execute_lane0_bypasser_integer_RS1_along_bypasses_0_hits;
  wire       [4:0]    _zz_toplevel_execute_ctrl2_integer_RS1_lane0_bypass;
  wire                toplevel_execute_lane0_bypasser_integer_RS1_along_bypasses_1_checks_0_selfHit;
  wire                toplevel_execute_lane0_bypasser_integer_RS1_along_bypasses_1_checks_0_hit;
  wire                toplevel_execute_lane0_bypasser_integer_RS1_along_bypasses_1_checks_1_selfHit;
  wire                toplevel_execute_lane0_bypasser_integer_RS1_along_bypasses_1_checks_1_hit;
  wire       [1:0]    toplevel_execute_lane0_bypasser_integer_RS1_along_bypasses_1_hits;
  wire       [2:0]    _zz_toplevel_execute_ctrl3_integer_RS1_lane0_bypass;
  wire                toplevel_execute_lane0_bypasser_integer_RS2_port_valid;
  wire       [4:0]    toplevel_execute_lane0_bypasser_integer_RS2_port_address;
  wire       [31:0]   toplevel_execute_lane0_bypasser_integer_RS2_port_data;
  reg        [8:0]    toplevel_execute_lane0_bypasser_integer_RS2_bypassEnables;
  wire       [8:0]    _zz_toplevel_execute_lane0_bypasser_integer_RS2_bypassEnables_bools_0;
  wire                toplevel_execute_lane0_bypasser_integer_RS2_bypassEnables_bools_0;
  wire                toplevel_execute_lane0_bypasser_integer_RS2_bypassEnables_bools_1;
  wire                toplevel_execute_lane0_bypasser_integer_RS2_bypassEnables_bools_2;
  wire                toplevel_execute_lane0_bypasser_integer_RS2_bypassEnables_bools_3;
  wire                toplevel_execute_lane0_bypasser_integer_RS2_bypassEnables_bools_4;
  wire                toplevel_execute_lane0_bypasser_integer_RS2_bypassEnables_bools_5;
  wire                toplevel_execute_lane0_bypasser_integer_RS2_bypassEnables_bools_6;
  wire                toplevel_execute_lane0_bypasser_integer_RS2_bypassEnables_bools_7;
  wire                toplevel_execute_lane0_bypasser_integer_RS2_bypassEnables_bools_8;
  reg        [8:0]    _zz_toplevel_execute_lane0_bypasser_integer_RS2_sel;
  wire                toplevel_execute_lane0_bypasser_integer_RS2_bypassEnables_range_0_to_1;
  wire                toplevel_execute_lane0_bypasser_integer_RS2_bypassEnables_range_0_to_2;
  wire                toplevel_execute_lane0_bypasser_integer_RS2_bypassEnables_range_0_to_3;
  wire                toplevel_execute_lane0_bypasser_integer_RS2_bypassEnables_range_4_to_5;
  wire                toplevel_execute_lane0_bypasser_integer_RS2_bypassEnables_range_4_to_6;
  wire                toplevel_execute_lane0_bypasser_integer_RS2_bypassEnables_range_4_to_7;
  wire       [8:0]    toplevel_execute_lane0_bypasser_integer_RS2_sel;
  wire       [7:0]    _zz_toplevel_execute_ctrl1_down_integer_RS2_lane0;
  (* keep , syn_keep *) reg        [31:0]   _zz_toplevel_execute_ctrl1_down_integer_RS2_lane0_1 /* synthesis syn_keep = 1 */ ;
  wire                when_ExecuteLanePlugin_l190_1;
  wire                toplevel_execute_lane0_bypasser_integer_RS2_along_bypasses_0_checks_0_selfHit;
  wire                toplevel_execute_lane0_bypasser_integer_RS2_along_bypasses_0_checks_0_hit;
  wire                toplevel_execute_lane0_bypasser_integer_RS2_along_bypasses_0_checks_1_selfHit;
  wire                toplevel_execute_lane0_bypasser_integer_RS2_along_bypasses_0_checks_1_youngerHits_0;
  wire                toplevel_execute_lane0_bypasser_integer_RS2_along_bypasses_0_checks_1_youngerHits_1;
  wire                toplevel_execute_lane0_bypasser_integer_RS2_along_bypasses_0_checks_1_hit;
  wire                toplevel_execute_lane0_bypasser_integer_RS2_along_bypasses_0_checks_2_selfHit;
  wire                toplevel_execute_lane0_bypasser_integer_RS2_along_bypasses_0_checks_2_hit;
  wire                toplevel_execute_lane0_bypasser_integer_RS2_along_bypasses_0_checks_3_selfHit;
  wire                toplevel_execute_lane0_bypasser_integer_RS2_along_bypasses_0_checks_3_youngerHits_0;
  wire                toplevel_execute_lane0_bypasser_integer_RS2_along_bypasses_0_checks_3_youngerHits_1;
  wire                toplevel_execute_lane0_bypasser_integer_RS2_along_bypasses_0_checks_3_hit;
  wire       [3:0]    toplevel_execute_lane0_bypasser_integer_RS2_along_bypasses_0_hits;
  wire       [4:0]    _zz_toplevel_execute_ctrl2_integer_RS2_lane0_bypass;
  wire                toplevel_execute_lane0_bypasser_integer_RS2_along_bypasses_1_checks_0_selfHit;
  wire                toplevel_execute_lane0_bypasser_integer_RS2_along_bypasses_1_checks_0_hit;
  wire                toplevel_execute_lane0_bypasser_integer_RS2_along_bypasses_1_checks_1_selfHit;
  wire                toplevel_execute_lane0_bypasser_integer_RS2_along_bypasses_1_checks_1_hit;
  wire       [1:0]    toplevel_execute_lane0_bypasser_integer_RS2_along_bypasses_1_hits;
  wire       [2:0]    _zz_toplevel_execute_ctrl3_integer_RS2_lane0_bypass;
  wire                execute_lane0_logic_completions_onCtrl_0_port_valid;
  wire       [15:0]   execute_lane0_logic_completions_onCtrl_0_port_payload_uopId;
  wire                execute_lane0_logic_completions_onCtrl_0_port_payload_trap;
  wire                execute_lane0_logic_completions_onCtrl_0_port_payload_commit;
  wire                execute_lane0_logic_completions_onCtrl_1_port_valid;
  wire       [15:0]   execute_lane0_logic_completions_onCtrl_1_port_payload_uopId;
  wire                execute_lane0_logic_completions_onCtrl_1_port_payload_trap;
  wire                execute_lane0_logic_completions_onCtrl_1_port_payload_commit;
  wire                execute_lane0_logic_completions_onCtrl_2_port_valid;
  wire       [15:0]   execute_lane0_logic_completions_onCtrl_2_port_payload_uopId;
  wire                execute_lane0_logic_completions_onCtrl_2_port_payload_trap;
  wire                execute_lane0_logic_completions_onCtrl_2_port_payload_commit;
  wire       [32:0]   execute_lane0_logic_decoding_decodingBits;
  wire                _zz_toplevel_execute_ctrl1_down_execute_lane0_logic_completions_onCtrl_0_ENABLE_lane0;
  wire                _zz_toplevel_execute_ctrl1_down_execute_lane0_logic_completions_onCtrl_0_ENABLE_lane0_1;
  wire                _zz_toplevel_execute_ctrl1_down_execute_lane0_logic_completions_onCtrl_0_ENABLE_lane0_2;
  wire                _zz_toplevel_execute_ctrl1_down_execute_lane0_logic_completions_onCtrl_0_ENABLE_lane0_3;
  wire                _zz_toplevel_execute_ctrl1_down_execute_lane0_logic_completions_onCtrl_1_ENABLE_lane0;
  wire                _zz_toplevel_execute_ctrl1_down_execute_lane0_logic_completions_onCtrl_1_ENABLE_lane0_1;
  wire                _zz_toplevel_execute_ctrl1_down_execute_lane0_logic_completions_onCtrl_1_ENABLE_lane0_2;
  wire                _zz_toplevel_execute_ctrl1_down_execute_lane0_logic_completions_onCtrl_0_ENABLE_lane0_4;
  wire                _zz_toplevel_execute_ctrl1_down_late0_BranchPlugin_SEL_lane0;
  wire                _zz_toplevel_execute_ctrl1_down_execute_lane0_logic_completions_onCtrl_2_ENABLE_lane0;
  wire                _zz_toplevel_execute_ctrl1_down_execute_lane0_logic_completions_onCtrl_2_ENABLE_lane0_1;
  wire                _zz_toplevel_execute_ctrl1_down_AguPlugin_LOAD_lane0;
  wire                _zz_toplevel_execute_ctrl1_down_lane0_integer_WriteBackPlugin_SEL_lane0;
  wire                _zz_toplevel_execute_ctrl1_down_AguPlugin_ATOMIC_lane0;
  wire                _zz_toplevel_execute_ctrl1_down_execute_lane0_logic_completions_onCtrl_0_ENABLE_lane0_5;
  wire                _zz_toplevel_execute_ctrl1_down_execute_lane0_logic_completions_onCtrl_0_ENABLE_lane0_6;
  wire                _zz_toplevel_execute_ctrl1_down_execute_lane0_logic_completions_onCtrl_1_ENABLE_lane0_3;
  wire                _zz_toplevel_execute_ctrl1_down_execute_lane0_logic_completions_onCtrl_1_ENABLE_lane0_4;
  wire                _zz_toplevel_execute_ctrl1_down_execute_lane0_logic_completions_onCtrl_1_ENABLE_lane0_5;
  wire                _zz_toplevel_execute_ctrl1_down_execute_lane0_logic_completions_onCtrl_2_ENABLE_lane0_2;
  wire                _zz_toplevel_execute_ctrl1_down_execute_lane0_logic_completions_onCtrl_2_ENABLE_lane0_3;
  wire                _zz_toplevel_execute_ctrl1_down_late0_IntAluPlugin_ALU_ADD_SUB_lane0;
  wire                _zz_toplevel_execute_ctrl1_down_late0_SrcPlugin_logic_SRC2_CTRL_lane0;
  wire                _zz_toplevel_execute_ctrl1_down_late0_IntAluPlugin_ALU_SLTX_lane0;
  wire                _zz_toplevel_execute_ctrl1_down_late0_IntAluPlugin_ALU_BITWISE_CTRL_lane0;
  wire                _zz_toplevel_execute_ctrl1_down_BarrelShifterPlugin_LEFT_lane0;
  wire                _zz_toplevel_execute_ctrl1_down_CsrAccessPlugin_CSR_CLEAR_lane0;
  wire       [1:0]    _zz_toplevel_execute_ctrl1_down_early0_IntAluPlugin_ALU_BITWISE_CTRL_lane0;
  wire       [1:0]    _zz_toplevel_execute_ctrl1_down_early0_IntAluPlugin_ALU_BITWISE_CTRL_lane0_1;
  wire       [1:0]    _zz_toplevel_execute_ctrl1_down_early0_IntAluPlugin_ALU_BITWISE_CTRL_lane0_2;
  wire                _zz_toplevel_execute_ctrl1_down_late0_SrcPlugin_logic_SRC2_CTRL_lane0_1;
  wire                _zz_toplevel_execute_ctrl1_down_AguPlugin_STORE_lane0;
  wire                _zz_toplevel_execute_ctrl1_down_BYPASSED_AT_3_lane0;
  wire                _zz_toplevel_execute_ctrl1_down_SrcStageables_UNSIGNED_lane0;
  wire       [1:0]    _zz_toplevel_execute_ctrl1_down_BranchPlugin_BRANCH_CTRL_lane0;
  wire       [1:0]    _zz_toplevel_execute_ctrl1_down_BranchPlugin_BRANCH_CTRL_lane0_1;
  wire       [1:0]    _zz_toplevel_execute_ctrl1_down_BranchPlugin_BRANCH_CTRL_lane0_2;
  wire                _zz_toplevel_execute_ctrl1_down_CsrAccessPlugin_CSR_MASK_lane0;
  wire                _zz_toplevel_execute_ctrl1_down_early0_EnvPlugin_OP_lane0;
  wire       [2:0]    _zz_toplevel_execute_ctrl1_down_early0_EnvPlugin_OP_lane0_1;
  wire       [2:0]    _zz_toplevel_execute_ctrl1_down_early0_EnvPlugin_OP_lane0_2;
  wire       [2:0]    _zz_toplevel_execute_ctrl1_down_early0_EnvPlugin_OP_lane0_3;
  wire       [1:0]    _zz_toplevel_execute_ctrl1_down_late0_IntAluPlugin_ALU_BITWISE_CTRL_lane0_1;
  wire       [1:0]    _zz_toplevel_execute_ctrl1_down_late0_IntAluPlugin_ALU_BITWISE_CTRL_lane0_2;
  wire       [1:0]    _zz_toplevel_execute_ctrl1_down_late0_IntAluPlugin_ALU_BITWISE_CTRL_lane0_3;
  wire                when_ExecuteLanePlugin_l300;
  wire                when_ExecuteLanePlugin_l300_1;
  wire                when_ExecuteLanePlugin_l300_2;
  wire                when_ExecuteLanePlugin_l300_3;
  wire                when_ExecuteLanePlugin_l300_4;
  wire                WhiteboxerPlugin_logic_csr_port_valid;
  wire       [15:0]   WhiteboxerPlugin_logic_csr_port_payload_uopId;
  wire       [11:0]   WhiteboxerPlugin_logic_csr_port_payload_address;
  wire       [31:0]   WhiteboxerPlugin_logic_csr_port_payload_write;
  wire       [31:0]   WhiteboxerPlugin_logic_csr_port_payload_read;
  wire                WhiteboxerPlugin_logic_csr_port_payload_writeDone;
  wire                WhiteboxerPlugin_logic_csr_port_payload_readDone;
  wire                WhiteboxerPlugin_logic_rfWrites_ports_0_valid;
  wire       [15:0]   WhiteboxerPlugin_logic_rfWrites_ports_0_payload_uopId;
  wire       [31:0]   WhiteboxerPlugin_logic_rfWrites_ports_0_payload_data;
  wire                WhiteboxerPlugin_logic_rfWrites_ports_1_valid;
  wire       [15:0]   WhiteboxerPlugin_logic_rfWrites_ports_1_payload_uopId;
  wire       [31:0]   WhiteboxerPlugin_logic_rfWrites_ports_1_payload_data;
  wire                WhiteboxerPlugin_logic_rfWrites_ports_2_valid;
  wire       [15:0]   WhiteboxerPlugin_logic_rfWrites_ports_2_payload_uopId;
  wire       [31:0]   WhiteboxerPlugin_logic_rfWrites_ports_2_payload_data;
  wire                WhiteboxerPlugin_logic_rfWrites_ports_3_valid;
  wire       [15:0]   WhiteboxerPlugin_logic_rfWrites_ports_3_payload_uopId;
  wire       [31:0]   WhiteboxerPlugin_logic_rfWrites_ports_3_payload_data;
  wire                WhiteboxerPlugin_logic_rfWrites_ports_4_valid;
  wire       [15:0]   WhiteboxerPlugin_logic_rfWrites_ports_4_payload_uopId;
  wire       [31:0]   WhiteboxerPlugin_logic_rfWrites_ports_4_payload_data;
  wire                WhiteboxerPlugin_logic_rfWrites_ports_5_valid;
  wire       [15:0]   WhiteboxerPlugin_logic_rfWrites_ports_5_payload_uopId;
  wire       [31:0]   WhiteboxerPlugin_logic_rfWrites_ports_5_payload_data;
  wire                WhiteboxerPlugin_logic_completions_ports_0_valid;
  wire       [15:0]   WhiteboxerPlugin_logic_completions_ports_0_payload_uopId;
  wire                WhiteboxerPlugin_logic_completions_ports_0_payload_trap;
  wire                WhiteboxerPlugin_logic_completions_ports_0_payload_commit;
  wire                WhiteboxerPlugin_logic_completions_ports_1_valid;
  wire       [15:0]   WhiteboxerPlugin_logic_completions_ports_1_payload_uopId;
  wire                WhiteboxerPlugin_logic_completions_ports_1_payload_trap;
  wire                WhiteboxerPlugin_logic_completions_ports_1_payload_commit;
  wire                WhiteboxerPlugin_logic_completions_ports_2_valid;
  wire       [15:0]   WhiteboxerPlugin_logic_completions_ports_2_payload_uopId;
  wire                WhiteboxerPlugin_logic_completions_ports_2_payload_trap;
  wire                WhiteboxerPlugin_logic_completions_ports_2_payload_commit;
  wire                WhiteboxerPlugin_logic_completions_ports_3_valid;
  wire       [15:0]   WhiteboxerPlugin_logic_completions_ports_3_payload_uopId;
  wire                WhiteboxerPlugin_logic_completions_ports_3_payload_trap;
  wire                WhiteboxerPlugin_logic_completions_ports_3_payload_commit;
  wire                WhiteboxerPlugin_logic_completions_ports_4_valid;
  wire       [15:0]   WhiteboxerPlugin_logic_completions_ports_4_payload_uopId;
  wire                WhiteboxerPlugin_logic_completions_ports_4_payload_trap;
  wire                WhiteboxerPlugin_logic_completions_ports_4_payload_commit;
  wire                fetch_logic_flushes_0_doIt;
  wire                fetch_logic_ctrls_1_throwWhen_FetchPipelinePlugin_l44;
  wire                fetch_logic_flushes_1_doIt;
  wire                fetch_logic_ctrls_2_forgetsSingleRequest_FetchPipelinePlugin_l46;
  reg        [8:0]    toplevel_execute_lane1_bypasser_integer_RS1_bypassEnables;
  wire       [8:0]    _zz_toplevel_execute_lane1_bypasser_integer_RS1_bypassEnables_bools_0;
  wire                toplevel_execute_lane1_bypasser_integer_RS1_bypassEnables_bools_0;
  wire                toplevel_execute_lane1_bypasser_integer_RS1_bypassEnables_bools_1;
  wire                toplevel_execute_lane1_bypasser_integer_RS1_bypassEnables_bools_2;
  wire                toplevel_execute_lane1_bypasser_integer_RS1_bypassEnables_bools_3;
  wire                toplevel_execute_lane1_bypasser_integer_RS1_bypassEnables_bools_4;
  wire                toplevel_execute_lane1_bypasser_integer_RS1_bypassEnables_bools_5;
  wire                toplevel_execute_lane1_bypasser_integer_RS1_bypassEnables_bools_6;
  wire                toplevel_execute_lane1_bypasser_integer_RS1_bypassEnables_bools_7;
  wire                toplevel_execute_lane1_bypasser_integer_RS1_bypassEnables_bools_8;
  reg        [8:0]    _zz_toplevel_execute_lane1_bypasser_integer_RS1_sel;
  wire                toplevel_execute_lane1_bypasser_integer_RS1_bypassEnables_range_0_to_1;
  wire                toplevel_execute_lane1_bypasser_integer_RS1_bypassEnables_range_0_to_2;
  wire                toplevel_execute_lane1_bypasser_integer_RS1_bypassEnables_range_0_to_3;
  wire                toplevel_execute_lane1_bypasser_integer_RS1_bypassEnables_range_4_to_5;
  wire                toplevel_execute_lane1_bypasser_integer_RS1_bypassEnables_range_4_to_6;
  wire                toplevel_execute_lane1_bypasser_integer_RS1_bypassEnables_range_4_to_7;
  wire       [8:0]    toplevel_execute_lane1_bypasser_integer_RS1_sel;
  wire       [7:0]    _zz_toplevel_execute_ctrl1_down_integer_RS1_lane1;
  (* keep , syn_keep *) reg        [31:0]   _zz_toplevel_execute_ctrl1_down_integer_RS1_lane1_1 /* synthesis syn_keep = 1 */ ;
  wire                when_ExecuteLanePlugin_l190_2;
  wire                toplevel_execute_lane1_bypasser_integer_RS1_along_bypasses_0_checks_0_selfHit;
  wire                toplevel_execute_lane1_bypasser_integer_RS1_along_bypasses_0_checks_0_hit;
  wire                toplevel_execute_lane1_bypasser_integer_RS1_along_bypasses_0_checks_1_selfHit;
  wire                toplevel_execute_lane1_bypasser_integer_RS1_along_bypasses_0_checks_1_youngerHits_0;
  wire                toplevel_execute_lane1_bypasser_integer_RS1_along_bypasses_0_checks_1_youngerHits_1;
  wire                toplevel_execute_lane1_bypasser_integer_RS1_along_bypasses_0_checks_1_hit;
  wire                toplevel_execute_lane1_bypasser_integer_RS1_along_bypasses_0_checks_2_selfHit;
  wire                toplevel_execute_lane1_bypasser_integer_RS1_along_bypasses_0_checks_2_hit;
  wire                toplevel_execute_lane1_bypasser_integer_RS1_along_bypasses_0_checks_3_selfHit;
  wire                toplevel_execute_lane1_bypasser_integer_RS1_along_bypasses_0_checks_3_youngerHits_0;
  wire                toplevel_execute_lane1_bypasser_integer_RS1_along_bypasses_0_checks_3_youngerHits_1;
  wire                toplevel_execute_lane1_bypasser_integer_RS1_along_bypasses_0_checks_3_hit;
  wire       [3:0]    toplevel_execute_lane1_bypasser_integer_RS1_along_bypasses_0_hits;
  wire       [4:0]    _zz_toplevel_execute_ctrl2_integer_RS1_lane1_bypass;
  wire                toplevel_execute_lane1_bypasser_integer_RS1_along_bypasses_1_checks_0_selfHit;
  wire                toplevel_execute_lane1_bypasser_integer_RS1_along_bypasses_1_checks_0_hit;
  wire                toplevel_execute_lane1_bypasser_integer_RS1_along_bypasses_1_checks_1_selfHit;
  wire                toplevel_execute_lane1_bypasser_integer_RS1_along_bypasses_1_checks_1_hit;
  wire       [1:0]    toplevel_execute_lane1_bypasser_integer_RS1_along_bypasses_1_hits;
  wire       [2:0]    _zz_toplevel_execute_ctrl3_integer_RS1_lane1_bypass;
  wire                toplevel_execute_lane1_bypasser_integer_RS2_port_valid;
  wire       [4:0]    toplevel_execute_lane1_bypasser_integer_RS2_port_address;
  wire       [31:0]   toplevel_execute_lane1_bypasser_integer_RS2_port_data;
  reg        [8:0]    toplevel_execute_lane1_bypasser_integer_RS2_bypassEnables;
  wire       [8:0]    _zz_toplevel_execute_lane1_bypasser_integer_RS2_bypassEnables_bools_0;
  wire                toplevel_execute_lane1_bypasser_integer_RS2_bypassEnables_bools_0;
  wire                toplevel_execute_lane1_bypasser_integer_RS2_bypassEnables_bools_1;
  wire                toplevel_execute_lane1_bypasser_integer_RS2_bypassEnables_bools_2;
  wire                toplevel_execute_lane1_bypasser_integer_RS2_bypassEnables_bools_3;
  wire                toplevel_execute_lane1_bypasser_integer_RS2_bypassEnables_bools_4;
  wire                toplevel_execute_lane1_bypasser_integer_RS2_bypassEnables_bools_5;
  wire                toplevel_execute_lane1_bypasser_integer_RS2_bypassEnables_bools_6;
  wire                toplevel_execute_lane1_bypasser_integer_RS2_bypassEnables_bools_7;
  wire                toplevel_execute_lane1_bypasser_integer_RS2_bypassEnables_bools_8;
  reg        [8:0]    _zz_toplevel_execute_lane1_bypasser_integer_RS2_sel;
  wire                toplevel_execute_lane1_bypasser_integer_RS2_bypassEnables_range_0_to_1;
  wire                toplevel_execute_lane1_bypasser_integer_RS2_bypassEnables_range_0_to_2;
  wire                toplevel_execute_lane1_bypasser_integer_RS2_bypassEnables_range_0_to_3;
  wire                toplevel_execute_lane1_bypasser_integer_RS2_bypassEnables_range_4_to_5;
  wire                toplevel_execute_lane1_bypasser_integer_RS2_bypassEnables_range_4_to_6;
  wire                toplevel_execute_lane1_bypasser_integer_RS2_bypassEnables_range_4_to_7;
  wire       [8:0]    toplevel_execute_lane1_bypasser_integer_RS2_sel;
  wire       [7:0]    _zz_toplevel_execute_ctrl1_down_integer_RS2_lane1;
  (* keep , syn_keep *) reg        [31:0]   _zz_toplevel_execute_ctrl1_down_integer_RS2_lane1_1 /* synthesis syn_keep = 1 */ ;
  wire                when_ExecuteLanePlugin_l190_3;
  wire                toplevel_execute_lane1_bypasser_integer_RS2_along_bypasses_0_checks_0_selfHit;
  wire                toplevel_execute_lane1_bypasser_integer_RS2_along_bypasses_0_checks_0_hit;
  wire                toplevel_execute_lane1_bypasser_integer_RS2_along_bypasses_0_checks_1_selfHit;
  wire                toplevel_execute_lane1_bypasser_integer_RS2_along_bypasses_0_checks_1_youngerHits_0;
  wire                toplevel_execute_lane1_bypasser_integer_RS2_along_bypasses_0_checks_1_youngerHits_1;
  wire                toplevel_execute_lane1_bypasser_integer_RS2_along_bypasses_0_checks_1_hit;
  wire                toplevel_execute_lane1_bypasser_integer_RS2_along_bypasses_0_checks_2_selfHit;
  wire                toplevel_execute_lane1_bypasser_integer_RS2_along_bypasses_0_checks_2_hit;
  wire                toplevel_execute_lane1_bypasser_integer_RS2_along_bypasses_0_checks_3_selfHit;
  wire                toplevel_execute_lane1_bypasser_integer_RS2_along_bypasses_0_checks_3_youngerHits_0;
  wire                toplevel_execute_lane1_bypasser_integer_RS2_along_bypasses_0_checks_3_youngerHits_1;
  wire                toplevel_execute_lane1_bypasser_integer_RS2_along_bypasses_0_checks_3_hit;
  wire       [3:0]    toplevel_execute_lane1_bypasser_integer_RS2_along_bypasses_0_hits;
  wire       [4:0]    _zz_toplevel_execute_ctrl2_integer_RS2_lane1_bypass;
  wire                toplevel_execute_lane1_bypasser_integer_RS2_along_bypasses_1_checks_0_selfHit;
  wire                toplevel_execute_lane1_bypasser_integer_RS2_along_bypasses_1_checks_0_hit;
  wire                toplevel_execute_lane1_bypasser_integer_RS2_along_bypasses_1_checks_1_selfHit;
  wire                toplevel_execute_lane1_bypasser_integer_RS2_along_bypasses_1_checks_1_hit;
  wire       [1:0]    toplevel_execute_lane1_bypasser_integer_RS2_along_bypasses_1_hits;
  wire       [2:0]    _zz_toplevel_execute_ctrl3_integer_RS2_lane1_bypass;
  wire                execute_lane1_logic_completions_onCtrl_0_port_valid;
  wire       [15:0]   execute_lane1_logic_completions_onCtrl_0_port_payload_uopId;
  wire                execute_lane1_logic_completions_onCtrl_0_port_payload_trap;
  wire                execute_lane1_logic_completions_onCtrl_0_port_payload_commit;
  wire                execute_lane1_logic_completions_onCtrl_1_port_valid;
  wire       [15:0]   execute_lane1_logic_completions_onCtrl_1_port_payload_uopId;
  wire                execute_lane1_logic_completions_onCtrl_1_port_payload_trap;
  wire                execute_lane1_logic_completions_onCtrl_1_port_payload_commit;
  wire                execute_lane1_logic_completions_onCtrl_2_port_valid;
  wire       [15:0]   execute_lane1_logic_completions_onCtrl_2_port_payload_uopId;
  wire                execute_lane1_logic_completions_onCtrl_2_port_payload_trap;
  wire                execute_lane1_logic_completions_onCtrl_2_port_payload_commit;
  wire       [32:0]   execute_lane1_logic_decoding_decodingBits;
  wire                _zz_toplevel_execute_ctrl1_down_execute_lane1_logic_completions_onCtrl_0_ENABLE_lane1;
  wire                _zz_toplevel_execute_ctrl1_down_execute_lane1_logic_completions_onCtrl_0_ENABLE_lane1_1;
  wire                _zz_toplevel_execute_ctrl1_down_execute_lane1_logic_completions_onCtrl_0_ENABLE_lane1_2;
  wire                _zz_toplevel_execute_ctrl1_down_execute_lane1_logic_completions_onCtrl_1_ENABLE_lane1;
  wire                _zz_toplevel_execute_ctrl1_down_late1_BranchPlugin_SEL_lane1;
  wire                _zz_toplevel_execute_ctrl1_down_late1_SrcPlugin_logic_SRC2_CTRL_lane1;
  wire                _zz_toplevel_execute_ctrl1_down_execute_lane1_logic_completions_onCtrl_1_ENABLE_lane1_1;
  wire                _zz_toplevel_execute_ctrl1_down_execute_lane1_logic_completions_onCtrl_2_ENABLE_lane1;
  wire                _zz_toplevel_execute_ctrl1_down_late1_IntAluPlugin_ALU_ADD_SUB_lane1;
  wire                _zz_toplevel_execute_ctrl1_down_late1_IntAluPlugin_ALU_SLTX_lane1;
  wire                _zz_toplevel_execute_ctrl1_down_late1_IntAluPlugin_ALU_BITWISE_CTRL_lane1;
  wire                _zz_toplevel_execute_ctrl1_down_BarrelShifterPlugin_LEFT_lane1;
  wire                _zz_toplevel_execute_ctrl1_down_late1_IntAluPlugin_ALU_BITWISE_CTRL_lane1_1;
  wire       [1:0]    _zz_toplevel_execute_ctrl1_down_early1_IntAluPlugin_ALU_BITWISE_CTRL_lane1;
  wire       [1:0]    _zz_toplevel_execute_ctrl1_down_early1_IntAluPlugin_ALU_BITWISE_CTRL_lane1_1;
  wire       [1:0]    _zz_toplevel_execute_ctrl1_down_early1_IntAluPlugin_ALU_BITWISE_CTRL_lane1_2;
  wire                _zz_toplevel_execute_ctrl1_down_SrcStageables_REVERT_lane1;
  wire                _zz_toplevel_execute_ctrl1_down_late1_SrcPlugin_logic_SRC2_CTRL_lane1_1;
  wire       [1:0]    _zz_toplevel_execute_ctrl1_down_BranchPlugin_BRANCH_CTRL_lane1;
  wire       [1:0]    _zz_toplevel_execute_ctrl1_down_BranchPlugin_BRANCH_CTRL_lane1_1;
  wire       [1:0]    _zz_toplevel_execute_ctrl1_down_BranchPlugin_BRANCH_CTRL_lane1_2;
  wire       [1:0]    _zz_toplevel_execute_ctrl1_down_late1_IntAluPlugin_ALU_BITWISE_CTRL_lane1_2;
  wire       [1:0]    _zz_toplevel_execute_ctrl1_down_late1_IntAluPlugin_ALU_BITWISE_CTRL_lane1_3;
  wire       [1:0]    _zz_toplevel_execute_ctrl1_down_late1_IntAluPlugin_ALU_BITWISE_CTRL_lane1_4;
  wire                when_ExecuteLanePlugin_l300_5;
  wire                when_ExecuteLanePlugin_l300_6;
  wire                when_ExecuteLanePlugin_l300_7;
  wire                when_ExecuteLanePlugin_l300_8;
  wire                when_ExecuteLanePlugin_l300_9;
  wire                integer_RegFilePlugin_logic_writeMerges_0_bus_valid;
  wire       [4:0]    integer_RegFilePlugin_logic_writeMerges_0_bus_address;
  wire       [31:0]   integer_RegFilePlugin_logic_writeMerges_0_bus_data;
  wire       [15:0]   integer_RegFilePlugin_logic_writeMerges_0_bus_uopId;
  wire                integer_RegFilePlugin_logic_writeMerges_1_bus_valid;
  wire       [4:0]    integer_RegFilePlugin_logic_writeMerges_1_bus_address;
  wire       [31:0]   integer_RegFilePlugin_logic_writeMerges_1_bus_data;
  wire       [15:0]   integer_RegFilePlugin_logic_writeMerges_1_bus_uopId;
  reg        [5:0]    integer_RegFilePlugin_logic_initalizer_counter;
  wire                integer_RegFilePlugin_logic_initalizer_done;
  wire                when_RegFilePlugin_l127;
  wire                integer_write_0_valid /* verilator public */ ;
  wire       [4:0]    integer_write_0_address /* verilator public */ ;
  wire       [31:0]   integer_write_0_data /* verilator public */ ;
  wire       [15:0]   integer_write_0_uopId /* verilator public */ ;
  wire                integer_write_1_valid /* verilator public */ ;
  wire       [4:0]    integer_write_1_address /* verilator public */ ;
  wire       [31:0]   integer_write_1_data /* verilator public */ ;
  wire       [15:0]   integer_write_1_uopId /* verilator public */ ;
  wire       [31:0]   FetchL1Plugin_pmaBuilder_addressBits;
  wire                _zz_FetchL1Plugin_logic_ctrl_pmaPort_rsp_io;
  wire                FetchL1Plugin_pmaBuilder_onTransfers_0_addressHit;
  wire                FetchL1Plugin_pmaBuilder_onTransfers_0_argsHit;
  wire                FetchL1Plugin_pmaBuilder_onTransfers_0_hit;
  wire       [31:0]   LsuPlugin_pmaBuilder_l1_addressBits;
  wire       [0:0]    LsuPlugin_pmaBuilder_l1_argsBits;
  wire                _zz_LsuPlugin_logic_onPma_cached_rsp_io;
  wire                LsuPlugin_pmaBuilder_l1_onTransfers_0_addressHit;
  wire                LsuPlugin_pmaBuilder_l1_onTransfers_0_argsHit;
  wire                LsuPlugin_pmaBuilder_l1_onTransfers_0_hit;
  wire       [31:0]   LsuPlugin_pmaBuilder_io_addressBits;
  wire       [2:0]    LsuPlugin_pmaBuilder_io_argsBits;
  wire                LsuPlugin_pmaBuilder_io_onTransfers_0_addressHit;
  wire                LsuPlugin_pmaBuilder_io_onTransfers_0_argsHit;
  wire                LsuPlugin_pmaBuilder_io_onTransfers_0_hit;
  wire                _zz_LsuPlugin_logic_onPma_io_rsp_io;
  wire                _zz_LsuPlugin_logic_onPma_io_rsp_io_1;
  wire                LsuPlugin_pmaBuilder_io_onTransfers_1_addressHit;
  wire                LsuPlugin_pmaBuilder_io_onTransfers_1_argsHit;
  wire                LsuPlugin_pmaBuilder_io_onTransfers_1_hit;
  wire                WhiteboxerPlugin_logic_completions_ports_5_valid;
  wire       [15:0]   WhiteboxerPlugin_logic_completions_ports_5_payload_uopId;
  wire                WhiteboxerPlugin_logic_completions_ports_5_payload_trap;
  wire                WhiteboxerPlugin_logic_completions_ports_5_payload_commit;
  wire                WhiteboxerPlugin_logic_completions_ports_6_valid;
  wire       [15:0]   WhiteboxerPlugin_logic_completions_ports_6_payload_uopId;
  wire                WhiteboxerPlugin_logic_completions_ports_6_payload_trap;
  wire                WhiteboxerPlugin_logic_completions_ports_6_payload_commit;
  wire                WhiteboxerPlugin_logic_completions_ports_7_valid;
  wire       [15:0]   WhiteboxerPlugin_logic_completions_ports_7_payload_uopId;
  wire                WhiteboxerPlugin_logic_completions_ports_7_payload_trap;
  wire                WhiteboxerPlugin_logic_completions_ports_7_payload_commit;
  wire                WhiteboxerPlugin_logic_commits_ports_0_oh_0;
  wire                WhiteboxerPlugin_logic_commits_ports_0_oh_1;
  wire                WhiteboxerPlugin_logic_commits_ports_0_valid;
  wire       [31:0]   WhiteboxerPlugin_logic_commits_ports_0_pc;
  wire       [31:0]   WhiteboxerPlugin_logic_commits_ports_0_uop;
  wire                WhiteboxerPlugin_logic_commits_ports_1_oh_0;
  wire                WhiteboxerPlugin_logic_commits_ports_1_oh_1;
  wire                WhiteboxerPlugin_logic_commits_ports_1_valid;
  wire       [31:0]   WhiteboxerPlugin_logic_commits_ports_1_pc;
  wire       [31:0]   WhiteboxerPlugin_logic_commits_ports_1_uop;
  wire                WhiteboxerPlugin_logic_reschedules_flushes_0_valid;
  wire                WhiteboxerPlugin_logic_reschedules_flushes_0_payload_self;
  wire                WhiteboxerPlugin_logic_reschedules_flushes_1_valid;
  wire       [15:0]   WhiteboxerPlugin_logic_reschedules_flushes_1_payload_uopId;
  wire       [0:0]    WhiteboxerPlugin_logic_reschedules_flushes_1_payload_laneAge;
  wire                WhiteboxerPlugin_logic_reschedules_flushes_1_payload_self;
  wire                WhiteboxerPlugin_logic_reschedules_flushes_2_valid;
  wire       [15:0]   WhiteboxerPlugin_logic_reschedules_flushes_2_payload_uopId;
  wire       [0:0]    WhiteboxerPlugin_logic_reschedules_flushes_2_payload_laneAge;
  wire                WhiteboxerPlugin_logic_reschedules_flushes_2_payload_self;
  wire                WhiteboxerPlugin_logic_reschedules_flushes_3_valid;
  wire       [15:0]   WhiteboxerPlugin_logic_reschedules_flushes_3_payload_uopId;
  wire       [0:0]    WhiteboxerPlugin_logic_reschedules_flushes_3_payload_laneAge;
  wire                WhiteboxerPlugin_logic_reschedules_flushes_3_payload_self;
  wire                WhiteboxerPlugin_logic_reschedules_flushes_4_valid;
  wire       [15:0]   WhiteboxerPlugin_logic_reschedules_flushes_4_payload_uopId;
  wire       [0:0]    WhiteboxerPlugin_logic_reschedules_flushes_4_payload_laneAge;
  wire                WhiteboxerPlugin_logic_reschedules_flushes_4_payload_self;
  wire                WhiteboxerPlugin_logic_reschedules_flushes_5_valid;
  wire       [15:0]   WhiteboxerPlugin_logic_reschedules_flushes_5_payload_uopId;
  wire       [0:0]    WhiteboxerPlugin_logic_reschedules_flushes_5_payload_laneAge;
  wire                WhiteboxerPlugin_logic_reschedules_flushes_5_payload_self;
  wire                WhiteboxerPlugin_logic_reschedules_flushes_6_valid;
  wire       [15:0]   WhiteboxerPlugin_logic_reschedules_flushes_6_payload_uopId;
  wire       [0:0]    WhiteboxerPlugin_logic_reschedules_flushes_6_payload_laneAge;
  wire                WhiteboxerPlugin_logic_reschedules_flushes_6_payload_self;
  wire                WhiteboxerPlugin_logic_reschedules_flushes_7_valid;
  wire       [15:0]   WhiteboxerPlugin_logic_reschedules_flushes_7_payload_uopId;
  wire       [0:0]    WhiteboxerPlugin_logic_reschedules_flushes_7_payload_laneAge;
  wire                WhiteboxerPlugin_logic_reschedules_flushes_7_payload_self;
  wire                WhiteboxerPlugin_logic_reschedules_flushes_8_valid;
  wire       [15:0]   WhiteboxerPlugin_logic_reschedules_flushes_8_payload_uopId;
  wire       [0:0]    WhiteboxerPlugin_logic_reschedules_flushes_8_payload_laneAge;
  wire                WhiteboxerPlugin_logic_reschedules_flushes_8_payload_self;
  wire                WhiteboxerPlugin_logic_reschedules_flushes_9_valid;
  wire       [15:0]   WhiteboxerPlugin_logic_reschedules_flushes_9_payload_uopId;
  wire       [0:0]    WhiteboxerPlugin_logic_reschedules_flushes_9_payload_laneAge;
  wire                WhiteboxerPlugin_logic_reschedules_flushes_9_payload_self;
  wire                WhiteboxerPlugin_logic_prediction_learns_0_valid;
  wire       [31:0]   WhiteboxerPlugin_logic_prediction_learns_0_payload_pcOnLastSlice;
  wire       [31:0]   WhiteboxerPlugin_logic_prediction_learns_0_payload_pcTarget;
  wire                WhiteboxerPlugin_logic_prediction_learns_0_payload_taken;
  wire                WhiteboxerPlugin_logic_prediction_learns_0_payload_isBranch;
  wire                WhiteboxerPlugin_logic_prediction_learns_0_payload_isPush;
  wire                WhiteboxerPlugin_logic_prediction_learns_0_payload_isPop;
  wire                WhiteboxerPlugin_logic_prediction_learns_0_payload_wasWrong;
  wire                WhiteboxerPlugin_logic_prediction_learns_0_payload_badPredictedTarget;
  wire       [11:0]   WhiteboxerPlugin_logic_prediction_learns_0_payload_history;
  wire       [15:0]   WhiteboxerPlugin_logic_prediction_learns_0_payload_uopId;
  wire       [1:0]    WhiteboxerPlugin_logic_prediction_learns_0_payload_ctx_GSharePlugin_GSHARE_COUNTER_0;
  wire       [1:0]    WhiteboxerPlugin_logic_prediction_learns_0_payload_ctx_GSharePlugin_GSHARE_COUNTER_1;
  wire       [1:0]    WhiteboxerPlugin_logic_prediction_learns_0_payload_ctx_GSharePlugin_GSHARE_COUNTER_2;
  wire       [1:0]    WhiteboxerPlugin_logic_prediction_learns_0_payload_ctx_GSharePlugin_GSHARE_COUNTER_3;
  wire                WhiteboxerPlugin_logic_prediction_learns_1_valid;
  wire       [31:0]   WhiteboxerPlugin_logic_prediction_learns_1_payload_pcOnLastSlice;
  wire       [31:0]   WhiteboxerPlugin_logic_prediction_learns_1_payload_pcTarget;
  wire                WhiteboxerPlugin_logic_prediction_learns_1_payload_taken;
  wire                WhiteboxerPlugin_logic_prediction_learns_1_payload_isBranch;
  wire                WhiteboxerPlugin_logic_prediction_learns_1_payload_isPush;
  wire                WhiteboxerPlugin_logic_prediction_learns_1_payload_isPop;
  wire                WhiteboxerPlugin_logic_prediction_learns_1_payload_wasWrong;
  wire                WhiteboxerPlugin_logic_prediction_learns_1_payload_badPredictedTarget;
  wire       [11:0]   WhiteboxerPlugin_logic_prediction_learns_1_payload_history;
  wire       [15:0]   WhiteboxerPlugin_logic_prediction_learns_1_payload_uopId;
  wire       [1:0]    WhiteboxerPlugin_logic_prediction_learns_1_payload_ctx_GSharePlugin_GSHARE_COUNTER_0;
  wire       [1:0]    WhiteboxerPlugin_logic_prediction_learns_1_payload_ctx_GSharePlugin_GSHARE_COUNTER_1;
  wire       [1:0]    WhiteboxerPlugin_logic_prediction_learns_1_payload_ctx_GSharePlugin_GSHARE_COUNTER_2;
  wire       [1:0]    WhiteboxerPlugin_logic_prediction_learns_1_payload_ctx_GSharePlugin_GSHARE_COUNTER_3;
  wire                WhiteboxerPlugin_logic_loadExecute_fire;
  wire       [15:0]   WhiteboxerPlugin_logic_loadExecute_uopId;
  wire       [1:0]    WhiteboxerPlugin_logic_loadExecute_size;
  wire       [31:0]   WhiteboxerPlugin_logic_loadExecute_address;
  wire       [31:0]   WhiteboxerPlugin_logic_loadExecute_data;
  wire                WhiteboxerPlugin_logic_storeCommit_fire;
  wire       [15:0]   WhiteboxerPlugin_logic_storeCommit_uopId;
  wire       [11:0]   WhiteboxerPlugin_logic_storeCommit_storeId;
  wire       [1:0]    WhiteboxerPlugin_logic_storeCommit_size;
  wire       [31:0]   WhiteboxerPlugin_logic_storeCommit_address;
  wire       [31:0]   WhiteboxerPlugin_logic_storeCommit_data;
  wire                WhiteboxerPlugin_logic_storeCommit_amo;
  wire                WhiteboxerPlugin_logic_storeConditional_fire;
  wire       [15:0]   WhiteboxerPlugin_logic_storeConditional_uopId;
  wire                WhiteboxerPlugin_logic_storeConditional_miss;
  wire                WhiteboxerPlugin_logic_storeBroadcast_fire;
  wire       [11:0]   WhiteboxerPlugin_logic_storeBroadcast_storeId;
  wire       [0:0]    WhiteboxerPlugin_logic_wfi;
  wire                WhiteboxerPlugin_logic_perf_executeFreezed;
  wire                WhiteboxerPlugin_logic_perf_dispatchHazards;
  wire       [1:0]    WhiteboxerPlugin_logic_perf_candidatesCount;
  wire       [1:0]    WhiteboxerPlugin_logic_perf_dispatchFeedCount;
  reg                 _zz_WhiteboxerPlugin_logic_perf_executeFreezedCounter;
  reg        [59:0]   _zz_WhiteboxerPlugin_logic_perf_executeFreezedCounter_1;
  reg        [59:0]   _zz_WhiteboxerPlugin_logic_perf_executeFreezedCounter_2;
  wire       [59:0]   WhiteboxerPlugin_logic_perf_executeFreezedCounter;
  reg                 _zz_WhiteboxerPlugin_logic_perf_dispatchHazardsCounter;
  reg        [59:0]   _zz_WhiteboxerPlugin_logic_perf_dispatchHazardsCounter_1;
  reg        [59:0]   _zz_WhiteboxerPlugin_logic_perf_dispatchHazardsCounter_2;
  wire       [59:0]   WhiteboxerPlugin_logic_perf_dispatchHazardsCounter;
  wire                when_Utils_l585;
  reg                 _zz_WhiteboxerPlugin_logic_perf_candidatesCountCounters_0;
  reg        [59:0]   _zz_WhiteboxerPlugin_logic_perf_candidatesCountCounters_0_1;
  reg        [59:0]   _zz_WhiteboxerPlugin_logic_perf_candidatesCountCounters_0_2;
  wire       [59:0]   WhiteboxerPlugin_logic_perf_candidatesCountCounters_0;
  wire                when_Utils_l585_1;
  reg                 _zz_WhiteboxerPlugin_logic_perf_candidatesCountCounters_1;
  reg        [59:0]   _zz_WhiteboxerPlugin_logic_perf_candidatesCountCounters_1_1;
  reg        [59:0]   _zz_WhiteboxerPlugin_logic_perf_candidatesCountCounters_1_2;
  wire       [59:0]   WhiteboxerPlugin_logic_perf_candidatesCountCounters_1;
  wire                when_Utils_l585_2;
  reg                 _zz_WhiteboxerPlugin_logic_perf_candidatesCountCounters_2;
  reg        [59:0]   _zz_WhiteboxerPlugin_logic_perf_candidatesCountCounters_2_1;
  reg        [59:0]   _zz_WhiteboxerPlugin_logic_perf_candidatesCountCounters_2_2;
  wire       [59:0]   WhiteboxerPlugin_logic_perf_candidatesCountCounters_2;
  wire                when_Utils_l585_3;
  reg                 _zz_WhiteboxerPlugin_logic_perf_candidatesCountCounters_3;
  reg        [59:0]   _zz_WhiteboxerPlugin_logic_perf_candidatesCountCounters_3_1;
  reg        [59:0]   _zz_WhiteboxerPlugin_logic_perf_candidatesCountCounters_3_2;
  wire       [59:0]   WhiteboxerPlugin_logic_perf_candidatesCountCounters_3;
  wire                when_Utils_l585_4;
  reg                 _zz_WhiteboxerPlugin_logic_perf_dispatchFeedCounters_0;
  reg        [59:0]   _zz_WhiteboxerPlugin_logic_perf_dispatchFeedCounters_0_1;
  reg        [59:0]   _zz_WhiteboxerPlugin_logic_perf_dispatchFeedCounters_0_2;
  wire       [59:0]   WhiteboxerPlugin_logic_perf_dispatchFeedCounters_0;
  wire                when_Utils_l585_5;
  reg                 _zz_WhiteboxerPlugin_logic_perf_dispatchFeedCounters_1;
  reg        [59:0]   _zz_WhiteboxerPlugin_logic_perf_dispatchFeedCounters_1_1;
  reg        [59:0]   _zz_WhiteboxerPlugin_logic_perf_dispatchFeedCounters_1_2;
  wire       [59:0]   WhiteboxerPlugin_logic_perf_dispatchFeedCounters_1;
  wire                when_Utils_l585_6;
  reg                 _zz_WhiteboxerPlugin_logic_perf_dispatchFeedCounters_2;
  reg        [59:0]   _zz_WhiteboxerPlugin_logic_perf_dispatchFeedCounters_2_1;
  reg        [59:0]   _zz_WhiteboxerPlugin_logic_perf_dispatchFeedCounters_2_2;
  wire       [59:0]   WhiteboxerPlugin_logic_perf_dispatchFeedCounters_2;
  wire                WhiteboxerPlugin_logic_trap_ports_0_valid;
  wire                WhiteboxerPlugin_logic_trap_ports_0_interrupt;
  wire       [3:0]    WhiteboxerPlugin_logic_trap_ports_0_cause;
  wire                fetch_logic_ctrls_2_up_forgetOne;
  wire                fetch_logic_ctrls_1_up_forgetOne;
  wire                when_CtrlLink_l150;
  wire                when_CtrlLink_l157;
  wire                when_StageLink_l67;
  wire                when_DecodePipelinePlugin_l68;
  wire                when_DecodePipelinePlugin_l68_1;
  reg        [1:0]    LsuPlugin_logic_flusher_stateReg;
  reg        [1:0]    LsuPlugin_logic_flusher_stateNext;
  wire                when_LsuPlugin_l297;
  wire                when_LsuPlugin_l305;
  reg        [3:0]    TrapPlugin_logic_harts_0_trap_fsm_stateReg;
  reg        [3:0]    TrapPlugin_logic_harts_0_trap_fsm_stateNext;
  wire                when_TrapPlugin_l393;
  reg        [2:0]    _zz_TrapPlugin_logic_harts_0_crsPorts_write_address;
  reg        [2:0]    _zz_TrapPlugin_logic_harts_0_crsPorts_write_address_1;
  reg        [2:0]    _zz_TrapPlugin_logic_harts_0_crsPorts_read_address;
  reg        [2:0]    _zz_TrapPlugin_logic_harts_0_crsPorts_read_address_1;
  wire                when_TrapPlugin_l637;
  wire       [1:0]    switch_TrapPlugin_l638;
  wire                when_TrapPlugin_l492;
  wire       [2:0]    switch_TrapPlugin_l494;
  wire                when_TrapPlugin_l348;
  reg        [2:0]    MmuPlugin_logic_refill_stateReg;
  reg        [2:0]    MmuPlugin_logic_refill_stateNext;
  wire                when_MmuPlugin_l454;
  wire                when_MmuPlugin_l454_1;
  wire                when_MmuPlugin_l463;
  wire                when_MmuPlugin_l439;
  wire                _zz_54;
  wire                when_MmuPlugin_l439_1;
  wire                when_MmuPlugin_l471;
  wire                when_MmuPlugin_l439_2;
  wire                when_MmuPlugin_l439_3;
  reg        [1:0]    CsrAccessPlugin_logic_fsm_stateReg;
  reg        [1:0]    CsrAccessPlugin_logic_fsm_stateNext;
  wire                when_CsrAccessPlugin_l308;
  wire                when_CsrAccessPlugin_l338;
  wire                when_CsrAccessPlugin_l224;
  `ifndef SYNTHESIS
  reg [39:0] toplevel_execute_ctrl3_down_late1_IntAluPlugin_ALU_BITWISE_CTRL_lane1_string;
  reg [39:0] toplevel_execute_ctrl3_down_late0_IntAluPlugin_ALU_BITWISE_CTRL_lane0_string;
  reg [39:0] toplevel_execute_ctrl4_up_late1_IntAluPlugin_ALU_BITWISE_CTRL_lane1_string;
  reg [31:0] toplevel_execute_ctrl4_up_BranchPlugin_BRANCH_CTRL_lane1_string;
  reg [39:0] toplevel_execute_ctrl4_up_late0_IntAluPlugin_ALU_BITWISE_CTRL_lane0_string;
  reg [31:0] toplevel_execute_ctrl4_up_BranchPlugin_BRANCH_CTRL_lane0_string;
  reg [39:0] toplevel_execute_ctrl2_down_late1_IntAluPlugin_ALU_BITWISE_CTRL_lane1_string;
  reg [39:0] toplevel_execute_ctrl2_down_late0_IntAluPlugin_ALU_BITWISE_CTRL_lane0_string;
  reg [39:0] toplevel_execute_ctrl3_up_late1_IntAluPlugin_ALU_BITWISE_CTRL_lane1_string;
  reg [31:0] toplevel_execute_ctrl3_up_BranchPlugin_BRANCH_CTRL_lane1_string;
  reg [39:0] toplevel_execute_ctrl3_up_late0_IntAluPlugin_ALU_BITWISE_CTRL_lane0_string;
  reg [31:0] toplevel_execute_ctrl3_up_BranchPlugin_BRANCH_CTRL_lane0_string;
  reg [39:0] toplevel_execute_ctrl2_up_late1_IntAluPlugin_ALU_BITWISE_CTRL_lane1_string;
  reg [31:0] toplevel_execute_ctrl2_up_BranchPlugin_BRANCH_CTRL_lane1_string;
  reg [39:0] toplevel_execute_ctrl2_up_early1_IntAluPlugin_ALU_BITWISE_CTRL_lane1_string;
  reg [39:0] toplevel_execute_ctrl2_up_late0_IntAluPlugin_ALU_BITWISE_CTRL_lane0_string;
  reg [79:0] toplevel_execute_ctrl2_up_early0_EnvPlugin_OP_lane0_string;
  reg [31:0] toplevel_execute_ctrl2_up_BranchPlugin_BRANCH_CTRL_lane0_string;
  reg [39:0] toplevel_execute_ctrl2_up_early0_IntAluPlugin_ALU_BITWISE_CTRL_lane0_string;
  reg [39:0] toplevel_execute_ctrl1_down_late1_IntAluPlugin_ALU_BITWISE_CTRL_lane1_string;
  reg [31:0] toplevel_execute_ctrl1_down_BranchPlugin_BRANCH_CTRL_lane1_string;
  reg [39:0] toplevel_execute_ctrl1_down_early1_IntAluPlugin_ALU_BITWISE_CTRL_lane1_string;
  reg [39:0] toplevel_execute_ctrl1_down_late0_IntAluPlugin_ALU_BITWISE_CTRL_lane0_string;
  reg [79:0] toplevel_execute_ctrl1_down_early0_EnvPlugin_OP_lane0_string;
  reg [31:0] toplevel_execute_ctrl1_down_BranchPlugin_BRANCH_CTRL_lane0_string;
  reg [39:0] toplevel_execute_ctrl1_down_early0_IntAluPlugin_ALU_BITWISE_CTRL_lane0_string;
  reg [31:0] toplevel_execute_ctrl4_down_BranchPlugin_BRANCH_CTRL_lane1_string;
  reg [31:0] toplevel_execute_ctrl4_down_BranchPlugin_BRANCH_CTRL_lane0_string;
  reg [31:0] toplevel_execute_ctrl3_down_BranchPlugin_BRANCH_CTRL_lane1_string;
  reg [79:0] toplevel_execute_ctrl2_down_early0_EnvPlugin_OP_lane0_string;
  reg [31:0] toplevel_execute_ctrl3_down_BranchPlugin_BRANCH_CTRL_lane0_string;
  reg [31:0] toplevel_execute_ctrl2_down_BranchPlugin_BRANCH_CTRL_lane1_string;
  reg [31:0] toplevel_execute_ctrl2_down_BranchPlugin_BRANCH_CTRL_lane0_string;
  reg [39:0] toplevel_execute_ctrl4_down_late1_IntAluPlugin_ALU_BITWISE_CTRL_lane1_string;
  reg [39:0] toplevel_execute_ctrl2_down_early1_IntAluPlugin_ALU_BITWISE_CTRL_lane1_string;
  reg [39:0] toplevel_execute_ctrl4_down_late0_IntAluPlugin_ALU_BITWISE_CTRL_lane0_string;
  reg [39:0] toplevel_execute_ctrl2_down_early0_IntAluPlugin_ALU_BITWISE_CTRL_lane0_string;
  reg [127:0] FetchL1TileLinkPlugin_logic_down_a_payload_opcode_string;
  reg [119:0] FetchL1TileLinkPlugin_logic_down_d_payload_opcode_string;
  reg [95:0] LsuPlugin_logic_onAddress0_ls_port_payload_op_string;
  reg [95:0] LsuPlugin_logic_onAddress0_access_port_payload_op_string;
  reg [95:0] LsuPlugin_logic_onAddress0_flush_port_payload_op_string;
  reg [127:0] LsuL1TileLinkPlugin_logic_down_a_payload_opcode_string;
  reg [119:0] LsuL1TileLinkPlugin_logic_down_d_payload_opcode_string;
  reg [127:0] LsuTileLinkPlugin_logic_bridge_down_a_payload_opcode_string;
  reg [119:0] LsuTileLinkPlugin_logic_bridge_down_d_payload_opcode_string;
  reg [127:0] _zz_LsuTileLinkPlugin_logic_bridge_down_a_payload_opcode_string;
  reg [39:0] _zz_toplevel_execute_ctrl1_down_early0_IntAluPlugin_ALU_BITWISE_CTRL_lane0_string;
  reg [39:0] _zz_toplevel_execute_ctrl1_down_early0_IntAluPlugin_ALU_BITWISE_CTRL_lane0_1_string;
  reg [39:0] _zz_toplevel_execute_ctrl1_down_early0_IntAluPlugin_ALU_BITWISE_CTRL_lane0_2_string;
  reg [31:0] _zz_toplevel_execute_ctrl1_down_BranchPlugin_BRANCH_CTRL_lane0_string;
  reg [31:0] _zz_toplevel_execute_ctrl1_down_BranchPlugin_BRANCH_CTRL_lane0_1_string;
  reg [31:0] _zz_toplevel_execute_ctrl1_down_BranchPlugin_BRANCH_CTRL_lane0_2_string;
  reg [79:0] _zz_toplevel_execute_ctrl1_down_early0_EnvPlugin_OP_lane0_1_string;
  reg [79:0] _zz_toplevel_execute_ctrl1_down_early0_EnvPlugin_OP_lane0_2_string;
  reg [79:0] _zz_toplevel_execute_ctrl1_down_early0_EnvPlugin_OP_lane0_3_string;
  reg [39:0] _zz_toplevel_execute_ctrl1_down_late0_IntAluPlugin_ALU_BITWISE_CTRL_lane0_1_string;
  reg [39:0] _zz_toplevel_execute_ctrl1_down_late0_IntAluPlugin_ALU_BITWISE_CTRL_lane0_2_string;
  reg [39:0] _zz_toplevel_execute_ctrl1_down_late0_IntAluPlugin_ALU_BITWISE_CTRL_lane0_3_string;
  reg [39:0] _zz_toplevel_execute_ctrl1_down_early1_IntAluPlugin_ALU_BITWISE_CTRL_lane1_string;
  reg [39:0] _zz_toplevel_execute_ctrl1_down_early1_IntAluPlugin_ALU_BITWISE_CTRL_lane1_1_string;
  reg [39:0] _zz_toplevel_execute_ctrl1_down_early1_IntAluPlugin_ALU_BITWISE_CTRL_lane1_2_string;
  reg [31:0] _zz_toplevel_execute_ctrl1_down_BranchPlugin_BRANCH_CTRL_lane1_string;
  reg [31:0] _zz_toplevel_execute_ctrl1_down_BranchPlugin_BRANCH_CTRL_lane1_1_string;
  reg [31:0] _zz_toplevel_execute_ctrl1_down_BranchPlugin_BRANCH_CTRL_lane1_2_string;
  reg [39:0] _zz_toplevel_execute_ctrl1_down_late1_IntAluPlugin_ALU_BITWISE_CTRL_lane1_2_string;
  reg [39:0] _zz_toplevel_execute_ctrl1_down_late1_IntAluPlugin_ALU_BITWISE_CTRL_lane1_3_string;
  reg [39:0] _zz_toplevel_execute_ctrl1_down_late1_IntAluPlugin_ALU_BITWISE_CTRL_lane1_4_string;
  reg [79:0] LsuPlugin_logic_flusher_stateReg_string;
  reg [79:0] LsuPlugin_logic_flusher_stateNext_string;
  reg [87:0] TrapPlugin_logic_harts_0_trap_fsm_stateReg_string;
  reg [87:0] TrapPlugin_logic_harts_0_trap_fsm_stateNext_string;
  reg [39:0] MmuPlugin_logic_refill_stateReg_string;
  reg [39:0] MmuPlugin_logic_refill_stateNext_string;
  reg [79:0] CsrAccessPlugin_logic_fsm_stateReg_string;
  reg [79:0] CsrAccessPlugin_logic_fsm_stateNext_string;
  `endif

  (* ram_style = "distributed" *) reg [30:0] BtbPlugin_logic_ras_mem_stack [0:3];
  reg [63:0] FetchL1Plugin_logic_banks_0_mem [0:511];
  reg [63:0] FetchL1Plugin_logic_banks_1_mem [0:511];
  reg [21:0] FetchL1Plugin_logic_ways_0_mem [0:63];
  reg [21:0] FetchL1Plugin_logic_ways_1_mem [0:63];
  reg [0:0] FetchL1Plugin_logic_plru_mem [0:63];
  reg [7:0] GSharePlugin_logic_mem_counter [0:4095];
  (* ram_style = "block" *) reg [50:0] BtbPlugin_logic_mem_symbol0 [0:255];
  (* ram_style = "block" *) reg [50:0] BtbPlugin_logic_mem_symbol1 [0:255];
  reg [50:0] _zz_BtbPlugin_logic_memsymbol_read;
  reg [50:0] _zz_BtbPlugin_logic_memsymbol_read_1;
  reg [7:0] LsuL1Plugin_logic_banks_0_mem_symbol0 [0:511];
  reg [7:0] LsuL1Plugin_logic_banks_0_mem_symbol1 [0:511];
  reg [7:0] LsuL1Plugin_logic_banks_0_mem_symbol2 [0:511];
  reg [7:0] LsuL1Plugin_logic_banks_0_mem_symbol3 [0:511];
  reg [7:0] LsuL1Plugin_logic_banks_0_mem_symbol4 [0:511];
  reg [7:0] LsuL1Plugin_logic_banks_0_mem_symbol5 [0:511];
  reg [7:0] LsuL1Plugin_logic_banks_0_mem_symbol6 [0:511];
  reg [7:0] LsuL1Plugin_logic_banks_0_mem_symbol7 [0:511];
  reg [7:0] _zz_LsuL1Plugin_logic_banks_0_memsymbol_read;
  reg [7:0] _zz_LsuL1Plugin_logic_banks_0_memsymbol_read_1;
  reg [7:0] _zz_LsuL1Plugin_logic_banks_0_memsymbol_read_2;
  reg [7:0] _zz_LsuL1Plugin_logic_banks_0_memsymbol_read_3;
  reg [7:0] _zz_LsuL1Plugin_logic_banks_0_memsymbol_read_4;
  reg [7:0] _zz_LsuL1Plugin_logic_banks_0_memsymbol_read_5;
  reg [7:0] _zz_LsuL1Plugin_logic_banks_0_memsymbol_read_6;
  reg [7:0] _zz_LsuL1Plugin_logic_banks_0_memsymbol_read_7;
  reg [7:0] LsuL1Plugin_logic_banks_1_mem_symbol0 [0:511];
  reg [7:0] LsuL1Plugin_logic_banks_1_mem_symbol1 [0:511];
  reg [7:0] LsuL1Plugin_logic_banks_1_mem_symbol2 [0:511];
  reg [7:0] LsuL1Plugin_logic_banks_1_mem_symbol3 [0:511];
  reg [7:0] LsuL1Plugin_logic_banks_1_mem_symbol4 [0:511];
  reg [7:0] LsuL1Plugin_logic_banks_1_mem_symbol5 [0:511];
  reg [7:0] LsuL1Plugin_logic_banks_1_mem_symbol6 [0:511];
  reg [7:0] LsuL1Plugin_logic_banks_1_mem_symbol7 [0:511];
  reg [7:0] _zz_LsuL1Plugin_logic_banks_1_memsymbol_read;
  reg [7:0] _zz_LsuL1Plugin_logic_banks_1_memsymbol_read_1;
  reg [7:0] _zz_LsuL1Plugin_logic_banks_1_memsymbol_read_2;
  reg [7:0] _zz_LsuL1Plugin_logic_banks_1_memsymbol_read_3;
  reg [7:0] _zz_LsuL1Plugin_logic_banks_1_memsymbol_read_4;
  reg [7:0] _zz_LsuL1Plugin_logic_banks_1_memsymbol_read_5;
  reg [7:0] _zz_LsuL1Plugin_logic_banks_1_memsymbol_read_6;
  reg [7:0] _zz_LsuL1Plugin_logic_banks_1_memsymbol_read_7;
  reg [21:0] LsuL1Plugin_logic_ways_0_mem [0:63];
  reg [21:0] LsuL1Plugin_logic_ways_1_mem [0:63];
  reg [2:0] LsuL1Plugin_logic_shared_mem [0:63];
  reg [63:0] LsuL1Plugin_logic_writeback_victimBuffer [0:7];
  (* ram_style = "distributed" *) reg [38:0] FetchL1Plugin_logic_translationStorage_logic_sl_0_ways_0 [0:63];
  (* ram_style = "distributed" *) reg [38:0] FetchL1Plugin_logic_translationStorage_logic_sl_0_ways_1 [0:63];
  (* ram_style = "distributed" *) reg [18:0] FetchL1Plugin_logic_translationStorage_logic_sl_1_ways_0 [0:63];
  (* ram_style = "distributed" *) reg [38:0] LsuPlugin_logic_translationStorage_logic_sl_0_ways_0 [0:63];
  (* ram_style = "distributed" *) reg [38:0] LsuPlugin_logic_translationStorage_logic_sl_0_ways_1 [0:63];
  (* ram_style = "distributed" *) reg [18:0] LsuPlugin_logic_translationStorage_logic_sl_1_ways_0 [0:63];
  reg [31:0] CsrRamPlugin_logic_mem [0:7];
  function [2:0] zz_FetchL1Plugin_logic_trapPort_payload_arg(input dummy);
    begin
      zz_FetchL1Plugin_logic_trapPort_payload_arg = 3'b000;
      zz_FetchL1Plugin_logic_trapPort_payload_arg[1 : 0] = 2'b10;
      zz_FetchL1Plugin_logic_trapPort_payload_arg[2 : 2] = 1'b0;
    end
  endfunction
  wire [2:0] _zz_59;

  assign _zz_when = (! FetchL1Plugin_logic_refill_slots_0_valid);
  assign _zz_early0_IntAluPlugin_logic_alu_result = (early0_IntAluPlugin_logic_alu_bitwise | _zz_early0_IntAluPlugin_logic_alu_result_1);
  assign _zz_early0_IntAluPlugin_logic_alu_result_1 = (toplevel_execute_ctrl2_down_early0_IntAluPlugin_ALU_ADD_SUB_lane0 ? toplevel_execute_ctrl2_down_early0_SrcPlugin_ADD_SUB_lane0 : 32'h0);
  assign _zz_early0_IntAluPlugin_logic_alu_result_2 = (toplevel_execute_ctrl2_down_early0_IntAluPlugin_ALU_SLTX_lane0 ? _zz_early0_IntAluPlugin_logic_alu_result_3 : 32'h0);
  assign _zz_early0_IntAluPlugin_logic_alu_result_3 = _zz_early0_IntAluPlugin_logic_alu_result_4;
  assign _zz_early0_IntAluPlugin_logic_alu_result_5 = toplevel_execute_ctrl2_down_early0_SrcPlugin_LESS_lane0;
  assign _zz_early0_IntAluPlugin_logic_alu_result_4 = {31'd0, _zz_early0_IntAluPlugin_logic_alu_result_5};
  assign _zz_early0_BarrelShifterPlugin_logic_shift_amplitude = toplevel_execute_ctrl2_down_early0_SrcPlugin_SRC2_lane0[4 : 0];
  assign _zz_early0_BarrelShifterPlugin_logic_shift_reversed = {toplevel_execute_ctrl2_down_early0_SrcPlugin_SRC1_lane0[0],{toplevel_execute_ctrl2_down_early0_SrcPlugin_SRC1_lane0[1],{toplevel_execute_ctrl2_down_early0_SrcPlugin_SRC1_lane0[2],{toplevel_execute_ctrl2_down_early0_SrcPlugin_SRC1_lane0[3],{toplevel_execute_ctrl2_down_early0_SrcPlugin_SRC1_lane0[4],{toplevel_execute_ctrl2_down_early0_SrcPlugin_SRC1_lane0[5],{toplevel_execute_ctrl2_down_early0_SrcPlugin_SRC1_lane0[6],{toplevel_execute_ctrl2_down_early0_SrcPlugin_SRC1_lane0[7],{toplevel_execute_ctrl2_down_early0_SrcPlugin_SRC1_lane0[8],{_zz_early0_BarrelShifterPlugin_logic_shift_reversed_1,{_zz_early0_BarrelShifterPlugin_logic_shift_reversed_2,_zz_early0_BarrelShifterPlugin_logic_shift_reversed_3}}}}}}}}}}};
  assign _zz_early0_BarrelShifterPlugin_logic_shift_shifted = ($signed(_zz_early0_BarrelShifterPlugin_logic_shift_shifted_1) >>> early0_BarrelShifterPlugin_logic_shift_amplitude);
  assign _zz_early0_BarrelShifterPlugin_logic_shift_shifted_1 = {(toplevel_execute_ctrl2_down_BarrelShifterPlugin_SIGNED_lane0 && toplevel_execute_ctrl2_down_early0_SrcPlugin_SRC1_lane0[31]),early0_BarrelShifterPlugin_logic_shift_reversed};
  assign _zz_early0_BarrelShifterPlugin_logic_shift_patched = {early0_BarrelShifterPlugin_logic_shift_shifted[0],{early0_BarrelShifterPlugin_logic_shift_shifted[1],{early0_BarrelShifterPlugin_logic_shift_shifted[2],{early0_BarrelShifterPlugin_logic_shift_shifted[3],{early0_BarrelShifterPlugin_logic_shift_shifted[4],{early0_BarrelShifterPlugin_logic_shift_shifted[5],{early0_BarrelShifterPlugin_logic_shift_shifted[6],{early0_BarrelShifterPlugin_logic_shift_shifted[7],{early0_BarrelShifterPlugin_logic_shift_shifted[8],{_zz_early0_BarrelShifterPlugin_logic_shift_patched_1,{_zz_early0_BarrelShifterPlugin_logic_shift_patched_2,_zz_early0_BarrelShifterPlugin_logic_shift_patched_3}}}}}}}}}}};
  assign _zz_toplevel_execute_ctrl2_down_MUL_SRC1_lane0 = {(toplevel_execute_ctrl2_down_RsUnsignedPlugin_RS1_SIGNED_lane0 && toplevel_execute_ctrl2_up_integer_RS1_lane0[31]),toplevel_execute_ctrl2_up_integer_RS1_lane0};
  assign _zz_toplevel_execute_ctrl2_down_MUL_SRC2_lane0 = {(toplevel_execute_ctrl2_down_RsUnsignedPlugin_RS2_SIGNED_lane0 && toplevel_execute_ctrl2_up_integer_RS2_lane0[31]),toplevel_execute_ctrl2_up_integer_RS2_lane0};
  assign _zz_toplevel_execute_ctrl3_down_early0_MulPlugin_logic_mul_VALUES_1_lane0_1 = ($signed(_zz_toplevel_execute_ctrl3_down_early0_MulPlugin_logic_mul_VALUES_1_lane0_2) * $signed(_zz_toplevel_execute_ctrl3_down_early0_MulPlugin_logic_mul_VALUES_1_lane0_3));
  assign _zz_toplevel_execute_ctrl3_down_early0_MulPlugin_logic_mul_VALUES_1_lane0 = {{13{_zz_toplevel_execute_ctrl3_down_early0_MulPlugin_logic_mul_VALUES_1_lane0_1[33]}}, _zz_toplevel_execute_ctrl3_down_early0_MulPlugin_logic_mul_VALUES_1_lane0_1};
  assign _zz_toplevel_execute_ctrl3_down_early0_MulPlugin_logic_mul_VALUES_1_lane0_2 = {1'b0,toplevel_execute_ctrl3_down_MUL_SRC1_lane0[16 : 0]};
  assign _zz_toplevel_execute_ctrl3_down_early0_MulPlugin_logic_mul_VALUES_1_lane0_3 = toplevel_execute_ctrl3_down_MUL_SRC2_lane0[32 : 17];
  assign _zz_toplevel_execute_ctrl3_down_early0_MulPlugin_logic_mul_VALUES_2_lane0_1 = ($signed(_zz_toplevel_execute_ctrl3_down_early0_MulPlugin_logic_mul_VALUES_2_lane0_2) * $signed(_zz_toplevel_execute_ctrl3_down_early0_MulPlugin_logic_mul_VALUES_2_lane0_3));
  assign _zz_toplevel_execute_ctrl3_down_early0_MulPlugin_logic_mul_VALUES_2_lane0 = {{13{_zz_toplevel_execute_ctrl3_down_early0_MulPlugin_logic_mul_VALUES_2_lane0_1[33]}}, _zz_toplevel_execute_ctrl3_down_early0_MulPlugin_logic_mul_VALUES_2_lane0_1};
  assign _zz_toplevel_execute_ctrl3_down_early0_MulPlugin_logic_mul_VALUES_2_lane0_2 = toplevel_execute_ctrl3_down_MUL_SRC1_lane0[32 : 17];
  assign _zz_toplevel_execute_ctrl3_down_early0_MulPlugin_logic_mul_VALUES_2_lane0_3 = {1'b0,toplevel_execute_ctrl3_down_MUL_SRC2_lane0[16 : 0]};
  assign _zz_toplevel_execute_ctrl3_down_early0_MulPlugin_logic_mul_VALUES_3_lane0_1 = ($signed(_zz_toplevel_execute_ctrl3_down_early0_MulPlugin_logic_mul_VALUES_3_lane0_2) * $signed(_zz_toplevel_execute_ctrl3_down_early0_MulPlugin_logic_mul_VALUES_3_lane0_3));
  assign _zz_toplevel_execute_ctrl3_down_early0_MulPlugin_logic_mul_VALUES_3_lane0 = _zz_toplevel_execute_ctrl3_down_early0_MulPlugin_logic_mul_VALUES_3_lane0_1[29:0];
  assign _zz_toplevel_execute_ctrl3_down_early0_MulPlugin_logic_mul_VALUES_3_lane0_2 = toplevel_execute_ctrl3_down_MUL_SRC1_lane0[32 : 17];
  assign _zz_toplevel_execute_ctrl3_down_early0_MulPlugin_logic_mul_VALUES_3_lane0_3 = toplevel_execute_ctrl3_down_MUL_SRC2_lane0[32 : 17];
  assign _zz_toplevel_execute_ctrl3_down_early0_MulPlugin_logic_steps_0_adders_0_lane0_3 = (_zz_toplevel_execute_ctrl3_down_early0_MulPlugin_logic_steps_0_adders_0_lane0_4 + _zz_toplevel_execute_ctrl3_down_early0_MulPlugin_logic_steps_0_adders_0_lane0_5);
  assign _zz_toplevel_execute_ctrl3_down_early0_MulPlugin_logic_steps_0_adders_0_lane0_4 = {2'd0, _zz_toplevel_execute_ctrl3_down_early0_MulPlugin_logic_steps_0_adders_0_lane0};
  assign _zz_toplevel_execute_ctrl3_down_early0_MulPlugin_logic_steps_0_adders_0_lane0_5 = {2'd0, _zz_toplevel_execute_ctrl3_down_early0_MulPlugin_logic_steps_0_adders_0_lane0_1};
  assign _zz_toplevel_execute_ctrl3_down_early0_MulPlugin_logic_steps_0_adders_0_lane0_6 = {2'd0, _zz_toplevel_execute_ctrl3_down_early0_MulPlugin_logic_steps_0_adders_0_lane0_2};
  assign _zz_toplevel_execute_ctrl3_down_early0_MulPlugin_logic_steps_0_adders_1_lane0_3 = (_zz_toplevel_execute_ctrl3_down_early0_MulPlugin_logic_steps_0_adders_1_lane0_4 + _zz_toplevel_execute_ctrl3_down_early0_MulPlugin_logic_steps_0_adders_1_lane0_5);
  assign _zz_toplevel_execute_ctrl3_down_early0_MulPlugin_logic_steps_0_adders_1_lane0_4 = {2'd0, _zz_toplevel_execute_ctrl3_down_early0_MulPlugin_logic_steps_0_adders_1_lane0};
  assign _zz_toplevel_execute_ctrl3_down_early0_MulPlugin_logic_steps_0_adders_1_lane0_5 = {2'd0, _zz_toplevel_execute_ctrl3_down_early0_MulPlugin_logic_steps_0_adders_1_lane0_1};
  assign _zz_toplevel_execute_ctrl3_down_early0_MulPlugin_logic_steps_0_adders_1_lane0_6 = {2'd0, _zz_toplevel_execute_ctrl3_down_early0_MulPlugin_logic_steps_0_adders_1_lane0_2};
  assign _zz_toplevel_execute_ctrl2_down_RsUnsignedPlugin_RS1_UNSIGNED_lane0_1 = toplevel_execute_ctrl2_down_RsUnsignedPlugin_RS1_REVERT_lane0;
  assign _zz_toplevel_execute_ctrl2_down_RsUnsignedPlugin_RS1_UNSIGNED_lane0 = {31'd0, _zz_toplevel_execute_ctrl2_down_RsUnsignedPlugin_RS1_UNSIGNED_lane0_1};
  assign _zz_toplevel_execute_ctrl2_down_RsUnsignedPlugin_RS2_UNSIGNED_lane0_1 = toplevel_execute_ctrl2_down_RsUnsignedPlugin_RS2_REVERT_lane0;
  assign _zz_toplevel_execute_ctrl2_down_RsUnsignedPlugin_RS2_UNSIGNED_lane0 = {31'd0, _zz_toplevel_execute_ctrl2_down_RsUnsignedPlugin_RS2_UNSIGNED_lane0_1};
  assign _zz_toplevel_execute_ctrl2_down_DivPlugin_DIV_RESULT_lane0_1 = ((early0_DivPlugin_logic_processing_divRevertResult ? (~ _zz_toplevel_execute_ctrl2_down_DivPlugin_DIV_RESULT_lane0) : _zz_toplevel_execute_ctrl2_down_DivPlugin_DIV_RESULT_lane0) + _zz_toplevel_execute_ctrl2_down_DivPlugin_DIV_RESULT_lane0_2);
  assign _zz_toplevel_execute_ctrl2_down_DivPlugin_DIV_RESULT_lane0_3 = early0_DivPlugin_logic_processing_divRevertResult;
  assign _zz_toplevel_execute_ctrl2_down_DivPlugin_DIV_RESULT_lane0_2 = {31'd0, _zz_toplevel_execute_ctrl2_down_DivPlugin_DIV_RESULT_lane0_3};
  assign _zz_late0_IntAluPlugin_logic_alu_result = (late0_IntAluPlugin_logic_alu_bitwise | _zz_late0_IntAluPlugin_logic_alu_result_1);
  assign _zz_late0_IntAluPlugin_logic_alu_result_1 = (toplevel_execute_ctrl4_down_late0_IntAluPlugin_ALU_ADD_SUB_lane0 ? toplevel_execute_ctrl4_down_late0_SrcPlugin_ADD_SUB_lane0 : 32'h0);
  assign _zz_late0_IntAluPlugin_logic_alu_result_2 = (toplevel_execute_ctrl4_down_late0_IntAluPlugin_ALU_SLTX_lane0 ? _zz_late0_IntAluPlugin_logic_alu_result_3 : 32'h0);
  assign _zz_late0_IntAluPlugin_logic_alu_result_3 = _zz_late0_IntAluPlugin_logic_alu_result_4;
  assign _zz_late0_IntAluPlugin_logic_alu_result_5 = toplevel_execute_ctrl4_down_late0_SrcPlugin_LESS_lane0;
  assign _zz_late0_IntAluPlugin_logic_alu_result_4 = {31'd0, _zz_late0_IntAluPlugin_logic_alu_result_5};
  assign _zz_late0_BarrelShifterPlugin_logic_shift_amplitude = toplevel_execute_ctrl4_down_late0_SrcPlugin_SRC2_lane0[4 : 0];
  assign _zz_late0_BarrelShifterPlugin_logic_shift_reversed = {toplevel_execute_ctrl4_down_late0_SrcPlugin_SRC1_lane0[0],{toplevel_execute_ctrl4_down_late0_SrcPlugin_SRC1_lane0[1],{toplevel_execute_ctrl4_down_late0_SrcPlugin_SRC1_lane0[2],{toplevel_execute_ctrl4_down_late0_SrcPlugin_SRC1_lane0[3],{toplevel_execute_ctrl4_down_late0_SrcPlugin_SRC1_lane0[4],{toplevel_execute_ctrl4_down_late0_SrcPlugin_SRC1_lane0[5],{toplevel_execute_ctrl4_down_late0_SrcPlugin_SRC1_lane0[6],{toplevel_execute_ctrl4_down_late0_SrcPlugin_SRC1_lane0[7],{toplevel_execute_ctrl4_down_late0_SrcPlugin_SRC1_lane0[8],{_zz_late0_BarrelShifterPlugin_logic_shift_reversed_1,{_zz_late0_BarrelShifterPlugin_logic_shift_reversed_2,_zz_late0_BarrelShifterPlugin_logic_shift_reversed_3}}}}}}}}}}};
  assign _zz_late0_BarrelShifterPlugin_logic_shift_shifted = ($signed(_zz_late0_BarrelShifterPlugin_logic_shift_shifted_1) >>> late0_BarrelShifterPlugin_logic_shift_amplitude);
  assign _zz_late0_BarrelShifterPlugin_logic_shift_shifted_1 = {(toplevel_execute_ctrl4_down_BarrelShifterPlugin_SIGNED_lane0 && toplevel_execute_ctrl4_down_late0_SrcPlugin_SRC1_lane0[31]),late0_BarrelShifterPlugin_logic_shift_reversed};
  assign _zz_late0_BarrelShifterPlugin_logic_shift_patched = {late0_BarrelShifterPlugin_logic_shift_shifted[0],{late0_BarrelShifterPlugin_logic_shift_shifted[1],{late0_BarrelShifterPlugin_logic_shift_shifted[2],{late0_BarrelShifterPlugin_logic_shift_shifted[3],{late0_BarrelShifterPlugin_logic_shift_shifted[4],{late0_BarrelShifterPlugin_logic_shift_shifted[5],{late0_BarrelShifterPlugin_logic_shift_shifted[6],{late0_BarrelShifterPlugin_logic_shift_shifted[7],{late0_BarrelShifterPlugin_logic_shift_shifted[8],{_zz_late0_BarrelShifterPlugin_logic_shift_patched_1,{_zz_late0_BarrelShifterPlugin_logic_shift_patched_2,_zz_late0_BarrelShifterPlugin_logic_shift_patched_3}}}}}}}}}}};
  assign _zz_early1_IntAluPlugin_logic_alu_result = (early1_IntAluPlugin_logic_alu_bitwise | _zz_early1_IntAluPlugin_logic_alu_result_1);
  assign _zz_early1_IntAluPlugin_logic_alu_result_1 = (toplevel_execute_ctrl2_down_early1_IntAluPlugin_ALU_ADD_SUB_lane1 ? toplevel_execute_ctrl2_down_early1_SrcPlugin_ADD_SUB_lane1 : 32'h0);
  assign _zz_early1_IntAluPlugin_logic_alu_result_2 = (toplevel_execute_ctrl2_down_early1_IntAluPlugin_ALU_SLTX_lane1 ? _zz_early1_IntAluPlugin_logic_alu_result_3 : 32'h0);
  assign _zz_early1_IntAluPlugin_logic_alu_result_3 = _zz_early1_IntAluPlugin_logic_alu_result_4;
  assign _zz_early1_IntAluPlugin_logic_alu_result_5 = toplevel_execute_ctrl2_down_early1_SrcPlugin_LESS_lane1;
  assign _zz_early1_IntAluPlugin_logic_alu_result_4 = {31'd0, _zz_early1_IntAluPlugin_logic_alu_result_5};
  assign _zz_early1_BarrelShifterPlugin_logic_shift_amplitude = toplevel_execute_ctrl2_down_early1_SrcPlugin_SRC2_lane1[4 : 0];
  assign _zz_early1_BarrelShifterPlugin_logic_shift_reversed = {toplevel_execute_ctrl2_down_early1_SrcPlugin_SRC1_lane1[0],{toplevel_execute_ctrl2_down_early1_SrcPlugin_SRC1_lane1[1],{toplevel_execute_ctrl2_down_early1_SrcPlugin_SRC1_lane1[2],{toplevel_execute_ctrl2_down_early1_SrcPlugin_SRC1_lane1[3],{toplevel_execute_ctrl2_down_early1_SrcPlugin_SRC1_lane1[4],{toplevel_execute_ctrl2_down_early1_SrcPlugin_SRC1_lane1[5],{toplevel_execute_ctrl2_down_early1_SrcPlugin_SRC1_lane1[6],{toplevel_execute_ctrl2_down_early1_SrcPlugin_SRC1_lane1[7],{toplevel_execute_ctrl2_down_early1_SrcPlugin_SRC1_lane1[8],{_zz_early1_BarrelShifterPlugin_logic_shift_reversed_1,{_zz_early1_BarrelShifterPlugin_logic_shift_reversed_2,_zz_early1_BarrelShifterPlugin_logic_shift_reversed_3}}}}}}}}}}};
  assign _zz_early1_BarrelShifterPlugin_logic_shift_shifted = ($signed(_zz_early1_BarrelShifterPlugin_logic_shift_shifted_1) >>> early1_BarrelShifterPlugin_logic_shift_amplitude);
  assign _zz_early1_BarrelShifterPlugin_logic_shift_shifted_1 = {(toplevel_execute_ctrl2_down_BarrelShifterPlugin_SIGNED_lane1 && toplevel_execute_ctrl2_down_early1_SrcPlugin_SRC1_lane1[31]),early1_BarrelShifterPlugin_logic_shift_reversed};
  assign _zz_early1_BarrelShifterPlugin_logic_shift_patched = {early1_BarrelShifterPlugin_logic_shift_shifted[0],{early1_BarrelShifterPlugin_logic_shift_shifted[1],{early1_BarrelShifterPlugin_logic_shift_shifted[2],{early1_BarrelShifterPlugin_logic_shift_shifted[3],{early1_BarrelShifterPlugin_logic_shift_shifted[4],{early1_BarrelShifterPlugin_logic_shift_shifted[5],{early1_BarrelShifterPlugin_logic_shift_shifted[6],{early1_BarrelShifterPlugin_logic_shift_shifted[7],{early1_BarrelShifterPlugin_logic_shift_shifted[8],{_zz_early1_BarrelShifterPlugin_logic_shift_patched_1,{_zz_early1_BarrelShifterPlugin_logic_shift_patched_2,_zz_early1_BarrelShifterPlugin_logic_shift_patched_3}}}}}}}}}}};
  assign _zz_late1_IntAluPlugin_logic_alu_result = (late1_IntAluPlugin_logic_alu_bitwise | _zz_late1_IntAluPlugin_logic_alu_result_1);
  assign _zz_late1_IntAluPlugin_logic_alu_result_1 = (toplevel_execute_ctrl4_down_late1_IntAluPlugin_ALU_ADD_SUB_lane1 ? toplevel_execute_ctrl4_down_late1_SrcPlugin_ADD_SUB_lane1 : 32'h0);
  assign _zz_late1_IntAluPlugin_logic_alu_result_2 = (toplevel_execute_ctrl4_down_late1_IntAluPlugin_ALU_SLTX_lane1 ? _zz_late1_IntAluPlugin_logic_alu_result_3 : 32'h0);
  assign _zz_late1_IntAluPlugin_logic_alu_result_3 = _zz_late1_IntAluPlugin_logic_alu_result_4;
  assign _zz_late1_IntAluPlugin_logic_alu_result_5 = toplevel_execute_ctrl4_down_late1_SrcPlugin_LESS_lane1;
  assign _zz_late1_IntAluPlugin_logic_alu_result_4 = {31'd0, _zz_late1_IntAluPlugin_logic_alu_result_5};
  assign _zz_late1_BarrelShifterPlugin_logic_shift_amplitude = toplevel_execute_ctrl4_down_late1_SrcPlugin_SRC2_lane1[4 : 0];
  assign _zz_late1_BarrelShifterPlugin_logic_shift_reversed = {toplevel_execute_ctrl4_down_late1_SrcPlugin_SRC1_lane1[0],{toplevel_execute_ctrl4_down_late1_SrcPlugin_SRC1_lane1[1],{toplevel_execute_ctrl4_down_late1_SrcPlugin_SRC1_lane1[2],{toplevel_execute_ctrl4_down_late1_SrcPlugin_SRC1_lane1[3],{toplevel_execute_ctrl4_down_late1_SrcPlugin_SRC1_lane1[4],{toplevel_execute_ctrl4_down_late1_SrcPlugin_SRC1_lane1[5],{toplevel_execute_ctrl4_down_late1_SrcPlugin_SRC1_lane1[6],{toplevel_execute_ctrl4_down_late1_SrcPlugin_SRC1_lane1[7],{toplevel_execute_ctrl4_down_late1_SrcPlugin_SRC1_lane1[8],{_zz_late1_BarrelShifterPlugin_logic_shift_reversed_1,{_zz_late1_BarrelShifterPlugin_logic_shift_reversed_2,_zz_late1_BarrelShifterPlugin_logic_shift_reversed_3}}}}}}}}}}};
  assign _zz_late1_BarrelShifterPlugin_logic_shift_shifted = ($signed(_zz_late1_BarrelShifterPlugin_logic_shift_shifted_1) >>> late1_BarrelShifterPlugin_logic_shift_amplitude);
  assign _zz_late1_BarrelShifterPlugin_logic_shift_shifted_1 = {(toplevel_execute_ctrl4_down_BarrelShifterPlugin_SIGNED_lane1 && toplevel_execute_ctrl4_down_late1_SrcPlugin_SRC1_lane1[31]),late1_BarrelShifterPlugin_logic_shift_reversed};
  assign _zz_late1_BarrelShifterPlugin_logic_shift_patched = {late1_BarrelShifterPlugin_logic_shift_shifted[0],{late1_BarrelShifterPlugin_logic_shift_shifted[1],{late1_BarrelShifterPlugin_logic_shift_shifted[2],{late1_BarrelShifterPlugin_logic_shift_shifted[3],{late1_BarrelShifterPlugin_logic_shift_shifted[4],{late1_BarrelShifterPlugin_logic_shift_shifted[5],{late1_BarrelShifterPlugin_logic_shift_shifted[6],{late1_BarrelShifterPlugin_logic_shift_shifted[7],{late1_BarrelShifterPlugin_logic_shift_shifted[8],{_zz_late1_BarrelShifterPlugin_logic_shift_patched_1,{_zz_late1_BarrelShifterPlugin_logic_shift_patched_2,_zz_late1_BarrelShifterPlugin_logic_shift_patched_3}}}}}}}}}}};
  assign _zz_early0_BranchPlugin_pcCalc_target_b = {{{{toplevel_execute_ctrl2_down_Decode_UOP_lane0[31],toplevel_execute_ctrl2_down_Decode_UOP_lane0[19 : 12]},toplevel_execute_ctrl2_down_Decode_UOP_lane0[20]},toplevel_execute_ctrl2_down_Decode_UOP_lane0[30 : 21]},1'b0};
  assign _zz_early0_BranchPlugin_pcCalc_target_b_1 = toplevel_execute_ctrl2_down_Decode_UOP_lane0[31 : 20];
  assign _zz_early0_BranchPlugin_pcCalc_target_b_2 = {{{{toplevel_execute_ctrl2_down_Decode_UOP_lane0[31],toplevel_execute_ctrl2_down_Decode_UOP_lane0[7]},toplevel_execute_ctrl2_down_Decode_UOP_lane0[30 : 25]},toplevel_execute_ctrl2_down_Decode_UOP_lane0[11 : 8]},1'b0};
  assign _zz_toplevel_execute_ctrl2_down_early0_BranchPlugin_pcCalc_PC_TRUE_lane0 = ($signed(early0_BranchPlugin_pcCalc_target_a) + $signed(early0_BranchPlugin_pcCalc_target_b));
  assign _zz_toplevel_execute_ctrl2_down_early0_BranchPlugin_pcCalc_PC_FALSE_lane0_1 = ({1'd0,early0_BranchPlugin_pcCalc_slices} <<< 1'd1);
  assign _zz_toplevel_execute_ctrl2_down_early0_BranchPlugin_pcCalc_PC_FALSE_lane0 = {29'd0, _zz_toplevel_execute_ctrl2_down_early0_BranchPlugin_pcCalc_PC_FALSE_lane0_1};
  assign _zz_toplevel_execute_ctrl2_down_early0_BranchPlugin_pcCalc_PC_LAST_SLICE_lane0_1 = ({1'd0,toplevel_execute_ctrl2_down_Decode_INSTRUCTION_SLICE_COUNT_lane0} <<< 1'd1);
  assign _zz_toplevel_execute_ctrl2_down_early0_BranchPlugin_pcCalc_PC_LAST_SLICE_lane0 = {30'd0, _zz_toplevel_execute_ctrl2_down_early0_BranchPlugin_pcCalc_PC_LAST_SLICE_lane0_1};
  assign _zz_early1_BranchPlugin_pcCalc_target_b = {{{{toplevel_execute_ctrl2_down_Decode_UOP_lane1[31],toplevel_execute_ctrl2_down_Decode_UOP_lane1[19 : 12]},toplevel_execute_ctrl2_down_Decode_UOP_lane1[20]},toplevel_execute_ctrl2_down_Decode_UOP_lane1[30 : 21]},1'b0};
  assign _zz_early1_BranchPlugin_pcCalc_target_b_1 = toplevel_execute_ctrl2_down_Decode_UOP_lane1[31 : 20];
  assign _zz_early1_BranchPlugin_pcCalc_target_b_2 = {{{{toplevel_execute_ctrl2_down_Decode_UOP_lane1[31],toplevel_execute_ctrl2_down_Decode_UOP_lane1[7]},toplevel_execute_ctrl2_down_Decode_UOP_lane1[30 : 25]},toplevel_execute_ctrl2_down_Decode_UOP_lane1[11 : 8]},1'b0};
  assign _zz_toplevel_execute_ctrl2_down_early1_BranchPlugin_pcCalc_PC_TRUE_lane1 = ($signed(early1_BranchPlugin_pcCalc_target_a) + $signed(early1_BranchPlugin_pcCalc_target_b));
  assign _zz_toplevel_execute_ctrl2_down_early1_BranchPlugin_pcCalc_PC_FALSE_lane1_1 = ({1'd0,early1_BranchPlugin_pcCalc_slices} <<< 1'd1);
  assign _zz_toplevel_execute_ctrl2_down_early1_BranchPlugin_pcCalc_PC_FALSE_lane1 = {29'd0, _zz_toplevel_execute_ctrl2_down_early1_BranchPlugin_pcCalc_PC_FALSE_lane1_1};
  assign _zz_toplevel_execute_ctrl2_down_early1_BranchPlugin_pcCalc_PC_LAST_SLICE_lane1_1 = ({1'd0,toplevel_execute_ctrl2_down_Decode_INSTRUCTION_SLICE_COUNT_lane1} <<< 1'd1);
  assign _zz_toplevel_execute_ctrl2_down_early1_BranchPlugin_pcCalc_PC_LAST_SLICE_lane1 = {30'd0, _zz_toplevel_execute_ctrl2_down_early1_BranchPlugin_pcCalc_PC_LAST_SLICE_lane1_1};
  assign _zz_fetch_logic_ctrls_2_down_AlignerPlugin_logic_FETCH_LAST = (4'b0001 <<< fetch_logic_ctrls_2_down_Prediction_WORD_JUMP_SLICE);
  assign _zz_AlignerPlugin_logic_extractors_0_redo_8 = ((((_zz_AlignerPlugin_logic_extractors_0_redo ? _zz_AlignerPlugin_logic_extractors_0_redo_9 : _zz_AlignerPlugin_logic_extractors_0_redo_10) | (_zz_AlignerPlugin_logic_extractors_0_redo_1 ? _zz_AlignerPlugin_logic_extractors_0_redo_11 : _zz_AlignerPlugin_logic_extractors_0_redo_12)) | ((_zz_AlignerPlugin_logic_extractors_0_redo_2 ? _zz_AlignerPlugin_logic_extractors_0_redo_13 : _zz_AlignerPlugin_logic_extractors_0_redo_14) | (_zz_AlignerPlugin_logic_extractors_0_redo_3 ? _zz_AlignerPlugin_logic_extractors_0_redo_15 : _zz_AlignerPlugin_logic_extractors_0_redo_16))) | (((_zz_AlignerPlugin_logic_extractors_0_redo_4 ? _zz_AlignerPlugin_logic_extractors_0_redo_17 : _zz_AlignerPlugin_logic_extractors_0_redo_18) | (_zz_AlignerPlugin_logic_extractors_0_redo_5 ? _zz_AlignerPlugin_logic_extractors_0_redo_19 : _zz_AlignerPlugin_logic_extractors_0_redo_20)) | ((_zz_AlignerPlugin_logic_extractors_0_redo_6 ? _zz_AlignerPlugin_logic_extractors_0_redo_21 : _zz_AlignerPlugin_logic_extractors_0_redo_22) | (_zz_AlignerPlugin_logic_extractors_0_redo_7 ? _zz_AlignerPlugin_logic_extractors_0_redo_23 : _zz_AlignerPlugin_logic_extractors_0_redo_24))));
  assign _zz_AlignerPlugin_logic_extractors_1_redo_7 = ((((_zz_AlignerPlugin_logic_extractors_1_redo ? _zz_AlignerPlugin_logic_extractors_1_redo_8 : _zz_AlignerPlugin_logic_extractors_1_redo_9) | (_zz_AlignerPlugin_logic_extractors_1_redo_1 ? _zz_AlignerPlugin_logic_extractors_1_redo_10 : _zz_AlignerPlugin_logic_extractors_1_redo_11)) | ((_zz_AlignerPlugin_logic_extractors_1_redo_2 ? _zz_AlignerPlugin_logic_extractors_1_redo_12 : _zz_AlignerPlugin_logic_extractors_1_redo_13) | (_zz_AlignerPlugin_logic_extractors_1_redo_3 ? _zz_AlignerPlugin_logic_extractors_1_redo_14 : _zz_AlignerPlugin_logic_extractors_1_redo_15))) | (((_zz_AlignerPlugin_logic_extractors_1_redo_4 ? _zz_AlignerPlugin_logic_extractors_1_redo_16 : _zz_AlignerPlugin_logic_extractors_1_redo_17) | (_zz_AlignerPlugin_logic_extractors_1_redo_5 ? _zz_AlignerPlugin_logic_extractors_1_redo_18 : _zz_AlignerPlugin_logic_extractors_1_redo_19)) | (_zz_AlignerPlugin_logic_extractors_1_redo_6 ? AlignerPlugin_logic_scanners_7_redo : 1'b0)));
  assign _zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_26 = {{_zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_10,AlignerPlugin_logic_extractors_0_ctx_instruction[6 : 2]},12'h0};
  assign _zz__zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_22_1 = {AlignerPlugin_logic_extractors_0_ctx_instruction[12],AlignerPlugin_logic_extractors_0_ctx_instruction[6 : 2]};
  assign _zz__zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_22 = {6'd0, _zz__zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_22_1};
  assign _zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_35 = {{{4'b0000,AlignerPlugin_logic_extractors_0_ctx_instruction[8 : 7]},AlignerPlugin_logic_extractors_0_ctx_instruction[12 : 9]},2'b00};
  assign _zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_36 = {{{4'b0000,AlignerPlugin_logic_extractors_0_ctx_instruction[8 : 7]},AlignerPlugin_logic_extractors_0_ctx_instruction[12 : 9]},2'b00};
  assign _zz__zz_toplevel_decode_ctrls_0_up_Decode_INSTRUCTION_SLICE_COUNT_0_5 = {_zz_toplevel_decode_ctrls_0_up_Decode_INSTRUCTION_SLICE_COUNT_0_4[0],_zz_toplevel_decode_ctrls_0_up_Decode_INSTRUCTION_SLICE_COUNT_0_4[1]};
  assign _zz_AlignerPlugin_logic_feeder_lanes_0_onBtb_pcLastSlice = {1'd0, toplevel_decode_ctrls_0_up_Decode_INSTRUCTION_SLICE_COUNT_0};
  assign _zz_AlignerPlugin_logic_feeder_lanes_1_withRvc_dec_inst_26 = {{_zz_AlignerPlugin_logic_feeder_lanes_1_withRvc_dec_inst_10,AlignerPlugin_logic_extractors_1_ctx_instruction[6 : 2]},12'h0};
  assign _zz__zz_AlignerPlugin_logic_feeder_lanes_1_withRvc_dec_inst_22_1 = {AlignerPlugin_logic_extractors_1_ctx_instruction[12],AlignerPlugin_logic_extractors_1_ctx_instruction[6 : 2]};
  assign _zz__zz_AlignerPlugin_logic_feeder_lanes_1_withRvc_dec_inst_22 = {6'd0, _zz__zz_AlignerPlugin_logic_feeder_lanes_1_withRvc_dec_inst_22_1};
  assign _zz_AlignerPlugin_logic_feeder_lanes_1_withRvc_dec_inst_35 = {{{4'b0000,AlignerPlugin_logic_extractors_1_ctx_instruction[8 : 7]},AlignerPlugin_logic_extractors_1_ctx_instruction[12 : 9]},2'b00};
  assign _zz_AlignerPlugin_logic_feeder_lanes_1_withRvc_dec_inst_36 = {{{4'b0000,AlignerPlugin_logic_extractors_1_ctx_instruction[8 : 7]},AlignerPlugin_logic_extractors_1_ctx_instruction[12 : 9]},2'b00};
  assign _zz__zz_toplevel_decode_ctrls_0_up_Decode_INSTRUCTION_SLICE_COUNT_1_5 = {_zz_toplevel_decode_ctrls_0_up_Decode_INSTRUCTION_SLICE_COUNT_1_4[0],_zz_toplevel_decode_ctrls_0_up_Decode_INSTRUCTION_SLICE_COUNT_1_4[1]};
  assign _zz_toplevel_decode_ctrls_0_up_Decode_DOP_ID_1_1 = toplevel_decode_ctrls_0_up_LANE_SEL_0;
  assign _zz_toplevel_decode_ctrls_0_up_Decode_DOP_ID_1 = {9'd0, _zz_toplevel_decode_ctrls_0_up_Decode_DOP_ID_1_1};
  assign _zz_AlignerPlugin_logic_feeder_lanes_1_onBtb_pcLastSlice = {1'd0, toplevel_decode_ctrls_0_up_Decode_INSTRUCTION_SLICE_COUNT_1};
  assign _zz_FetchL1Plugin_logic_hits_w_0_indirect_bypassHits = (fetch_logic_ctrls_1_down_Fetch_WORD_PC >>> 4'd12);
  assign _zz_FetchL1Plugin_logic_hits_w_1_indirect_bypassHits = (fetch_logic_ctrls_1_down_Fetch_WORD_PC >>> 4'd12);
  assign _zz_FetchL1Plugin_logic_ctrl_dataAccessFault = ((fetch_logic_ctrls_2_down_FetchL1Plugin_logic_WAYS_HITS_0 ? fetch_logic_ctrls_2_down_FetchL1Plugin_logic_WAYS_TAGS_0_error : 1'b0) | (fetch_logic_ctrls_2_down_FetchL1Plugin_logic_WAYS_HITS_1 ? fetch_logic_ctrls_2_down_FetchL1Plugin_logic_WAYS_TAGS_1_error : 1'b0));
  assign _zz_FetchL1Plugin_logic_plru_write_payload_data_0 = 1'b0;
  assign _zz_BtbPlugin_logic_ras_ptr_push = (BtbPlugin_logic_ras_ptr_push + _zz_BtbPlugin_logic_ras_ptr_push_1);
  assign _zz_BtbPlugin_logic_ras_ptr_push_2 = BtbPlugin_logic_ras_ptr_pushIt;
  assign _zz_BtbPlugin_logic_ras_ptr_push_1 = {1'd0, _zz_BtbPlugin_logic_ras_ptr_push_2};
  assign _zz_BtbPlugin_logic_ras_ptr_push_4 = BtbPlugin_logic_ras_ptr_popIt;
  assign _zz_BtbPlugin_logic_ras_ptr_push_3 = {1'd0, _zz_BtbPlugin_logic_ras_ptr_push_4};
  assign _zz_BtbPlugin_logic_ras_ptr_pop_aheadValue = (BtbPlugin_logic_ras_ptr_pop + _zz_BtbPlugin_logic_ras_ptr_pop_aheadValue_1);
  assign _zz_BtbPlugin_logic_ras_ptr_pop_aheadValue_2 = BtbPlugin_logic_ras_ptr_pushIt;
  assign _zz_BtbPlugin_logic_ras_ptr_pop_aheadValue_1 = {1'd0, _zz_BtbPlugin_logic_ras_ptr_pop_aheadValue_2};
  assign _zz_BtbPlugin_logic_ras_ptr_pop_aheadValue_4 = BtbPlugin_logic_ras_ptr_popIt;
  assign _zz_BtbPlugin_logic_ras_ptr_pop_aheadValue_3 = {1'd0, _zz_BtbPlugin_logic_ras_ptr_pop_aheadValue_4};
  assign _zz_WhiteboxerPlugin_logic_decodes_0_pc = {32'd0, toplevel_decode_ctrls_0_down_PC_0};
  assign _zz_WhiteboxerPlugin_logic_decodes_1_pc = {32'd0, toplevel_decode_ctrls_0_down_PC_1};
  assign _zz_early0_BranchPlugin_logic_alu_expectedMsb = toplevel_execute_ctrl2_down_early0_SrcPlugin_SRC1_lane0;
  assign _zz_early0_BranchPlugin_logic_jumpLogic_history_fromFetch_shifter_1 = {early0_BranchPlugin_logic_jumpLogic_history_fromFetch_shifter,toplevel_execute_ctrl3_down_Prediction_ALIGNED_SLICES_TAKEN_lane0[0]};
  assign _zz_early0_BranchPlugin_logic_jumpLogic_history_fromFetch_shifter_2 = {early0_BranchPlugin_logic_jumpLogic_history_fromFetch_shifter_1,toplevel_execute_ctrl3_down_Prediction_ALIGNED_SLICES_TAKEN_lane0[1]};
  assign _zz_early0_BranchPlugin_logic_jumpLogic_history_fromFetch_shifter_3 = {early0_BranchPlugin_logic_jumpLogic_history_fromFetch_shifter_2,toplevel_execute_ctrl3_down_Prediction_ALIGNED_SLICES_TAKEN_lane0[2]};
  assign _zz_early0_BranchPlugin_logic_jumpLogic_history_fromFetch_shifter_4 = {early0_BranchPlugin_logic_jumpLogic_history_fromFetch_shifter_3,toplevel_execute_ctrl3_down_early0_BranchPlugin_logic_jumpLogic_COND_lane0};
  assign _zz_early0_EnvPlugin_logic_trapPort_payload_code = {2'd0, early0_EnvPlugin_logic_exe_privilege};
  assign _zz_early1_BranchPlugin_logic_alu_expectedMsb = toplevel_execute_ctrl2_down_early1_SrcPlugin_SRC1_lane1;
  assign _zz_early1_BranchPlugin_logic_jumpLogic_history_fromFetch_shifter_1 = {early1_BranchPlugin_logic_jumpLogic_history_fromFetch_shifter,toplevel_execute_ctrl3_down_Prediction_ALIGNED_SLICES_TAKEN_lane1[0]};
  assign _zz_early1_BranchPlugin_logic_jumpLogic_history_fromFetch_shifter_2 = {early1_BranchPlugin_logic_jumpLogic_history_fromFetch_shifter_1,toplevel_execute_ctrl3_down_Prediction_ALIGNED_SLICES_TAKEN_lane1[1]};
  assign _zz_early1_BranchPlugin_logic_jumpLogic_history_fromFetch_shifter_3 = {early1_BranchPlugin_logic_jumpLogic_history_fromFetch_shifter_2,toplevel_execute_ctrl3_down_Prediction_ALIGNED_SLICES_TAKEN_lane1[2]};
  assign _zz_early1_BranchPlugin_logic_jumpLogic_history_fromFetch_shifter_4 = {early1_BranchPlugin_logic_jumpLogic_history_fromFetch_shifter_3,toplevel_execute_ctrl3_down_early1_BranchPlugin_logic_jumpLogic_COND_lane1};
  assign _zz__zz_toplevel_execute_ctrl1_down_early0_SrcPlugin_SRC2_lane0 = toplevel_execute_ctrl1_down_Decode_UOP_lane0[31 : 20];
  assign _zz__zz_toplevel_execute_ctrl1_down_early0_SrcPlugin_SRC2_lane0_1 = {toplevel_execute_ctrl1_down_Decode_UOP_lane0[31 : 25],toplevel_execute_ctrl1_down_Decode_UOP_lane0[11 : 7]};
  assign _zz_toplevel_execute_ctrl2_down_early0_SrcPlugin_ADD_SUB_lane0 = ($signed(toplevel_execute_ctrl2_down_early0_SrcPlugin_SRC1_lane0) + $signed(early0_SrcPlugin_logic_addsub_combined_rs2Patched));
  assign _zz_toplevel_execute_ctrl2_down_early0_SrcPlugin_ADD_SUB_lane0_1 = _zz_toplevel_execute_ctrl2_down_early0_SrcPlugin_ADD_SUB_lane0_2;
  assign _zz_toplevel_execute_ctrl2_down_early0_SrcPlugin_ADD_SUB_lane0_3 = toplevel_execute_ctrl2_down_SrcStageables_REVERT_lane0;
  assign _zz_toplevel_execute_ctrl2_down_early0_SrcPlugin_ADD_SUB_lane0_2 = {31'd0, _zz_toplevel_execute_ctrl2_down_early0_SrcPlugin_ADD_SUB_lane0_3};
  assign _zz__zz_toplevel_execute_ctrl3_down_late0_SrcPlugin_SRC2_lane0 = toplevel_execute_ctrl3_down_Decode_UOP_lane0[31 : 20];
  assign _zz_toplevel_execute_ctrl4_down_late0_SrcPlugin_ADD_SUB_lane0 = ($signed(toplevel_execute_ctrl4_down_late0_SrcPlugin_SRC1_lane0) + $signed(late0_SrcPlugin_logic_addsub_combined_rs2Patched));
  assign _zz_toplevel_execute_ctrl4_down_late0_SrcPlugin_ADD_SUB_lane0_1 = _zz_toplevel_execute_ctrl4_down_late0_SrcPlugin_ADD_SUB_lane0_2;
  assign _zz_toplevel_execute_ctrl4_down_late0_SrcPlugin_ADD_SUB_lane0_3 = toplevel_execute_ctrl4_down_SrcStageables_REVERT_lane0;
  assign _zz_toplevel_execute_ctrl4_down_late0_SrcPlugin_ADD_SUB_lane0_2 = {31'd0, _zz_toplevel_execute_ctrl4_down_late0_SrcPlugin_ADD_SUB_lane0_3};
  assign _zz__zz_toplevel_execute_ctrl1_down_early1_SrcPlugin_SRC2_lane1 = toplevel_execute_ctrl1_down_Decode_UOP_lane1[31 : 20];
  assign _zz_toplevel_execute_ctrl2_down_early1_SrcPlugin_ADD_SUB_lane1 = ($signed(toplevel_execute_ctrl2_down_early1_SrcPlugin_SRC1_lane1) + $signed(early1_SrcPlugin_logic_addsub_combined_rs2Patched));
  assign _zz_toplevel_execute_ctrl2_down_early1_SrcPlugin_ADD_SUB_lane1_1 = _zz_toplevel_execute_ctrl2_down_early1_SrcPlugin_ADD_SUB_lane1_2;
  assign _zz_toplevel_execute_ctrl2_down_early1_SrcPlugin_ADD_SUB_lane1_3 = toplevel_execute_ctrl2_down_SrcStageables_REVERT_lane1;
  assign _zz_toplevel_execute_ctrl2_down_early1_SrcPlugin_ADD_SUB_lane1_2 = {31'd0, _zz_toplevel_execute_ctrl2_down_early1_SrcPlugin_ADD_SUB_lane1_3};
  assign _zz__zz_toplevel_execute_ctrl3_down_late1_SrcPlugin_SRC2_lane1 = toplevel_execute_ctrl3_down_Decode_UOP_lane1[31 : 20];
  assign _zz_toplevel_execute_ctrl4_down_late1_SrcPlugin_ADD_SUB_lane1 = ($signed(toplevel_execute_ctrl4_down_late1_SrcPlugin_SRC1_lane1) + $signed(late1_SrcPlugin_logic_addsub_combined_rs2Patched));
  assign _zz_toplevel_execute_ctrl4_down_late1_SrcPlugin_ADD_SUB_lane1_1 = _zz_toplevel_execute_ctrl4_down_late1_SrcPlugin_ADD_SUB_lane1_2;
  assign _zz_toplevel_execute_ctrl4_down_late1_SrcPlugin_ADD_SUB_lane1_3 = toplevel_execute_ctrl4_down_SrcStageables_REVERT_lane1;
  assign _zz_toplevel_execute_ctrl4_down_late1_SrcPlugin_ADD_SUB_lane1_2 = {31'd0, _zz_toplevel_execute_ctrl4_down_late1_SrcPlugin_ADD_SUB_lane1_3};
  assign _zz_late0_BranchPlugin_logic_alu_expectedMsb = toplevel_execute_ctrl4_down_late0_SrcPlugin_SRC1_lane0;
  assign _zz_late0_BranchPlugin_logic_jumpLogic_history_fromFetch_shifter_1 = {late0_BranchPlugin_logic_jumpLogic_history_fromFetch_shifter,toplevel_execute_ctrl4_down_Prediction_ALIGNED_SLICES_TAKEN_lane0[0]};
  assign _zz_late0_BranchPlugin_logic_jumpLogic_history_fromFetch_shifter_2 = {late0_BranchPlugin_logic_jumpLogic_history_fromFetch_shifter_1,toplevel_execute_ctrl4_down_Prediction_ALIGNED_SLICES_TAKEN_lane0[1]};
  assign _zz_late0_BranchPlugin_logic_jumpLogic_history_fromFetch_shifter_3 = {late0_BranchPlugin_logic_jumpLogic_history_fromFetch_shifter_2,toplevel_execute_ctrl4_down_Prediction_ALIGNED_SLICES_TAKEN_lane0[2]};
  assign _zz_late0_BranchPlugin_logic_jumpLogic_history_fromFetch_shifter_4 = {late0_BranchPlugin_logic_jumpLogic_history_fromFetch_shifter_3,toplevel_execute_ctrl4_down_late0_BranchPlugin_logic_jumpLogic_COND_lane0};
  assign _zz_late1_BranchPlugin_logic_alu_expectedMsb = toplevel_execute_ctrl4_down_late1_SrcPlugin_SRC1_lane1;
  assign _zz_late1_BranchPlugin_logic_jumpLogic_history_fromFetch_shifter_1 = {late1_BranchPlugin_logic_jumpLogic_history_fromFetch_shifter,toplevel_execute_ctrl4_down_Prediction_ALIGNED_SLICES_TAKEN_lane1[0]};
  assign _zz_late1_BranchPlugin_logic_jumpLogic_history_fromFetch_shifter_2 = {late1_BranchPlugin_logic_jumpLogic_history_fromFetch_shifter_1,toplevel_execute_ctrl4_down_Prediction_ALIGNED_SLICES_TAKEN_lane1[1]};
  assign _zz_late1_BranchPlugin_logic_jumpLogic_history_fromFetch_shifter_3 = {late1_BranchPlugin_logic_jumpLogic_history_fromFetch_shifter_2,toplevel_execute_ctrl4_down_Prediction_ALIGNED_SLICES_TAKEN_lane1[2]};
  assign _zz_late1_BranchPlugin_logic_jumpLogic_history_fromFetch_shifter_4 = {late1_BranchPlugin_logic_jumpLogic_history_fromFetch_shifter_3,toplevel_execute_ctrl4_down_late1_BranchPlugin_logic_jumpLogic_COND_lane1};
  assign _zz_BtbPlugin_logic_onLearn_port_payload_address = (LearnPlugin_logic_learn_payload_pcOnLastSlice >>> 2'd3);
  assign _zz_toplevel_decode_ctrls_1_down_RS1_ENABLE_0 = (|{((toplevel_decode_ctrls_1_down_Decode_INSTRUCTION_0 & 32'h00000044) == 32'h0),{_zz_toplevel_decode_ctrls_1_down_DispatchPlugin_MAY_FLUSH_0,{((toplevel_decode_ctrls_1_down_Decode_INSTRUCTION_0 & 32'h00006004) == 32'h00002000),{((toplevel_decode_ctrls_1_down_Decode_INSTRUCTION_0 & 32'h00005004) == 32'h00001000),((toplevel_decode_ctrls_1_down_Decode_INSTRUCTION_0 & 32'h00002050) == 32'h00002000)}}}});
  assign _zz_toplevel_decode_ctrls_1_down_RS2_ENABLE_0 = (|{((toplevel_decode_ctrls_1_down_Decode_INSTRUCTION_0 & 32'h00000034) == 32'h00000020),{((toplevel_decode_ctrls_1_down_Decode_INSTRUCTION_0 & 32'h00000064) == 32'h00000020),{((toplevel_decode_ctrls_1_down_Decode_INSTRUCTION_0 & 32'h08000070) == 32'h08000020),((toplevel_decode_ctrls_1_down_Decode_INSTRUCTION_0 & 32'h10000070) == 32'h00000020)}}});
  assign _zz_toplevel_decode_ctrls_1_down_RD_ENABLE_0 = (|{_zz_toplevel_decode_ctrls_1_down_DispatchPlugin_logic_LANES_LAYER_HIT_3_0,{((toplevel_decode_ctrls_1_down_Decode_INSTRUCTION_0 & 32'h00001010) == 32'h00001010),{((toplevel_decode_ctrls_1_down_Decode_INSTRUCTION_0 & 32'h00002010) == 32'h00002010),{((toplevel_decode_ctrls_1_down_Decode_INSTRUCTION_0 & _zz_toplevel_decode_ctrls_1_down_RD_ENABLE_0_1) == 32'h00002008),{(_zz_toplevel_decode_ctrls_1_down_RD_ENABLE_0_2 == _zz_toplevel_decode_ctrls_1_down_RD_ENABLE_0_3),{_zz_toplevel_decode_ctrls_1_down_DispatchPlugin_logic_LANES_LAYER_HIT_0_0,_zz_toplevel_decode_ctrls_1_down_RD_ENABLE_0_4}}}}}});
  assign _zz_DecoderPlugin_logic_laneLogic_0_fixer_isJb = (|_zz_toplevel_decode_ctrls_1_down_DispatchPlugin_logic_LANES_LAYER_HIT_0_0_1);
  assign _zz_DecoderPlugin_logic_forgetPort_payload_pcOnLastSlice_1 = ((! toplevel_decode_ctrls_1_down_Prediction_ALIGN_REDO_0) ? _zz_DecoderPlugin_logic_forgetPort_payload_pcOnLastSlice_2 : 2'b00);
  assign _zz_DecoderPlugin_logic_forgetPort_payload_pcOnLastSlice = {30'd0, _zz_DecoderPlugin_logic_forgetPort_payload_pcOnLastSlice_1};
  assign _zz_DecoderPlugin_logic_forgetPort_payload_pcOnLastSlice_2 = ({1'd0,toplevel_decode_ctrls_1_down_Decode_INSTRUCTION_SLICE_COUNT_0} <<< 1'd1);
  assign _zz_toplevel_decode_ctrls_1_down_RS1_ENABLE_1 = (|{((toplevel_decode_ctrls_1_down_Decode_INSTRUCTION_1 & 32'h00000044) == 32'h0),{_zz_toplevel_decode_ctrls_1_down_DispatchPlugin_MAY_FLUSH_1,{((toplevel_decode_ctrls_1_down_Decode_INSTRUCTION_1 & 32'h00006004) == 32'h00002000),{((toplevel_decode_ctrls_1_down_Decode_INSTRUCTION_1 & 32'h00005004) == 32'h00001000),((toplevel_decode_ctrls_1_down_Decode_INSTRUCTION_1 & 32'h00002050) == 32'h00002000)}}}});
  assign _zz_toplevel_decode_ctrls_1_down_RS2_ENABLE_1 = (|{((toplevel_decode_ctrls_1_down_Decode_INSTRUCTION_1 & 32'h00000034) == 32'h00000020),{((toplevel_decode_ctrls_1_down_Decode_INSTRUCTION_1 & 32'h00000064) == 32'h00000020),{((toplevel_decode_ctrls_1_down_Decode_INSTRUCTION_1 & 32'h08000070) == 32'h08000020),((toplevel_decode_ctrls_1_down_Decode_INSTRUCTION_1 & 32'h10000070) == 32'h00000020)}}});
  assign _zz_toplevel_decode_ctrls_1_down_RD_ENABLE_1 = (|{_zz_toplevel_decode_ctrls_1_down_DispatchPlugin_logic_LANES_LAYER_HIT_3_1,{((toplevel_decode_ctrls_1_down_Decode_INSTRUCTION_1 & 32'h00001010) == 32'h00001010),{((toplevel_decode_ctrls_1_down_Decode_INSTRUCTION_1 & 32'h00002010) == 32'h00002010),{((toplevel_decode_ctrls_1_down_Decode_INSTRUCTION_1 & _zz_toplevel_decode_ctrls_1_down_RD_ENABLE_1_1) == 32'h00002008),{(_zz_toplevel_decode_ctrls_1_down_RD_ENABLE_1_2 == _zz_toplevel_decode_ctrls_1_down_RD_ENABLE_1_3),{_zz_toplevel_decode_ctrls_1_down_DispatchPlugin_logic_LANES_LAYER_HIT_0_1,_zz_toplevel_decode_ctrls_1_down_RD_ENABLE_1_4}}}}}});
  assign _zz_DecoderPlugin_logic_laneLogic_1_fixer_isJb = (|_zz_toplevel_decode_ctrls_1_down_DispatchPlugin_logic_LANES_LAYER_HIT_0_1_1);
  assign _zz_DecoderPlugin_logic_forgetPort_payload_pcOnLastSlice_4 = ((! toplevel_decode_ctrls_1_down_Prediction_ALIGN_REDO_1) ? _zz_DecoderPlugin_logic_forgetPort_payload_pcOnLastSlice_5 : 2'b00);
  assign _zz_DecoderPlugin_logic_forgetPort_payload_pcOnLastSlice_3 = {30'd0, _zz_DecoderPlugin_logic_forgetPort_payload_pcOnLastSlice_4};
  assign _zz_DecoderPlugin_logic_forgetPort_payload_pcOnLastSlice_5 = ({1'd0,toplevel_decode_ctrls_1_down_Decode_INSTRUCTION_SLICE_COUNT_1} <<< 1'd1);
  assign _zz_toplevel_decode_ctrls_1_down_DispatchPlugin_logic_LANES_LAYER_HIT_0_0_2 = _zz_toplevel_decode_ctrls_1_down_DispatchPlugin_logic_LANES_LAYER_HIT_0_0_3[0];
  assign _zz_toplevel_decode_ctrls_1_down_DispatchPlugin_logic_LANES_LAYER_HIT_0_0_3 = (|{_zz_toplevel_decode_ctrls_1_down_DispatchPlugin_logic_LANES_LAYER_HIT_3_0_2,{_zz_toplevel_decode_ctrls_1_down_DispatchPlugin_logic_LANES_LAYER_HIT_0_0_1,{_zz_toplevel_decode_ctrls_1_down_DispatchPlugin_logic_LANES_LAYER_HIT_0_0,_zz_toplevel_decode_ctrls_1_down_DispatchPlugin_logic_LANES_LAYER_HIT_3_0_1}}});
  assign _zz_toplevel_decode_ctrls_1_down_DispatchPlugin_logic_LANES_LAYER_HIT_1_0 = _zz_toplevel_decode_ctrls_1_down_DispatchPlugin_logic_LANES_LAYER_HIT_1_0_1[0];
  assign _zz_toplevel_decode_ctrls_1_down_DispatchPlugin_logic_LANES_LAYER_HIT_1_0_1 = (|_zz_toplevel_decode_ctrls_1_down_DispatchPlugin_logic_hcs_3_onRs_1_ENABLES_0_0);
  assign _zz_toplevel_decode_ctrls_1_down_DispatchPlugin_logic_LANES_LAYER_HIT_2_0 = _zz_toplevel_decode_ctrls_1_down_DispatchPlugin_logic_LANES_LAYER_HIT_2_0_1[0];
  assign _zz_toplevel_decode_ctrls_1_down_DispatchPlugin_logic_LANES_LAYER_HIT_2_0_1 = (|{_zz_toplevel_decode_ctrls_1_down_DispatchPlugin_logic_LANES_LAYER_HIT_3_0,{_zz_toplevel_decode_ctrls_1_down_DispatchPlugin_logic_LANES_LAYER_HIT_3_0_2,{_zz_toplevel_decode_ctrls_1_down_DispatchPlugin_logic_LANES_LAYER_HIT_3_0_4,{_zz_toplevel_decode_ctrls_1_down_DispatchPlugin_logic_LANES_LAYER_HIT_3_0_1,_zz_toplevel_decode_ctrls_1_down_DispatchPlugin_logic_LANES_LAYER_HIT_3_0_3}}}});
  assign _zz_toplevel_decode_ctrls_1_down_DispatchPlugin_logic_LANES_LAYER_HIT_3_0_5 = _zz_toplevel_decode_ctrls_1_down_DispatchPlugin_logic_LANES_LAYER_HIT_3_0_6[0];
  assign _zz_toplevel_decode_ctrls_1_down_DispatchPlugin_logic_LANES_LAYER_HIT_3_0_6 = (|{_zz_toplevel_decode_ctrls_1_down_DispatchPlugin_logic_LANES_LAYER_HIT_3_0,{_zz_toplevel_decode_ctrls_1_down_DispatchPlugin_logic_LANES_LAYER_HIT_3_0_2,{_zz_toplevel_decode_ctrls_1_down_DispatchPlugin_logic_LANES_LAYER_HIT_3_0_4,{_zz_toplevel_decode_ctrls_1_down_DispatchPlugin_logic_LANES_LAYER_HIT_3_0_1,_zz_toplevel_decode_ctrls_1_down_DispatchPlugin_logic_LANES_LAYER_HIT_3_0_3}}}});
  assign _zz_toplevel_decode_ctrls_1_down_DispatchPlugin_MAY_FLUSH_0_1 = _zz_toplevel_decode_ctrls_1_down_DispatchPlugin_MAY_FLUSH_0_2[0];
  assign _zz_toplevel_decode_ctrls_1_down_DispatchPlugin_MAY_FLUSH_0_2 = (|{_zz_toplevel_decode_ctrls_1_down_DispatchPlugin_logic_hcs_1_onRs_1_ENABLES_0_0,{((toplevel_decode_ctrls_1_down_Decode_INSTRUCTION_0 & 32'h00002010) == 32'h00002000),{((toplevel_decode_ctrls_1_down_Decode_INSTRUCTION_0 & 32'h00001010) == 32'h00001000),_zz_toplevel_decode_ctrls_1_down_DispatchPlugin_MAY_FLUSH_0}}});
  assign _zz_toplevel_decode_ctrls_1_down_DispatchPlugin_DONT_FLUSH_0 = _zz_toplevel_decode_ctrls_1_down_DispatchPlugin_DONT_FLUSH_0_1[0];
  assign _zz_toplevel_decode_ctrls_1_down_DispatchPlugin_DONT_FLUSH_0_1 = (|{_zz_toplevel_decode_ctrls_1_down_DONT_FLUSH_PRECISE_4_0_1,_zz_toplevel_decode_ctrls_1_down_DONT_FLUSH_PRECISE_4_0});
  assign _zz_toplevel_decode_ctrls_1_down_DispatchPlugin_DONT_FLUSH_FROM_LANES_0 = _zz_toplevel_decode_ctrls_1_down_DispatchPlugin_DONT_FLUSH_FROM_LANES_0_1[0];
  assign _zz_toplevel_decode_ctrls_1_down_DispatchPlugin_DONT_FLUSH_FROM_LANES_0_1 = (|{_zz_toplevel_decode_ctrls_1_down_DONT_FLUSH_PRECISE_4_0_1,_zz_toplevel_decode_ctrls_1_down_DONT_FLUSH_PRECISE_4_0});
  assign _zz_toplevel_decode_ctrls_1_down_DispatchPlugin_FENCE_OLDER_0 = _zz_toplevel_decode_ctrls_1_down_DispatchPlugin_FENCE_OLDER_0_1[0];
  assign _zz_toplevel_decode_ctrls_1_down_DispatchPlugin_FENCE_OLDER_0_1 = (|{_zz_toplevel_decode_ctrls_1_down_DONT_FLUSH_PRECISE_4_0_1,_zz_toplevel_decode_ctrls_1_down_DONT_FLUSH_PRECISE_4_0});
  assign _zz_toplevel_decode_ctrls_1_down_DONT_FLUSH_PRECISE_3_0 = _zz_toplevel_decode_ctrls_1_down_DONT_FLUSH_PRECISE_3_0_1[0];
  assign _zz_toplevel_decode_ctrls_1_down_DONT_FLUSH_PRECISE_3_0_1 = (|{_zz_toplevel_decode_ctrls_1_down_DONT_FLUSH_PRECISE_4_0_1,_zz_toplevel_decode_ctrls_1_down_DONT_FLUSH_PRECISE_4_0});
  assign _zz_toplevel_decode_ctrls_1_down_DONT_FLUSH_PRECISE_4_0_2 = _zz_toplevel_decode_ctrls_1_down_DONT_FLUSH_PRECISE_4_0_3[0];
  assign _zz_toplevel_decode_ctrls_1_down_DONT_FLUSH_PRECISE_4_0_3 = (|{_zz_toplevel_decode_ctrls_1_down_DONT_FLUSH_PRECISE_4_0_1,_zz_toplevel_decode_ctrls_1_down_DONT_FLUSH_PRECISE_4_0});
  assign _zz_toplevel_decode_ctrls_1_down_DecoderPlugin_logic_NEED_FPU_0 = _zz_toplevel_decode_ctrls_1_down_DecoderPlugin_logic_NEED_FPU_0_1[0];
  assign _zz_toplevel_decode_ctrls_1_down_DecoderPlugin_logic_NEED_FPU_0_1 = 1'b0;
  assign _zz_toplevel_decode_ctrls_1_down_DecoderPlugin_logic_NEED_RM_0 = _zz_toplevel_decode_ctrls_1_down_DecoderPlugin_logic_NEED_RM_0_1[0];
  assign _zz_toplevel_decode_ctrls_1_down_DecoderPlugin_logic_NEED_RM_0_1 = 1'b0;
  assign _zz_toplevel_decode_ctrls_1_down_DispatchPlugin_logic_hcs_0_onRs_0_ENABLES_0_0 = _zz_toplevel_decode_ctrls_1_down_DispatchPlugin_logic_hcs_0_onRs_0_ENABLES_0_0_1[0];
  assign _zz_toplevel_decode_ctrls_1_down_DispatchPlugin_logic_hcs_0_onRs_0_ENABLES_0_0_1 = (|_zz_toplevel_decode_ctrls_1_down_DispatchPlugin_logic_hcs_3_onRs_1_ENABLES_0_0);
  assign _zz_toplevel_decode_ctrls_1_down_DispatchPlugin_logic_hcs_0_onRs_1_ENABLES_0_0 = _zz_toplevel_decode_ctrls_1_down_DispatchPlugin_logic_hcs_0_onRs_1_ENABLES_0_0_1[0];
  assign _zz_toplevel_decode_ctrls_1_down_DispatchPlugin_logic_hcs_0_onRs_1_ENABLES_0_0_1 = (|_zz_toplevel_decode_ctrls_1_down_DispatchPlugin_logic_hcs_3_onRs_1_ENABLES_0_0);
  assign _zz_toplevel_decode_ctrls_1_down_DispatchPlugin_logic_hcs_1_onRs_0_ENABLES_0_0 = _zz_toplevel_decode_ctrls_1_down_DispatchPlugin_logic_hcs_1_onRs_0_ENABLES_0_0_1[0];
  assign _zz_toplevel_decode_ctrls_1_down_DispatchPlugin_logic_hcs_1_onRs_0_ENABLES_0_0_1 = (|_zz_toplevel_decode_ctrls_1_down_DispatchPlugin_logic_hcs_3_onRs_1_ENABLES_0_0);
  assign _zz_toplevel_decode_ctrls_1_down_DispatchPlugin_logic_hcs_1_onRs_1_ENABLES_0_0_1 = _zz_toplevel_decode_ctrls_1_down_DispatchPlugin_logic_hcs_1_onRs_1_ENABLES_0_0_2[0];
  assign _zz_toplevel_decode_ctrls_1_down_DispatchPlugin_logic_hcs_1_onRs_1_ENABLES_0_0_2 = (|{_zz_toplevel_decode_ctrls_1_down_DispatchPlugin_logic_hcs_1_onRs_1_ENABLES_0_0,((toplevel_decode_ctrls_1_down_Decode_INSTRUCTION_0 & 32'h00000010) == 32'h00000010)});
  assign _zz_toplevel_decode_ctrls_1_down_DispatchPlugin_logic_hcs_1_onRs_1_ENABLES_1_0 = _zz_toplevel_decode_ctrls_1_down_DispatchPlugin_logic_hcs_1_onRs_1_ENABLES_1_0_1[0];
  assign _zz_toplevel_decode_ctrls_1_down_DispatchPlugin_logic_hcs_1_onRs_1_ENABLES_1_0_1 = (|_zz_toplevel_decode_ctrls_1_down_DispatchPlugin_logic_hcs_3_onRs_1_ENABLES_0_0);
  assign _zz_toplevel_decode_ctrls_1_down_DispatchPlugin_logic_hcs_2_onRs_0_ENABLES_0_0 = _zz_toplevel_decode_ctrls_1_down_DispatchPlugin_logic_hcs_2_onRs_0_ENABLES_0_0_1[0];
  assign _zz_toplevel_decode_ctrls_1_down_DispatchPlugin_logic_hcs_2_onRs_0_ENABLES_0_0_1 = (|_zz_toplevel_decode_ctrls_1_down_DispatchPlugin_logic_hcs_3_onRs_1_ENABLES_0_0);
  assign _zz_toplevel_decode_ctrls_1_down_DispatchPlugin_logic_hcs_2_onRs_1_ENABLES_0_0 = _zz_toplevel_decode_ctrls_1_down_DispatchPlugin_logic_hcs_2_onRs_1_ENABLES_0_0_1[0];
  assign _zz_toplevel_decode_ctrls_1_down_DispatchPlugin_logic_hcs_2_onRs_1_ENABLES_0_0_1 = (|_zz_toplevel_decode_ctrls_1_down_DispatchPlugin_logic_hcs_3_onRs_1_ENABLES_0_0);
  assign _zz_toplevel_decode_ctrls_1_down_DispatchPlugin_logic_hcs_3_onRs_0_ENABLES_0_0 = _zz_toplevel_decode_ctrls_1_down_DispatchPlugin_logic_hcs_3_onRs_0_ENABLES_0_0_1[0];
  assign _zz_toplevel_decode_ctrls_1_down_DispatchPlugin_logic_hcs_3_onRs_0_ENABLES_0_0_1 = (|_zz_toplevel_decode_ctrls_1_down_DispatchPlugin_logic_hcs_3_onRs_1_ENABLES_0_0);
  assign _zz_toplevel_decode_ctrls_1_down_DispatchPlugin_logic_hcs_3_onRs_1_ENABLES_0_0_1 = _zz_toplevel_decode_ctrls_1_down_DispatchPlugin_logic_hcs_3_onRs_1_ENABLES_0_0_2[0];
  assign _zz_toplevel_decode_ctrls_1_down_DispatchPlugin_logic_hcs_3_onRs_1_ENABLES_0_0_2 = (|_zz_toplevel_decode_ctrls_1_down_DispatchPlugin_logic_hcs_3_onRs_1_ENABLES_0_0);
  assign _zz_toplevel_decode_ctrls_1_down_DispatchPlugin_logic_LANES_LAYER_HIT_0_1_2 = _zz_toplevel_decode_ctrls_1_down_DispatchPlugin_logic_LANES_LAYER_HIT_0_1_3[0];
  assign _zz_toplevel_decode_ctrls_1_down_DispatchPlugin_logic_LANES_LAYER_HIT_0_1_3 = (|{_zz_toplevel_decode_ctrls_1_down_DispatchPlugin_logic_LANES_LAYER_HIT_3_1_2,{_zz_toplevel_decode_ctrls_1_down_DispatchPlugin_logic_LANES_LAYER_HIT_0_1_1,{_zz_toplevel_decode_ctrls_1_down_DispatchPlugin_logic_LANES_LAYER_HIT_0_1,_zz_toplevel_decode_ctrls_1_down_DispatchPlugin_logic_LANES_LAYER_HIT_3_1_1}}});
  assign _zz_toplevel_decode_ctrls_1_down_DispatchPlugin_logic_LANES_LAYER_HIT_1_1 = _zz_toplevel_decode_ctrls_1_down_DispatchPlugin_logic_LANES_LAYER_HIT_1_1_1[0];
  assign _zz_toplevel_decode_ctrls_1_down_DispatchPlugin_logic_LANES_LAYER_HIT_1_1_1 = (|_zz_toplevel_decode_ctrls_1_down_DispatchPlugin_logic_hcs_3_onRs_1_ENABLES_0_1);
  assign _zz_toplevel_decode_ctrls_1_down_DispatchPlugin_logic_LANES_LAYER_HIT_2_1 = _zz_toplevel_decode_ctrls_1_down_DispatchPlugin_logic_LANES_LAYER_HIT_2_1_1[0];
  assign _zz_toplevel_decode_ctrls_1_down_DispatchPlugin_logic_LANES_LAYER_HIT_2_1_1 = (|{_zz_toplevel_decode_ctrls_1_down_DispatchPlugin_logic_LANES_LAYER_HIT_3_1,{_zz_toplevel_decode_ctrls_1_down_DispatchPlugin_logic_LANES_LAYER_HIT_3_1_2,{_zz_toplevel_decode_ctrls_1_down_DispatchPlugin_logic_LANES_LAYER_HIT_3_1_4,{_zz_toplevel_decode_ctrls_1_down_DispatchPlugin_logic_LANES_LAYER_HIT_3_1_1,_zz_toplevel_decode_ctrls_1_down_DispatchPlugin_logic_LANES_LAYER_HIT_3_1_3}}}});
  assign _zz_toplevel_decode_ctrls_1_down_DispatchPlugin_logic_LANES_LAYER_HIT_3_1_5 = _zz_toplevel_decode_ctrls_1_down_DispatchPlugin_logic_LANES_LAYER_HIT_3_1_6[0];
  assign _zz_toplevel_decode_ctrls_1_down_DispatchPlugin_logic_LANES_LAYER_HIT_3_1_6 = (|{_zz_toplevel_decode_ctrls_1_down_DispatchPlugin_logic_LANES_LAYER_HIT_3_1,{_zz_toplevel_decode_ctrls_1_down_DispatchPlugin_logic_LANES_LAYER_HIT_3_1_2,{_zz_toplevel_decode_ctrls_1_down_DispatchPlugin_logic_LANES_LAYER_HIT_3_1_4,{_zz_toplevel_decode_ctrls_1_down_DispatchPlugin_logic_LANES_LAYER_HIT_3_1_1,_zz_toplevel_decode_ctrls_1_down_DispatchPlugin_logic_LANES_LAYER_HIT_3_1_3}}}});
  assign _zz_toplevel_decode_ctrls_1_down_DispatchPlugin_MAY_FLUSH_1_1 = _zz_toplevel_decode_ctrls_1_down_DispatchPlugin_MAY_FLUSH_1_2[0];
  assign _zz_toplevel_decode_ctrls_1_down_DispatchPlugin_MAY_FLUSH_1_2 = (|{_zz_toplevel_decode_ctrls_1_down_DispatchPlugin_logic_hcs_1_onRs_1_ENABLES_0_1,{((toplevel_decode_ctrls_1_down_Decode_INSTRUCTION_1 & 32'h00002010) == 32'h00002000),{((toplevel_decode_ctrls_1_down_Decode_INSTRUCTION_1 & 32'h00001010) == 32'h00001000),_zz_toplevel_decode_ctrls_1_down_DispatchPlugin_MAY_FLUSH_1}}});
  assign _zz_toplevel_decode_ctrls_1_down_DispatchPlugin_DONT_FLUSH_1 = _zz_toplevel_decode_ctrls_1_down_DispatchPlugin_DONT_FLUSH_1_1[0];
  assign _zz_toplevel_decode_ctrls_1_down_DispatchPlugin_DONT_FLUSH_1_1 = (|{_zz_toplevel_decode_ctrls_1_down_DONT_FLUSH_PRECISE_4_1_1,_zz_toplevel_decode_ctrls_1_down_DONT_FLUSH_PRECISE_4_1});
  assign _zz_toplevel_decode_ctrls_1_down_DispatchPlugin_DONT_FLUSH_FROM_LANES_1 = _zz_toplevel_decode_ctrls_1_down_DispatchPlugin_DONT_FLUSH_FROM_LANES_1_1[0];
  assign _zz_toplevel_decode_ctrls_1_down_DispatchPlugin_DONT_FLUSH_FROM_LANES_1_1 = (|{_zz_toplevel_decode_ctrls_1_down_DONT_FLUSH_PRECISE_4_1_1,_zz_toplevel_decode_ctrls_1_down_DONT_FLUSH_PRECISE_4_1});
  assign _zz_toplevel_decode_ctrls_1_down_DispatchPlugin_FENCE_OLDER_1 = _zz_toplevel_decode_ctrls_1_down_DispatchPlugin_FENCE_OLDER_1_1[0];
  assign _zz_toplevel_decode_ctrls_1_down_DispatchPlugin_FENCE_OLDER_1_1 = (|{_zz_toplevel_decode_ctrls_1_down_DONT_FLUSH_PRECISE_4_1_1,_zz_toplevel_decode_ctrls_1_down_DONT_FLUSH_PRECISE_4_1});
  assign _zz_toplevel_decode_ctrls_1_down_DONT_FLUSH_PRECISE_3_1 = _zz_toplevel_decode_ctrls_1_down_DONT_FLUSH_PRECISE_3_1_1[0];
  assign _zz_toplevel_decode_ctrls_1_down_DONT_FLUSH_PRECISE_3_1_1 = (|{_zz_toplevel_decode_ctrls_1_down_DONT_FLUSH_PRECISE_4_1_1,_zz_toplevel_decode_ctrls_1_down_DONT_FLUSH_PRECISE_4_1});
  assign _zz_toplevel_decode_ctrls_1_down_DONT_FLUSH_PRECISE_4_1_2 = _zz_toplevel_decode_ctrls_1_down_DONT_FLUSH_PRECISE_4_1_3[0];
  assign _zz_toplevel_decode_ctrls_1_down_DONT_FLUSH_PRECISE_4_1_3 = (|{_zz_toplevel_decode_ctrls_1_down_DONT_FLUSH_PRECISE_4_1_1,_zz_toplevel_decode_ctrls_1_down_DONT_FLUSH_PRECISE_4_1});
  assign _zz_toplevel_decode_ctrls_1_down_DecoderPlugin_logic_NEED_FPU_1 = _zz_toplevel_decode_ctrls_1_down_DecoderPlugin_logic_NEED_FPU_1_1[0];
  assign _zz_toplevel_decode_ctrls_1_down_DecoderPlugin_logic_NEED_FPU_1_1 = 1'b0;
  assign _zz_toplevel_decode_ctrls_1_down_DecoderPlugin_logic_NEED_RM_1 = _zz_toplevel_decode_ctrls_1_down_DecoderPlugin_logic_NEED_RM_1_1[0];
  assign _zz_toplevel_decode_ctrls_1_down_DecoderPlugin_logic_NEED_RM_1_1 = 1'b0;
  assign _zz_toplevel_decode_ctrls_1_down_DispatchPlugin_logic_hcs_0_onRs_0_ENABLES_0_1 = _zz_toplevel_decode_ctrls_1_down_DispatchPlugin_logic_hcs_0_onRs_0_ENABLES_0_1_1[0];
  assign _zz_toplevel_decode_ctrls_1_down_DispatchPlugin_logic_hcs_0_onRs_0_ENABLES_0_1_1 = (|_zz_toplevel_decode_ctrls_1_down_DispatchPlugin_logic_hcs_3_onRs_1_ENABLES_0_1);
  assign _zz_toplevel_decode_ctrls_1_down_DispatchPlugin_logic_hcs_0_onRs_1_ENABLES_0_1 = _zz_toplevel_decode_ctrls_1_down_DispatchPlugin_logic_hcs_0_onRs_1_ENABLES_0_1_1[0];
  assign _zz_toplevel_decode_ctrls_1_down_DispatchPlugin_logic_hcs_0_onRs_1_ENABLES_0_1_1 = (|_zz_toplevel_decode_ctrls_1_down_DispatchPlugin_logic_hcs_3_onRs_1_ENABLES_0_1);
  assign _zz_toplevel_decode_ctrls_1_down_DispatchPlugin_logic_hcs_1_onRs_0_ENABLES_0_1 = _zz_toplevel_decode_ctrls_1_down_DispatchPlugin_logic_hcs_1_onRs_0_ENABLES_0_1_1[0];
  assign _zz_toplevel_decode_ctrls_1_down_DispatchPlugin_logic_hcs_1_onRs_0_ENABLES_0_1_1 = (|_zz_toplevel_decode_ctrls_1_down_DispatchPlugin_logic_hcs_3_onRs_1_ENABLES_0_1);
  assign _zz_toplevel_decode_ctrls_1_down_DispatchPlugin_logic_hcs_1_onRs_1_ENABLES_0_1_1 = _zz_toplevel_decode_ctrls_1_down_DispatchPlugin_logic_hcs_1_onRs_1_ENABLES_0_1_2[0];
  assign _zz_toplevel_decode_ctrls_1_down_DispatchPlugin_logic_hcs_1_onRs_1_ENABLES_0_1_2 = (|{_zz_toplevel_decode_ctrls_1_down_DispatchPlugin_logic_hcs_1_onRs_1_ENABLES_0_1,((toplevel_decode_ctrls_1_down_Decode_INSTRUCTION_1 & 32'h00000010) == 32'h00000010)});
  assign _zz_toplevel_decode_ctrls_1_down_DispatchPlugin_logic_hcs_1_onRs_1_ENABLES_1_1 = _zz_toplevel_decode_ctrls_1_down_DispatchPlugin_logic_hcs_1_onRs_1_ENABLES_1_1_1[0];
  assign _zz_toplevel_decode_ctrls_1_down_DispatchPlugin_logic_hcs_1_onRs_1_ENABLES_1_1_1 = (|_zz_toplevel_decode_ctrls_1_down_DispatchPlugin_logic_hcs_3_onRs_1_ENABLES_0_1);
  assign _zz_toplevel_decode_ctrls_1_down_DispatchPlugin_logic_hcs_2_onRs_0_ENABLES_0_1 = _zz_toplevel_decode_ctrls_1_down_DispatchPlugin_logic_hcs_2_onRs_0_ENABLES_0_1_1[0];
  assign _zz_toplevel_decode_ctrls_1_down_DispatchPlugin_logic_hcs_2_onRs_0_ENABLES_0_1_1 = (|_zz_toplevel_decode_ctrls_1_down_DispatchPlugin_logic_hcs_3_onRs_1_ENABLES_0_1);
  assign _zz_toplevel_decode_ctrls_1_down_DispatchPlugin_logic_hcs_2_onRs_1_ENABLES_0_1 = _zz_toplevel_decode_ctrls_1_down_DispatchPlugin_logic_hcs_2_onRs_1_ENABLES_0_1_1[0];
  assign _zz_toplevel_decode_ctrls_1_down_DispatchPlugin_logic_hcs_2_onRs_1_ENABLES_0_1_1 = (|_zz_toplevel_decode_ctrls_1_down_DispatchPlugin_logic_hcs_3_onRs_1_ENABLES_0_1);
  assign _zz_toplevel_decode_ctrls_1_down_DispatchPlugin_logic_hcs_3_onRs_0_ENABLES_0_1 = _zz_toplevel_decode_ctrls_1_down_DispatchPlugin_logic_hcs_3_onRs_0_ENABLES_0_1_1[0];
  assign _zz_toplevel_decode_ctrls_1_down_DispatchPlugin_logic_hcs_3_onRs_0_ENABLES_0_1_1 = (|_zz_toplevel_decode_ctrls_1_down_DispatchPlugin_logic_hcs_3_onRs_1_ENABLES_0_1);
  assign _zz_toplevel_decode_ctrls_1_down_DispatchPlugin_logic_hcs_3_onRs_1_ENABLES_0_1_1 = _zz_toplevel_decode_ctrls_1_down_DispatchPlugin_logic_hcs_3_onRs_1_ENABLES_0_1_2[0];
  assign _zz_toplevel_decode_ctrls_1_down_DispatchPlugin_logic_hcs_3_onRs_1_ENABLES_0_1_2 = (|_zz_toplevel_decode_ctrls_1_down_DispatchPlugin_logic_hcs_3_onRs_1_ENABLES_0_1);
  assign _zz_BtbPlugin_logic_onLearn_port_payload_address_1 = (DecoderPlugin_logic_forgetPort_payload_pcOnLastSlice >>> 2'd3);
  assign _zz_BtbPlugin_logic_readPort_cmd_payload = (fetch_logic_ctrls_0_down_Fetch_WORD_PC >>> 2'd3);
  assign _zz_BtbPlugin_logic_ras_write_payload_data = (BtbPlugin_logic_applyIt_rasLogic_pushPc + 32'h00000002);
  assign _zz_DispatchPlugin_logic_inserter_0_trap = (((_zz_toplevel_execute_ctrl0_up_LANE_AGE_lane0 ? DispatchPlugin_logic_candidates_0_ctx_hm_TRAP : 1'b0) | (_zz_toplevel_execute_ctrl0_up_LANE_AGE_lane0_1 ? DispatchPlugin_logic_candidates_1_ctx_hm_TRAP : 1'b0)) | (_zz_toplevel_execute_ctrl0_up_LANE_AGE_lane0_2 ? DispatchPlugin_logic_candidates_2_ctx_hm_TRAP : 1'b0));
  assign _zz_toplevel_execute_ctrl0_up_LANE_SEL_lane0 = (((_zz_toplevel_execute_ctrl0_up_LANE_AGE_lane0 ? DispatchPlugin_logic_candidates_0_cancel : 1'b0) | (_zz_toplevel_execute_ctrl0_up_LANE_AGE_lane0_1 ? DispatchPlugin_logic_candidates_1_cancel : 1'b0)) | (_zz_toplevel_execute_ctrl0_up_LANE_AGE_lane0_2 ? DispatchPlugin_logic_candidates_2_cancel : 1'b0));
  assign _zz_toplevel_execute_ctrl0_up_Prediction_ALIGNED_JUMPED_lane0 = (((_zz_toplevel_execute_ctrl0_up_LANE_AGE_lane0 ? DispatchPlugin_logic_candidates_0_ctx_hm_Prediction_ALIGNED_JUMPED : 1'b0) | (_zz_toplevel_execute_ctrl0_up_LANE_AGE_lane0_1 ? DispatchPlugin_logic_candidates_1_ctx_hm_Prediction_ALIGNED_JUMPED : 1'b0)) | (_zz_toplevel_execute_ctrl0_up_LANE_AGE_lane0_2 ? DispatchPlugin_logic_candidates_2_ctx_hm_Prediction_ALIGNED_JUMPED : 1'b0));
  assign _zz_toplevel_execute_ctrl0_up_DispatchPlugin_FENCE_OLDER_lane0 = (((_zz_toplevel_execute_ctrl0_up_LANE_AGE_lane0 ? DispatchPlugin_logic_candidates_0_ctx_hm_DispatchPlugin_FENCE_OLDER : 1'b0) | (_zz_toplevel_execute_ctrl0_up_LANE_AGE_lane0_1 ? DispatchPlugin_logic_candidates_1_ctx_hm_DispatchPlugin_FENCE_OLDER : 1'b0)) | (_zz_toplevel_execute_ctrl0_up_LANE_AGE_lane0_2 ? DispatchPlugin_logic_candidates_2_ctx_hm_DispatchPlugin_FENCE_OLDER : 1'b0));
  assign _zz_toplevel_execute_ctrl0_up_DispatchPlugin_MAY_FLUSH_lane0 = (((_zz_toplevel_execute_ctrl0_up_LANE_AGE_lane0 ? DispatchPlugin_logic_candidates_0_ctx_hm_DispatchPlugin_MAY_FLUSH : 1'b0) | (_zz_toplevel_execute_ctrl0_up_LANE_AGE_lane0_1 ? DispatchPlugin_logic_candidates_1_ctx_hm_DispatchPlugin_MAY_FLUSH : 1'b0)) | (_zz_toplevel_execute_ctrl0_up_LANE_AGE_lane0_2 ? DispatchPlugin_logic_candidates_2_ctx_hm_DispatchPlugin_MAY_FLUSH : 1'b0));
  assign _zz_toplevel_execute_ctrl0_up_DispatchPlugin_DONT_FLUSH_lane0 = (((_zz_toplevel_execute_ctrl0_up_LANE_AGE_lane0 ? DispatchPlugin_logic_candidates_0_ctx_hm_DispatchPlugin_DONT_FLUSH : 1'b0) | (_zz_toplevel_execute_ctrl0_up_LANE_AGE_lane0_1 ? DispatchPlugin_logic_candidates_1_ctx_hm_DispatchPlugin_DONT_FLUSH : 1'b0)) | (_zz_toplevel_execute_ctrl0_up_LANE_AGE_lane0_2 ? DispatchPlugin_logic_candidates_2_ctx_hm_DispatchPlugin_DONT_FLUSH : 1'b0));
  assign _zz_toplevel_execute_ctrl0_up_DispatchPlugin_DONT_FLUSH_FROM_LANES_lane0 = (((_zz_toplevel_execute_ctrl0_up_LANE_AGE_lane0 ? DispatchPlugin_logic_candidates_0_ctx_hm_DispatchPlugin_DONT_FLUSH_FROM_LANES : 1'b0) | (_zz_toplevel_execute_ctrl0_up_LANE_AGE_lane0_1 ? DispatchPlugin_logic_candidates_1_ctx_hm_DispatchPlugin_DONT_FLUSH_FROM_LANES : 1'b0)) | (_zz_toplevel_execute_ctrl0_up_LANE_AGE_lane0_2 ? DispatchPlugin_logic_candidates_2_ctx_hm_DispatchPlugin_DONT_FLUSH_FROM_LANES : 1'b0));
  assign _zz_toplevel_execute_ctrl0_up_DONT_FLUSH_PRECISE_3_lane0 = (((_zz_toplevel_execute_ctrl0_up_LANE_AGE_lane0 ? DispatchPlugin_logic_candidates_0_ctx_hm_DONT_FLUSH_PRECISE_3 : 1'b0) | (_zz_toplevel_execute_ctrl0_up_LANE_AGE_lane0_1 ? DispatchPlugin_logic_candidates_1_ctx_hm_DONT_FLUSH_PRECISE_3 : 1'b0)) | (_zz_toplevel_execute_ctrl0_up_LANE_AGE_lane0_2 ? DispatchPlugin_logic_candidates_2_ctx_hm_DONT_FLUSH_PRECISE_3 : 1'b0));
  assign _zz_toplevel_execute_ctrl0_up_DONT_FLUSH_PRECISE_4_lane0 = (((_zz_toplevel_execute_ctrl0_up_LANE_AGE_lane0 ? DispatchPlugin_logic_candidates_0_ctx_hm_DONT_FLUSH_PRECISE_4 : 1'b0) | (_zz_toplevel_execute_ctrl0_up_LANE_AGE_lane0_1 ? DispatchPlugin_logic_candidates_1_ctx_hm_DONT_FLUSH_PRECISE_4 : 1'b0)) | (_zz_toplevel_execute_ctrl0_up_LANE_AGE_lane0_2 ? DispatchPlugin_logic_candidates_2_ctx_hm_DONT_FLUSH_PRECISE_4 : 1'b0));
  assign _zz_toplevel_execute_ctrl0_up_TRAP_lane0 = (((_zz_toplevel_execute_ctrl0_up_LANE_AGE_lane0 ? DispatchPlugin_logic_candidates_0_ctx_hm_TRAP : 1'b0) | (_zz_toplevel_execute_ctrl0_up_LANE_AGE_lane0_1 ? DispatchPlugin_logic_candidates_1_ctx_hm_TRAP : 1'b0)) | (_zz_toplevel_execute_ctrl0_up_LANE_AGE_lane0_2 ? DispatchPlugin_logic_candidates_2_ctx_hm_TRAP : 1'b0));
  assign _zz_toplevel_execute_ctrl0_up_RS1_ENABLE_lane0 = (((_zz_toplevel_execute_ctrl0_up_LANE_AGE_lane0 ? DispatchPlugin_logic_candidates_0_ctx_hm_RS1_ENABLE : 1'b0) | (_zz_toplevel_execute_ctrl0_up_LANE_AGE_lane0_1 ? DispatchPlugin_logic_candidates_1_ctx_hm_RS1_ENABLE : 1'b0)) | (_zz_toplevel_execute_ctrl0_up_LANE_AGE_lane0_2 ? DispatchPlugin_logic_candidates_2_ctx_hm_RS1_ENABLE : 1'b0));
  assign _zz_toplevel_execute_ctrl0_up_RS2_ENABLE_lane0 = (((_zz_toplevel_execute_ctrl0_up_LANE_AGE_lane0 ? DispatchPlugin_logic_candidates_0_ctx_hm_RS2_ENABLE : 1'b0) | (_zz_toplevel_execute_ctrl0_up_LANE_AGE_lane0_1 ? DispatchPlugin_logic_candidates_1_ctx_hm_RS2_ENABLE : 1'b0)) | (_zz_toplevel_execute_ctrl0_up_LANE_AGE_lane0_2 ? DispatchPlugin_logic_candidates_2_ctx_hm_RS2_ENABLE : 1'b0));
  assign _zz_toplevel_execute_ctrl0_up_RD_ENABLE_lane0 = (((_zz_toplevel_execute_ctrl0_up_LANE_AGE_lane0 ? DispatchPlugin_logic_candidates_0_ctx_hm_RD_ENABLE : 1'b0) | (_zz_toplevel_execute_ctrl0_up_LANE_AGE_lane0_1 ? DispatchPlugin_logic_candidates_1_ctx_hm_RD_ENABLE : 1'b0)) | (_zz_toplevel_execute_ctrl0_up_LANE_AGE_lane0_2 ? DispatchPlugin_logic_candidates_2_ctx_hm_RD_ENABLE : 1'b0));
  assign _zz_toplevel_execute_ctrl0_up_DispatchPlugin_logic_hcs_0_onRs_0_ENABLES_0_lane0 = (((_zz_toplevel_execute_ctrl0_up_LANE_AGE_lane0 ? DispatchPlugin_logic_candidates_0_ctx_hm_DispatchPlugin_logic_hcs_0_onRs_0_ENABLES_0 : 1'b0) | (_zz_toplevel_execute_ctrl0_up_LANE_AGE_lane0_1 ? DispatchPlugin_logic_candidates_1_ctx_hm_DispatchPlugin_logic_hcs_0_onRs_0_ENABLES_0 : 1'b0)) | (_zz_toplevel_execute_ctrl0_up_LANE_AGE_lane0_2 ? DispatchPlugin_logic_candidates_2_ctx_hm_DispatchPlugin_logic_hcs_0_onRs_0_ENABLES_0 : 1'b0));
  assign _zz_toplevel_execute_ctrl0_up_DispatchPlugin_logic_hcs_0_onRs_1_ENABLES_0_lane0 = (((_zz_toplevel_execute_ctrl0_up_LANE_AGE_lane0 ? DispatchPlugin_logic_candidates_0_ctx_hm_DispatchPlugin_logic_hcs_0_onRs_1_ENABLES_0 : 1'b0) | (_zz_toplevel_execute_ctrl0_up_LANE_AGE_lane0_1 ? DispatchPlugin_logic_candidates_1_ctx_hm_DispatchPlugin_logic_hcs_0_onRs_1_ENABLES_0 : 1'b0)) | (_zz_toplevel_execute_ctrl0_up_LANE_AGE_lane0_2 ? DispatchPlugin_logic_candidates_2_ctx_hm_DispatchPlugin_logic_hcs_0_onRs_1_ENABLES_0 : 1'b0));
  assign _zz_toplevel_execute_ctrl0_up_DispatchPlugin_logic_hcs_1_onRs_0_ENABLES_0_lane0 = (((_zz_toplevel_execute_ctrl0_up_LANE_AGE_lane0 ? DispatchPlugin_logic_candidates_0_ctx_hm_DispatchPlugin_logic_hcs_1_onRs_0_ENABLES_0 : 1'b0) | (_zz_toplevel_execute_ctrl0_up_LANE_AGE_lane0_1 ? DispatchPlugin_logic_candidates_1_ctx_hm_DispatchPlugin_logic_hcs_1_onRs_0_ENABLES_0 : 1'b0)) | (_zz_toplevel_execute_ctrl0_up_LANE_AGE_lane0_2 ? DispatchPlugin_logic_candidates_2_ctx_hm_DispatchPlugin_logic_hcs_1_onRs_0_ENABLES_0 : 1'b0));
  assign _zz_toplevel_execute_ctrl0_up_DispatchPlugin_logic_hcs_1_onRs_1_ENABLES_0_lane0 = (((_zz_toplevel_execute_ctrl0_up_LANE_AGE_lane0 ? DispatchPlugin_logic_candidates_0_ctx_hm_DispatchPlugin_logic_hcs_1_onRs_1_ENABLES_0 : 1'b0) | (_zz_toplevel_execute_ctrl0_up_LANE_AGE_lane0_1 ? DispatchPlugin_logic_candidates_1_ctx_hm_DispatchPlugin_logic_hcs_1_onRs_1_ENABLES_0 : 1'b0)) | (_zz_toplevel_execute_ctrl0_up_LANE_AGE_lane0_2 ? DispatchPlugin_logic_candidates_2_ctx_hm_DispatchPlugin_logic_hcs_1_onRs_1_ENABLES_0 : 1'b0));
  assign _zz_toplevel_execute_ctrl0_up_DispatchPlugin_logic_hcs_1_onRs_1_ENABLES_1_lane0 = (((_zz_toplevel_execute_ctrl0_up_LANE_AGE_lane0 ? DispatchPlugin_logic_candidates_0_ctx_hm_DispatchPlugin_logic_hcs_1_onRs_1_ENABLES_1 : 1'b0) | (_zz_toplevel_execute_ctrl0_up_LANE_AGE_lane0_1 ? DispatchPlugin_logic_candidates_1_ctx_hm_DispatchPlugin_logic_hcs_1_onRs_1_ENABLES_1 : 1'b0)) | (_zz_toplevel_execute_ctrl0_up_LANE_AGE_lane0_2 ? DispatchPlugin_logic_candidates_2_ctx_hm_DispatchPlugin_logic_hcs_1_onRs_1_ENABLES_1 : 1'b0));
  assign _zz_toplevel_execute_ctrl0_up_DispatchPlugin_logic_hcs_2_onRs_0_ENABLES_0_lane0 = (((_zz_toplevel_execute_ctrl0_up_LANE_AGE_lane0 ? DispatchPlugin_logic_candidates_0_ctx_hm_DispatchPlugin_logic_hcs_2_onRs_0_ENABLES_0 : 1'b0) | (_zz_toplevel_execute_ctrl0_up_LANE_AGE_lane0_1 ? DispatchPlugin_logic_candidates_1_ctx_hm_DispatchPlugin_logic_hcs_2_onRs_0_ENABLES_0 : 1'b0)) | (_zz_toplevel_execute_ctrl0_up_LANE_AGE_lane0_2 ? DispatchPlugin_logic_candidates_2_ctx_hm_DispatchPlugin_logic_hcs_2_onRs_0_ENABLES_0 : 1'b0));
  assign _zz_toplevel_execute_ctrl0_up_DispatchPlugin_logic_hcs_2_onRs_1_ENABLES_0_lane0 = (((_zz_toplevel_execute_ctrl0_up_LANE_AGE_lane0 ? DispatchPlugin_logic_candidates_0_ctx_hm_DispatchPlugin_logic_hcs_2_onRs_1_ENABLES_0 : 1'b0) | (_zz_toplevel_execute_ctrl0_up_LANE_AGE_lane0_1 ? DispatchPlugin_logic_candidates_1_ctx_hm_DispatchPlugin_logic_hcs_2_onRs_1_ENABLES_0 : 1'b0)) | (_zz_toplevel_execute_ctrl0_up_LANE_AGE_lane0_2 ? DispatchPlugin_logic_candidates_2_ctx_hm_DispatchPlugin_logic_hcs_2_onRs_1_ENABLES_0 : 1'b0));
  assign _zz_toplevel_execute_ctrl0_up_DispatchPlugin_logic_hcs_3_onRs_0_ENABLES_0_lane0 = (((_zz_toplevel_execute_ctrl0_up_LANE_AGE_lane0 ? DispatchPlugin_logic_candidates_0_ctx_hm_DispatchPlugin_logic_hcs_3_onRs_0_ENABLES_0 : 1'b0) | (_zz_toplevel_execute_ctrl0_up_LANE_AGE_lane0_1 ? DispatchPlugin_logic_candidates_1_ctx_hm_DispatchPlugin_logic_hcs_3_onRs_0_ENABLES_0 : 1'b0)) | (_zz_toplevel_execute_ctrl0_up_LANE_AGE_lane0_2 ? DispatchPlugin_logic_candidates_2_ctx_hm_DispatchPlugin_logic_hcs_3_onRs_0_ENABLES_0 : 1'b0));
  assign _zz_toplevel_execute_ctrl0_up_DispatchPlugin_logic_hcs_3_onRs_1_ENABLES_0_lane0 = (((_zz_toplevel_execute_ctrl0_up_LANE_AGE_lane0 ? DispatchPlugin_logic_candidates_0_ctx_hm_DispatchPlugin_logic_hcs_3_onRs_1_ENABLES_0 : 1'b0) | (_zz_toplevel_execute_ctrl0_up_LANE_AGE_lane0_1 ? DispatchPlugin_logic_candidates_1_ctx_hm_DispatchPlugin_logic_hcs_3_onRs_1_ENABLES_0 : 1'b0)) | (_zz_toplevel_execute_ctrl0_up_LANE_AGE_lane0_2 ? DispatchPlugin_logic_candidates_2_ctx_hm_DispatchPlugin_logic_hcs_3_onRs_1_ENABLES_0 : 1'b0));
  assign _zz_DispatchPlugin_logic_inserter_1_trap = (((_zz_toplevel_execute_ctrl0_up_LANE_AGE_lane1 ? DispatchPlugin_logic_candidates_0_ctx_hm_TRAP : 1'b0) | (_zz_toplevel_execute_ctrl0_up_LANE_AGE_lane1_1 ? DispatchPlugin_logic_candidates_1_ctx_hm_TRAP : 1'b0)) | (_zz_toplevel_execute_ctrl0_up_LANE_AGE_lane1_2 ? DispatchPlugin_logic_candidates_2_ctx_hm_TRAP : 1'b0));
  assign _zz_toplevel_execute_ctrl0_up_LANE_SEL_lane1 = (((_zz_toplevel_execute_ctrl0_up_LANE_AGE_lane1 ? DispatchPlugin_logic_candidates_0_cancel : 1'b0) | (_zz_toplevel_execute_ctrl0_up_LANE_AGE_lane1_1 ? DispatchPlugin_logic_candidates_1_cancel : 1'b0)) | (_zz_toplevel_execute_ctrl0_up_LANE_AGE_lane1_2 ? DispatchPlugin_logic_candidates_2_cancel : 1'b0));
  assign _zz_toplevel_execute_ctrl0_up_Prediction_ALIGNED_JUMPED_lane1 = (((_zz_toplevel_execute_ctrl0_up_LANE_AGE_lane1 ? DispatchPlugin_logic_candidates_0_ctx_hm_Prediction_ALIGNED_JUMPED : 1'b0) | (_zz_toplevel_execute_ctrl0_up_LANE_AGE_lane1_1 ? DispatchPlugin_logic_candidates_1_ctx_hm_Prediction_ALIGNED_JUMPED : 1'b0)) | (_zz_toplevel_execute_ctrl0_up_LANE_AGE_lane1_2 ? DispatchPlugin_logic_candidates_2_ctx_hm_Prediction_ALIGNED_JUMPED : 1'b0));
  assign _zz_toplevel_execute_ctrl0_up_DispatchPlugin_FENCE_OLDER_lane1 = (((_zz_toplevel_execute_ctrl0_up_LANE_AGE_lane1 ? DispatchPlugin_logic_candidates_0_ctx_hm_DispatchPlugin_FENCE_OLDER : 1'b0) | (_zz_toplevel_execute_ctrl0_up_LANE_AGE_lane1_1 ? DispatchPlugin_logic_candidates_1_ctx_hm_DispatchPlugin_FENCE_OLDER : 1'b0)) | (_zz_toplevel_execute_ctrl0_up_LANE_AGE_lane1_2 ? DispatchPlugin_logic_candidates_2_ctx_hm_DispatchPlugin_FENCE_OLDER : 1'b0));
  assign _zz_toplevel_execute_ctrl0_up_DispatchPlugin_MAY_FLUSH_lane1 = (((_zz_toplevel_execute_ctrl0_up_LANE_AGE_lane1 ? DispatchPlugin_logic_candidates_0_ctx_hm_DispatchPlugin_MAY_FLUSH : 1'b0) | (_zz_toplevel_execute_ctrl0_up_LANE_AGE_lane1_1 ? DispatchPlugin_logic_candidates_1_ctx_hm_DispatchPlugin_MAY_FLUSH : 1'b0)) | (_zz_toplevel_execute_ctrl0_up_LANE_AGE_lane1_2 ? DispatchPlugin_logic_candidates_2_ctx_hm_DispatchPlugin_MAY_FLUSH : 1'b0));
  assign _zz_toplevel_execute_ctrl0_up_DispatchPlugin_DONT_FLUSH_lane1 = (((_zz_toplevel_execute_ctrl0_up_LANE_AGE_lane1 ? DispatchPlugin_logic_candidates_0_ctx_hm_DispatchPlugin_DONT_FLUSH : 1'b0) | (_zz_toplevel_execute_ctrl0_up_LANE_AGE_lane1_1 ? DispatchPlugin_logic_candidates_1_ctx_hm_DispatchPlugin_DONT_FLUSH : 1'b0)) | (_zz_toplevel_execute_ctrl0_up_LANE_AGE_lane1_2 ? DispatchPlugin_logic_candidates_2_ctx_hm_DispatchPlugin_DONT_FLUSH : 1'b0));
  assign _zz_toplevel_execute_ctrl0_up_DispatchPlugin_DONT_FLUSH_FROM_LANES_lane1 = (((_zz_toplevel_execute_ctrl0_up_LANE_AGE_lane1 ? DispatchPlugin_logic_candidates_0_ctx_hm_DispatchPlugin_DONT_FLUSH_FROM_LANES : 1'b0) | (_zz_toplevel_execute_ctrl0_up_LANE_AGE_lane1_1 ? DispatchPlugin_logic_candidates_1_ctx_hm_DispatchPlugin_DONT_FLUSH_FROM_LANES : 1'b0)) | (_zz_toplevel_execute_ctrl0_up_LANE_AGE_lane1_2 ? DispatchPlugin_logic_candidates_2_ctx_hm_DispatchPlugin_DONT_FLUSH_FROM_LANES : 1'b0));
  assign _zz_toplevel_execute_ctrl0_up_DONT_FLUSH_PRECISE_3_lane1 = (((_zz_toplevel_execute_ctrl0_up_LANE_AGE_lane1 ? DispatchPlugin_logic_candidates_0_ctx_hm_DONT_FLUSH_PRECISE_3 : 1'b0) | (_zz_toplevel_execute_ctrl0_up_LANE_AGE_lane1_1 ? DispatchPlugin_logic_candidates_1_ctx_hm_DONT_FLUSH_PRECISE_3 : 1'b0)) | (_zz_toplevel_execute_ctrl0_up_LANE_AGE_lane1_2 ? DispatchPlugin_logic_candidates_2_ctx_hm_DONT_FLUSH_PRECISE_3 : 1'b0));
  assign _zz_toplevel_execute_ctrl0_up_DONT_FLUSH_PRECISE_4_lane1 = (((_zz_toplevel_execute_ctrl0_up_LANE_AGE_lane1 ? DispatchPlugin_logic_candidates_0_ctx_hm_DONT_FLUSH_PRECISE_4 : 1'b0) | (_zz_toplevel_execute_ctrl0_up_LANE_AGE_lane1_1 ? DispatchPlugin_logic_candidates_1_ctx_hm_DONT_FLUSH_PRECISE_4 : 1'b0)) | (_zz_toplevel_execute_ctrl0_up_LANE_AGE_lane1_2 ? DispatchPlugin_logic_candidates_2_ctx_hm_DONT_FLUSH_PRECISE_4 : 1'b0));
  assign _zz_toplevel_execute_ctrl0_up_TRAP_lane1 = (((_zz_toplevel_execute_ctrl0_up_LANE_AGE_lane1 ? DispatchPlugin_logic_candidates_0_ctx_hm_TRAP : 1'b0) | (_zz_toplevel_execute_ctrl0_up_LANE_AGE_lane1_1 ? DispatchPlugin_logic_candidates_1_ctx_hm_TRAP : 1'b0)) | (_zz_toplevel_execute_ctrl0_up_LANE_AGE_lane1_2 ? DispatchPlugin_logic_candidates_2_ctx_hm_TRAP : 1'b0));
  assign _zz_toplevel_execute_ctrl0_up_RS1_ENABLE_lane1 = (((_zz_toplevel_execute_ctrl0_up_LANE_AGE_lane1 ? DispatchPlugin_logic_candidates_0_ctx_hm_RS1_ENABLE : 1'b0) | (_zz_toplevel_execute_ctrl0_up_LANE_AGE_lane1_1 ? DispatchPlugin_logic_candidates_1_ctx_hm_RS1_ENABLE : 1'b0)) | (_zz_toplevel_execute_ctrl0_up_LANE_AGE_lane1_2 ? DispatchPlugin_logic_candidates_2_ctx_hm_RS1_ENABLE : 1'b0));
  assign _zz_toplevel_execute_ctrl0_up_RS2_ENABLE_lane1 = (((_zz_toplevel_execute_ctrl0_up_LANE_AGE_lane1 ? DispatchPlugin_logic_candidates_0_ctx_hm_RS2_ENABLE : 1'b0) | (_zz_toplevel_execute_ctrl0_up_LANE_AGE_lane1_1 ? DispatchPlugin_logic_candidates_1_ctx_hm_RS2_ENABLE : 1'b0)) | (_zz_toplevel_execute_ctrl0_up_LANE_AGE_lane1_2 ? DispatchPlugin_logic_candidates_2_ctx_hm_RS2_ENABLE : 1'b0));
  assign _zz_toplevel_execute_ctrl0_up_RD_ENABLE_lane1 = (((_zz_toplevel_execute_ctrl0_up_LANE_AGE_lane1 ? DispatchPlugin_logic_candidates_0_ctx_hm_RD_ENABLE : 1'b0) | (_zz_toplevel_execute_ctrl0_up_LANE_AGE_lane1_1 ? DispatchPlugin_logic_candidates_1_ctx_hm_RD_ENABLE : 1'b0)) | (_zz_toplevel_execute_ctrl0_up_LANE_AGE_lane1_2 ? DispatchPlugin_logic_candidates_2_ctx_hm_RD_ENABLE : 1'b0));
  assign _zz_toplevel_execute_ctrl0_up_DispatchPlugin_logic_hcs_0_onRs_0_ENABLES_0_lane1 = (((_zz_toplevel_execute_ctrl0_up_LANE_AGE_lane1 ? DispatchPlugin_logic_candidates_0_ctx_hm_DispatchPlugin_logic_hcs_0_onRs_0_ENABLES_0 : 1'b0) | (_zz_toplevel_execute_ctrl0_up_LANE_AGE_lane1_1 ? DispatchPlugin_logic_candidates_1_ctx_hm_DispatchPlugin_logic_hcs_0_onRs_0_ENABLES_0 : 1'b0)) | (_zz_toplevel_execute_ctrl0_up_LANE_AGE_lane1_2 ? DispatchPlugin_logic_candidates_2_ctx_hm_DispatchPlugin_logic_hcs_0_onRs_0_ENABLES_0 : 1'b0));
  assign _zz_toplevel_execute_ctrl0_up_DispatchPlugin_logic_hcs_0_onRs_1_ENABLES_0_lane1 = (((_zz_toplevel_execute_ctrl0_up_LANE_AGE_lane1 ? DispatchPlugin_logic_candidates_0_ctx_hm_DispatchPlugin_logic_hcs_0_onRs_1_ENABLES_0 : 1'b0) | (_zz_toplevel_execute_ctrl0_up_LANE_AGE_lane1_1 ? DispatchPlugin_logic_candidates_1_ctx_hm_DispatchPlugin_logic_hcs_0_onRs_1_ENABLES_0 : 1'b0)) | (_zz_toplevel_execute_ctrl0_up_LANE_AGE_lane1_2 ? DispatchPlugin_logic_candidates_2_ctx_hm_DispatchPlugin_logic_hcs_0_onRs_1_ENABLES_0 : 1'b0));
  assign _zz_toplevel_execute_ctrl0_up_DispatchPlugin_logic_hcs_1_onRs_0_ENABLES_0_lane1 = (((_zz_toplevel_execute_ctrl0_up_LANE_AGE_lane1 ? DispatchPlugin_logic_candidates_0_ctx_hm_DispatchPlugin_logic_hcs_1_onRs_0_ENABLES_0 : 1'b0) | (_zz_toplevel_execute_ctrl0_up_LANE_AGE_lane1_1 ? DispatchPlugin_logic_candidates_1_ctx_hm_DispatchPlugin_logic_hcs_1_onRs_0_ENABLES_0 : 1'b0)) | (_zz_toplevel_execute_ctrl0_up_LANE_AGE_lane1_2 ? DispatchPlugin_logic_candidates_2_ctx_hm_DispatchPlugin_logic_hcs_1_onRs_0_ENABLES_0 : 1'b0));
  assign _zz_toplevel_execute_ctrl0_up_DispatchPlugin_logic_hcs_1_onRs_1_ENABLES_0_lane1 = (((_zz_toplevel_execute_ctrl0_up_LANE_AGE_lane1 ? DispatchPlugin_logic_candidates_0_ctx_hm_DispatchPlugin_logic_hcs_1_onRs_1_ENABLES_0 : 1'b0) | (_zz_toplevel_execute_ctrl0_up_LANE_AGE_lane1_1 ? DispatchPlugin_logic_candidates_1_ctx_hm_DispatchPlugin_logic_hcs_1_onRs_1_ENABLES_0 : 1'b0)) | (_zz_toplevel_execute_ctrl0_up_LANE_AGE_lane1_2 ? DispatchPlugin_logic_candidates_2_ctx_hm_DispatchPlugin_logic_hcs_1_onRs_1_ENABLES_0 : 1'b0));
  assign _zz_toplevel_execute_ctrl0_up_DispatchPlugin_logic_hcs_1_onRs_1_ENABLES_1_lane1 = (((_zz_toplevel_execute_ctrl0_up_LANE_AGE_lane1 ? DispatchPlugin_logic_candidates_0_ctx_hm_DispatchPlugin_logic_hcs_1_onRs_1_ENABLES_1 : 1'b0) | (_zz_toplevel_execute_ctrl0_up_LANE_AGE_lane1_1 ? DispatchPlugin_logic_candidates_1_ctx_hm_DispatchPlugin_logic_hcs_1_onRs_1_ENABLES_1 : 1'b0)) | (_zz_toplevel_execute_ctrl0_up_LANE_AGE_lane1_2 ? DispatchPlugin_logic_candidates_2_ctx_hm_DispatchPlugin_logic_hcs_1_onRs_1_ENABLES_1 : 1'b0));
  assign _zz_toplevel_execute_ctrl0_up_DispatchPlugin_logic_hcs_2_onRs_0_ENABLES_0_lane1 = (((_zz_toplevel_execute_ctrl0_up_LANE_AGE_lane1 ? DispatchPlugin_logic_candidates_0_ctx_hm_DispatchPlugin_logic_hcs_2_onRs_0_ENABLES_0 : 1'b0) | (_zz_toplevel_execute_ctrl0_up_LANE_AGE_lane1_1 ? DispatchPlugin_logic_candidates_1_ctx_hm_DispatchPlugin_logic_hcs_2_onRs_0_ENABLES_0 : 1'b0)) | (_zz_toplevel_execute_ctrl0_up_LANE_AGE_lane1_2 ? DispatchPlugin_logic_candidates_2_ctx_hm_DispatchPlugin_logic_hcs_2_onRs_0_ENABLES_0 : 1'b0));
  assign _zz_toplevel_execute_ctrl0_up_DispatchPlugin_logic_hcs_2_onRs_1_ENABLES_0_lane1 = (((_zz_toplevel_execute_ctrl0_up_LANE_AGE_lane1 ? DispatchPlugin_logic_candidates_0_ctx_hm_DispatchPlugin_logic_hcs_2_onRs_1_ENABLES_0 : 1'b0) | (_zz_toplevel_execute_ctrl0_up_LANE_AGE_lane1_1 ? DispatchPlugin_logic_candidates_1_ctx_hm_DispatchPlugin_logic_hcs_2_onRs_1_ENABLES_0 : 1'b0)) | (_zz_toplevel_execute_ctrl0_up_LANE_AGE_lane1_2 ? DispatchPlugin_logic_candidates_2_ctx_hm_DispatchPlugin_logic_hcs_2_onRs_1_ENABLES_0 : 1'b0));
  assign _zz_toplevel_execute_ctrl0_up_DispatchPlugin_logic_hcs_3_onRs_0_ENABLES_0_lane1 = (((_zz_toplevel_execute_ctrl0_up_LANE_AGE_lane1 ? DispatchPlugin_logic_candidates_0_ctx_hm_DispatchPlugin_logic_hcs_3_onRs_0_ENABLES_0 : 1'b0) | (_zz_toplevel_execute_ctrl0_up_LANE_AGE_lane1_1 ? DispatchPlugin_logic_candidates_1_ctx_hm_DispatchPlugin_logic_hcs_3_onRs_0_ENABLES_0 : 1'b0)) | (_zz_toplevel_execute_ctrl0_up_LANE_AGE_lane1_2 ? DispatchPlugin_logic_candidates_2_ctx_hm_DispatchPlugin_logic_hcs_3_onRs_0_ENABLES_0 : 1'b0));
  assign _zz_toplevel_execute_ctrl0_up_DispatchPlugin_logic_hcs_3_onRs_1_ENABLES_0_lane1 = (((_zz_toplevel_execute_ctrl0_up_LANE_AGE_lane1 ? DispatchPlugin_logic_candidates_0_ctx_hm_DispatchPlugin_logic_hcs_3_onRs_1_ENABLES_0 : 1'b0) | (_zz_toplevel_execute_ctrl0_up_LANE_AGE_lane1_1 ? DispatchPlugin_logic_candidates_1_ctx_hm_DispatchPlugin_logic_hcs_3_onRs_1_ENABLES_0 : 1'b0)) | (_zz_toplevel_execute_ctrl0_up_LANE_AGE_lane1_2 ? DispatchPlugin_logic_candidates_2_ctx_hm_DispatchPlugin_logic_hcs_3_onRs_1_ENABLES_0 : 1'b0));
  assign _zz_LsuL1Plugin_logic_shared_lsuRead_rsp_plru_0_1 = _zz_LsuL1Plugin_logic_shared_lsuRead_rsp_plru_0[0 : 0];
  assign _zz_LsuL1Plugin_logic_writeback_read_wordIndex_1 = LsuL1Plugin_logic_writeback_read_slotRead_valid;
  assign _zz_LsuL1Plugin_logic_writeback_read_wordIndex = {2'd0, _zz_LsuL1Plugin_logic_writeback_read_wordIndex_1};
  assign _zz_LsuL1Plugin_logic_writeback_write_wordIndex_1 = (LsuL1Plugin_logic_writeback_write_bufferRead_fire && 1'b1);
  assign _zz_LsuL1Plugin_logic_writeback_write_wordIndex = {2'd0, _zz_LsuL1Plugin_logic_writeback_write_wordIndex_1};
  assign _zz_LsuL1Plugin_logic_ls_ctrl_refillWayNeedWriteback = ({toplevel_execute_ctrl4_down_LsuL1Plugin_logic_WAYS_TAGS_lane0_1_loaded,toplevel_execute_ctrl4_down_LsuL1Plugin_logic_WAYS_TAGS_lane0_0_loaded} & toplevel_execute_ctrl4_down_LsuL1Plugin_logic_SHARED_lane0_dirty);
  assign _zz_LsuL1Plugin_logic_ls_ctrl_doWrite = ((_zz_toplevel_execute_ctrl4_down_LsuL1Plugin_logic_MUXED_DATA_lane0 ? (1'b1 && (! toplevel_execute_ctrl4_down_LsuL1Plugin_logic_WAYS_TAGS_lane0_0_fault)) : 1'b0) | (_zz_toplevel_execute_ctrl4_down_LsuL1Plugin_logic_MUXED_DATA_lane0_1 ? (1'b1 && (! toplevel_execute_ctrl4_down_LsuL1Plugin_logic_WAYS_TAGS_lane0_1_fault)) : 1'b0));
  assign _zz_LsuL1Plugin_logic_shared_write_payload_data_dirty = (2'b01 <<< LsuL1Plugin_logic_ls_ctrl_refillWayWithoutUpdate);
  assign _zz_LsuL1Plugin_logic_shared_write_payload_data_plru_0_1 = _zz_LsuL1Plugin_logic_shared_write_payload_data_plru_0[0 : 0];
  assign _zz_LsuPlugin_logic_onAddress0_ls_storeId_1 = LsuPlugin_logic_onAddress0_ls_port_fire;
  assign _zz_LsuPlugin_logic_onAddress0_ls_storeId = {11'd0, _zz_LsuPlugin_logic_onAddress0_ls_storeId_1};
  assign _zz_LsuPlugin_logic_onAddress0_flush_port_payload_address = ({6'd0,LsuPlugin_logic_flusher_cmdCounter} <<< 3'd6);
  assign _zz_LsuPlugin_logic_onPma_addressExtension = toplevel_execute_ctrl3_down_early0_SrcPlugin_ADD_SUB_lane0;
  assign _zz_LsuPlugin_logic_onCtrl_rva_alu_addSub = ($signed(_zz_LsuPlugin_logic_onCtrl_rva_alu_addSub_1) + $signed(_zz_LsuPlugin_logic_onCtrl_rva_alu_addSub_4));
  assign _zz_LsuPlugin_logic_onCtrl_rva_alu_addSub_1 = ($signed(_zz_LsuPlugin_logic_onCtrl_rva_alu_addSub_2) + $signed(_zz_LsuPlugin_logic_onCtrl_rva_alu_addSub_3));
  assign _zz_LsuPlugin_logic_onCtrl_rva_alu_addSub_2 = toplevel_execute_ctrl4_down_integer_RS2_lane0;
  assign _zz_LsuPlugin_logic_onCtrl_rva_alu_addSub_3 = (LsuPlugin_logic_onCtrl_rva_alu_compare ? (~ LsuPlugin_logic_onCtrl_rva_srcBuffer) : LsuPlugin_logic_onCtrl_rva_srcBuffer);
  assign _zz_LsuPlugin_logic_onCtrl_rva_alu_addSub_5 = (LsuPlugin_logic_onCtrl_rva_alu_compare ? 2'b01 : 2'b00);
  assign _zz_LsuPlugin_logic_onCtrl_rva_alu_addSub_4 = {{30{_zz_LsuPlugin_logic_onCtrl_rva_alu_addSub_5[1]}}, _zz_LsuPlugin_logic_onCtrl_rva_alu_addSub_5};
  assign _zz_LsuPlugin_logic_onCtrl_rva_nc_age_1 = (! execute_freeze_valid);
  assign _zz_LsuPlugin_logic_onCtrl_rva_nc_age = {5'd0, _zz_LsuPlugin_logic_onCtrl_rva_nc_age_1};
  assign _zz_LsuPlugin_logic_trapPort_payload_code = (toplevel_execute_ctrl4_down_LsuPlugin_logic_preCtrl_MISS_ALIGNED_lane0 ? (toplevel_execute_ctrl4_down_AguPlugin_STORE_lane0 ? 3'b110 : 3'b100) : 3'b000);
  assign _zz_LsuPlugin_logic_flusher_cmdCounter = toplevel_execute_ctrl4_down_LsuL1_MIXED_ADDRESS_lane0[11 : 6];
  assign _zz_TrapPlugin_logic_harts_0_trap_pending_slices_1 = ((_zz_TrapPlugin_logic_harts_0_trap_pending_pc ? toplevel_execute_ctrl4_down_Decode_INSTRUCTION_SLICE_COUNT_lane0 : 1'b0) | (_zz_TrapPlugin_logic_harts_0_trap_pending_pc_1 ? toplevel_execute_ctrl4_down_Decode_INSTRUCTION_SLICE_COUNT_lane1 : 1'b0));
  assign _zz_TrapPlugin_logic_harts_0_trap_pending_slices = {1'd0, _zz_TrapPlugin_logic_harts_0_trap_pending_slices_1};
  assign _zz_TrapPlugin_logic_harts_0_trap_fsm_jumpTarget_1 = ({1'd0,TrapPlugin_logic_harts_0_trap_fsm_jumpOffset} <<< 1'd1);
  assign _zz_TrapPlugin_logic_harts_0_trap_fsm_jumpTarget = {29'd0, _zz_TrapPlugin_logic_harts_0_trap_fsm_jumpTarget_1};
  assign _zz_LsuPlugin_logic_onAddress0_translationPort_logic_ctrl_lineAllowExecute_3 = (((_zz_LsuPlugin_logic_onAddress0_translationPort_logic_ctrl_lineAllowExecute ? toplevel_execute_ctrl3_down_MMU_L0_ENTRIES_lane0_0_allowExecute : 1'b0) | (_zz_LsuPlugin_logic_onAddress0_translationPort_logic_ctrl_lineAllowExecute_1 ? toplevel_execute_ctrl3_down_MMU_L0_ENTRIES_lane0_1_allowExecute : 1'b0)) | (_zz_LsuPlugin_logic_onAddress0_translationPort_logic_ctrl_lineAllowExecute_2 ? toplevel_execute_ctrl3_down_MMU_L1_ENTRIES_lane0_0_allowExecute : 1'b0));
  assign _zz_LsuPlugin_logic_onAddress0_translationPort_logic_ctrl_lineAllowRead = (((_zz_LsuPlugin_logic_onAddress0_translationPort_logic_ctrl_lineAllowExecute ? toplevel_execute_ctrl3_down_MMU_L0_ENTRIES_lane0_0_allowRead : 1'b0) | (_zz_LsuPlugin_logic_onAddress0_translationPort_logic_ctrl_lineAllowExecute_1 ? toplevel_execute_ctrl3_down_MMU_L0_ENTRIES_lane0_1_allowRead : 1'b0)) | (_zz_LsuPlugin_logic_onAddress0_translationPort_logic_ctrl_lineAllowExecute_2 ? toplevel_execute_ctrl3_down_MMU_L1_ENTRIES_lane0_0_allowRead : 1'b0));
  assign _zz_LsuPlugin_logic_onAddress0_translationPort_logic_ctrl_lineAllowWrite = (((_zz_LsuPlugin_logic_onAddress0_translationPort_logic_ctrl_lineAllowExecute ? toplevel_execute_ctrl3_down_MMU_L0_ENTRIES_lane0_0_allowWrite : 1'b0) | (_zz_LsuPlugin_logic_onAddress0_translationPort_logic_ctrl_lineAllowExecute_1 ? toplevel_execute_ctrl3_down_MMU_L0_ENTRIES_lane0_1_allowWrite : 1'b0)) | (_zz_LsuPlugin_logic_onAddress0_translationPort_logic_ctrl_lineAllowExecute_2 ? toplevel_execute_ctrl3_down_MMU_L1_ENTRIES_lane0_0_allowWrite : 1'b0));
  assign _zz_LsuPlugin_logic_onAddress0_translationPort_logic_ctrl_lineAllowUser = (((_zz_LsuPlugin_logic_onAddress0_translationPort_logic_ctrl_lineAllowExecute ? toplevel_execute_ctrl3_down_MMU_L0_ENTRIES_lane0_0_allowUser : 1'b0) | (_zz_LsuPlugin_logic_onAddress0_translationPort_logic_ctrl_lineAllowExecute_1 ? toplevel_execute_ctrl3_down_MMU_L0_ENTRIES_lane0_1_allowUser : 1'b0)) | (_zz_LsuPlugin_logic_onAddress0_translationPort_logic_ctrl_lineAllowExecute_2 ? toplevel_execute_ctrl3_down_MMU_L1_ENTRIES_lane0_0_allowUser : 1'b0));
  assign _zz_FetchL1Plugin_logic_translationPort_logic_ctrl_lineAllowExecute_3 = (((_zz_FetchL1Plugin_logic_translationPort_logic_ctrl_lineAllowExecute ? fetch_logic_ctrls_1_down_MMU_L0_ENTRIES_0_allowExecute : 1'b0) | (_zz_FetchL1Plugin_logic_translationPort_logic_ctrl_lineAllowExecute_1 ? fetch_logic_ctrls_1_down_MMU_L0_ENTRIES_1_allowExecute : 1'b0)) | (_zz_FetchL1Plugin_logic_translationPort_logic_ctrl_lineAllowExecute_2 ? fetch_logic_ctrls_1_down_MMU_L1_ENTRIES_0_allowExecute : 1'b0));
  assign _zz_FetchL1Plugin_logic_translationPort_logic_ctrl_lineAllowRead = (((_zz_FetchL1Plugin_logic_translationPort_logic_ctrl_lineAllowExecute ? fetch_logic_ctrls_1_down_MMU_L0_ENTRIES_0_allowRead : 1'b0) | (_zz_FetchL1Plugin_logic_translationPort_logic_ctrl_lineAllowExecute_1 ? fetch_logic_ctrls_1_down_MMU_L0_ENTRIES_1_allowRead : 1'b0)) | (_zz_FetchL1Plugin_logic_translationPort_logic_ctrl_lineAllowExecute_2 ? fetch_logic_ctrls_1_down_MMU_L1_ENTRIES_0_allowRead : 1'b0));
  assign _zz_FetchL1Plugin_logic_translationPort_logic_ctrl_lineAllowWrite = (((_zz_FetchL1Plugin_logic_translationPort_logic_ctrl_lineAllowExecute ? fetch_logic_ctrls_1_down_MMU_L0_ENTRIES_0_allowWrite : 1'b0) | (_zz_FetchL1Plugin_logic_translationPort_logic_ctrl_lineAllowExecute_1 ? fetch_logic_ctrls_1_down_MMU_L0_ENTRIES_1_allowWrite : 1'b0)) | (_zz_FetchL1Plugin_logic_translationPort_logic_ctrl_lineAllowExecute_2 ? fetch_logic_ctrls_1_down_MMU_L1_ENTRIES_0_allowWrite : 1'b0));
  assign _zz_FetchL1Plugin_logic_translationPort_logic_ctrl_lineAllowUser = (((_zz_FetchL1Plugin_logic_translationPort_logic_ctrl_lineAllowExecute ? fetch_logic_ctrls_1_down_MMU_L0_ENTRIES_0_allowUser : 1'b0) | (_zz_FetchL1Plugin_logic_translationPort_logic_ctrl_lineAllowExecute_1 ? fetch_logic_ctrls_1_down_MMU_L0_ENTRIES_1_allowUser : 1'b0)) | (_zz_FetchL1Plugin_logic_translationPort_logic_ctrl_lineAllowExecute_2 ? fetch_logic_ctrls_1_down_MMU_L1_ENTRIES_0_allowUser : 1'b0));
  assign _zz_PcPlugin_logic_harts_0_self_pc_1 = (PcPlugin_logic_harts_0_self_increment ? 4'b1000 : 4'b0000);
  assign _zz_PcPlugin_logic_harts_0_self_pc = {28'd0, _zz_PcPlugin_logic_harts_0_self_pc_1};
  assign _zz_PcPlugin_logic_harts_0_aggregator_fault = ((((_zz_PcPlugin_logic_harts_0_aggregator_target ? TrapPlugin_logic_harts_0_trap_pcPort_payload_fault : 1'b0) | (_zz_PcPlugin_logic_harts_0_aggregator_target_1 ? late0_BranchPlugin_logic_pcPort_payload_fault : 1'b0)) | ((_zz_PcPlugin_logic_harts_0_aggregator_target_2 ? late1_BranchPlugin_logic_pcPort_payload_fault : 1'b0) | (_zz_PcPlugin_logic_harts_0_aggregator_target_3 ? early0_BranchPlugin_logic_pcPort_payload_fault : 1'b0))) | (((_zz_PcPlugin_logic_harts_0_aggregator_target_4 ? early1_BranchPlugin_logic_pcPort_payload_fault : 1'b0) | (_zz_PcPlugin_logic_harts_0_aggregator_target_5 ? BtbPlugin_logic_pcPort_payload_fault : 1'b0)) | (_zz_PcPlugin_logic_harts_0_aggregator_target_6 ? PcPlugin_logic_harts_0_self_flow_payload_fault : 1'b0)));
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_15 = ((when_CsrService_l188 && REG_CSR_3858) ? 6'h2e : 6'h0);
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_14 = {26'd0, _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_15};
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_19 = ({7'd0,(_zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_1 ? PrivilegedPlugin_logic_harts_0_m_status_mpie : 1'b0)} <<< 3'd7);
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_18 = {24'd0, _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_19};
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_22 = ({3'd0,(_zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_1 ? PrivilegedPlugin_logic_harts_0_m_status_mie : 1'b0)} <<< 2'd3);
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_21 = {28'd0, _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_22};
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_24 = ({11'd0,(_zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_1 ? PrivilegedPlugin_logic_harts_0_m_status_mpp : 2'b00)} <<< 4'd11);
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_23 = {19'd0, _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_24};
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_26 = ({31'd0,(_zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_1 ? PrivilegedPlugin_logic_harts_0_m_status_sd : 1'b0)} <<< 5'd31);
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_28 = ({13'd0,(_zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_1 ? PrivilegedPlugin_logic_harts_0_m_status_fs : 2'b00)} <<< 4'd13);
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_27 = {17'd0, _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_28};
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_31 = ({22'd0,(_zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_1 ? PrivilegedPlugin_logic_harts_0_m_status_tsr : 1'b0)} <<< 5'd22);
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_30 = {9'd0, _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_31};
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_33 = ({20'd0,(_zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_1 ? PrivilegedPlugin_logic_harts_0_m_status_tvm : 1'b0)} <<< 5'd20);
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_32 = {11'd0, _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_33};
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_36 = ({21'd0,(_zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_1 ? PrivilegedPlugin_logic_harts_0_m_status_tw : 1'b0)} <<< 5'd21);
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_35 = {10'd0, _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_36};
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_37 = ({31'd0,(_zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_2 ? PrivilegedPlugin_logic_harts_0_m_cause_interrupt : 1'b0)} <<< 5'd31);
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_40 = (_zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_2 ? PrivilegedPlugin_logic_harts_0_m_cause_code : 4'b0000);
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_39 = {28'd0, _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_40};
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_42 = ({11'd0,(_zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_3 ? PrivilegedPlugin_logic_harts_0_m_ip_meip : 1'b0)} <<< 4'd11);
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_41 = {20'd0, _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_42};
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_45 = ({7'd0,(_zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_3 ? PrivilegedPlugin_logic_harts_0_m_ip_mtip : 1'b0)} <<< 3'd7);
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_44 = {24'd0, _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_45};
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_47 = ({3'd0,(_zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_3 ? PrivilegedPlugin_logic_harts_0_m_ip_msip : 1'b0)} <<< 2'd3);
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_46 = {28'd0, _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_47};
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_50 = ({11'd0,(_zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_4 ? PrivilegedPlugin_logic_harts_0_m_ie_meie : 1'b0)} <<< 4'd11);
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_49 = {20'd0, _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_50};
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_52 = ({7'd0,(_zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_4 ? PrivilegedPlugin_logic_harts_0_m_ie_mtie : 1'b0)} <<< 3'd7);
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_51 = {24'd0, _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_52};
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_55 = ({3'd0,(_zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_4 ? PrivilegedPlugin_logic_harts_0_m_ie_msie : 1'b0)} <<< 2'd3);
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_54 = {28'd0, _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_55};
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_57 = (_zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_5 ? PrivilegedPlugin_logic_harts_0_m_edeleg_iam : 1'b0);
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_56 = {31'd0, _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_57};
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_60 = ({3'd0,(_zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_5 ? PrivilegedPlugin_logic_harts_0_m_edeleg_bp : 1'b0)} <<< 2'd3);
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_59 = {28'd0, _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_60};
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_62 = ({8'd0,(_zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_5 ? PrivilegedPlugin_logic_harts_0_m_edeleg_eu : 1'b0)} <<< 4'd8);
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_61 = {23'd0, _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_62};
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_65 = ({9'd0,(_zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_5 ? PrivilegedPlugin_logic_harts_0_m_edeleg_es : 1'b0)} <<< 4'd9);
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_64 = {22'd0, _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_65};
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_67 = ({12'd0,(_zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_5 ? PrivilegedPlugin_logic_harts_0_m_edeleg_ipf : 1'b0)} <<< 4'd12);
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_66 = {19'd0, _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_67};
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_70 = ({13'd0,(_zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_5 ? PrivilegedPlugin_logic_harts_0_m_edeleg_lpf : 1'b0)} <<< 4'd13);
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_69 = {18'd0, _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_70};
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_72 = ({15'd0,(_zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_5 ? PrivilegedPlugin_logic_harts_0_m_edeleg_spf : 1'b0)} <<< 4'd15);
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_71 = {16'd0, _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_72};
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_75 = ({9'd0,(_zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_6 ? PrivilegedPlugin_logic_harts_0_m_ideleg_se : 1'b0)} <<< 4'd9);
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_74 = {22'd0, _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_75};
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_77 = ({5'd0,(_zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_6 ? PrivilegedPlugin_logic_harts_0_m_ideleg_st : 1'b0)} <<< 3'd5);
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_76 = {26'd0, _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_77};
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_80 = ({1'd0,(_zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_6 ? PrivilegedPlugin_logic_harts_0_m_ideleg_ss : 1'b0)} <<< 1'd1);
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_79 = {30'd0, _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_80};
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_81 = ({31'd0,(_zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_7 ? PrivilegedPlugin_logic_harts_0_s_cause_interrupt : 1'b0)} <<< 5'd31);
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_84 = (_zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_7 ? PrivilegedPlugin_logic_harts_0_s_cause_code : 4'b0000);
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_83 = {28'd0, _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_84};
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_85 = ({31'd0,(_zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_9 ? PrivilegedPlugin_logic_harts_0_m_status_sd : 1'b0)} <<< 5'd31);
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_88 = ({8'd0,(_zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_1 ? PrivilegedPlugin_logic_harts_0_s_status_spp : 1'b0)} <<< 4'd8);
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_87 = {23'd0, _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_88};
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_90 = ({5'd0,(_zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_1 ? PrivilegedPlugin_logic_harts_0_s_status_spie : 1'b0)} <<< 3'd5);
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_89 = {26'd0, _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_90};
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_93 = ({1'd0,(_zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_1 ? PrivilegedPlugin_logic_harts_0_s_status_sie : 1'b0)} <<< 1'd1);
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_92 = {30'd0, _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_93};
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_95 = ({8'd0,(_zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_9 ? PrivilegedPlugin_logic_harts_0_s_status_spp : 1'b0)} <<< 4'd8);
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_94 = {23'd0, _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_95};
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_98 = ({5'd0,(_zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_9 ? PrivilegedPlugin_logic_harts_0_s_status_spie : 1'b0)} <<< 3'd5);
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_97 = {26'd0, _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_98};
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_100 = ({1'd0,(_zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_9 ? PrivilegedPlugin_logic_harts_0_s_status_sie : 1'b0)} <<< 1'd1);
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_99 = {30'd0, _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_100};
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_103 = ({13'd0,(_zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_9 ? PrivilegedPlugin_logic_harts_0_m_status_fs : 2'b00)} <<< 4'd13);
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_102 = {17'd0, _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_103};
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_105 = ({9'd0,(_zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_4 ? PrivilegedPlugin_logic_harts_0_s_ie_seie : 1'b0)} <<< 4'd9);
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_104 = {22'd0, _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_105};
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_108 = ({9'd0,(_zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_10 ? (PrivilegedPlugin_logic_harts_0_s_ie_seie && PrivilegedPlugin_logic_harts_0_m_ideleg_se) : 1'b0)} <<< 4'd9);
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_107 = {22'd0, _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_108};
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_110 = ({5'd0,(_zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_4 ? PrivilegedPlugin_logic_harts_0_s_ie_stie : 1'b0)} <<< 3'd5);
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_109 = {26'd0, _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_110};
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_113 = ({5'd0,(_zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_10 ? (PrivilegedPlugin_logic_harts_0_s_ie_stie && PrivilegedPlugin_logic_harts_0_m_ideleg_st) : 1'b0)} <<< 3'd5);
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_112 = {26'd0, _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_113};
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_115 = ({1'd0,(_zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_4 ? PrivilegedPlugin_logic_harts_0_s_ie_ssie : 1'b0)} <<< 1'd1);
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_114 = {30'd0, _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_115};
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_118 = ({1'd0,(_zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_10 ? (PrivilegedPlugin_logic_harts_0_s_ie_ssie && PrivilegedPlugin_logic_harts_0_m_ideleg_ss) : 1'b0)} <<< 1'd1);
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_117 = {30'd0, _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_118};
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_120 = ({9'd0,(_zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_3 ? PrivilegedPlugin_logic_harts_0_s_ip_seipOr : 1'b0)} <<< 4'd9);
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_119 = {22'd0, _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_120};
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_123 = ({9'd0,(_zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_11 ? (PrivilegedPlugin_logic_harts_0_s_ip_seipOr && PrivilegedPlugin_logic_harts_0_m_ideleg_se) : 1'b0)} <<< 4'd9);
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_122 = {22'd0, _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_123};
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_125 = ({5'd0,(_zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_3 ? PrivilegedPlugin_logic_harts_0_s_ip_stip : 1'b0)} <<< 3'd5);
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_124 = {26'd0, _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_125};
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_128 = ({5'd0,(_zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_11 ? (PrivilegedPlugin_logic_harts_0_s_ip_stip && PrivilegedPlugin_logic_harts_0_m_ideleg_st) : 1'b0)} <<< 3'd5);
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_127 = {26'd0, _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_128};
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_130 = ({1'd0,(_zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_3 ? PrivilegedPlugin_logic_harts_0_s_ip_ssip : 1'b0)} <<< 1'd1);
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_129 = {30'd0, _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_130};
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_133 = ({1'd0,(_zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_11 ? (PrivilegedPlugin_logic_harts_0_s_ip_ssip && PrivilegedPlugin_logic_harts_0_m_ideleg_ss) : 1'b0)} <<< 1'd1);
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_132 = {30'd0, _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_133};
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_136 = ({19'd0,(_zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue ? MmuPlugin_logic_status_mxr : 1'b0)} <<< 5'd19);
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_135 = {12'd0, _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_136};
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_139 = ({18'd0,(_zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue ? MmuPlugin_logic_status_sum : 1'b0)} <<< 5'd18);
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_138 = {13'd0, _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_139};
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_141 = ({19'd0,(_zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_8 ? MmuPlugin_logic_status_mxr : 1'b0)} <<< 5'd19);
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_140 = {12'd0, _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_141};
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_144 = ({18'd0,(_zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_8 ? MmuPlugin_logic_status_sum : 1'b0)} <<< 5'd18);
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_143 = {13'd0, _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_144};
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_146 = ({17'd0,(_zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue ? MmuPlugin_logic_status_mprv : 1'b0)} <<< 5'd17);
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_145 = {14'd0, _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_146};
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_148 = ({31'd0,(_zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_12 ? MmuPlugin_logic_satp_mode : 1'b0)} <<< 5'd31);
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_150 = (_zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_12 ? MmuPlugin_logic_satp_ppn : 20'h0);
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_149 = {12'd0, _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_150};
  assign _zz_CsrAccessPlugin_logic_fsm_writeLogic_alu_mask_1 = CsrAccessPlugin_logic_fsm_regs_uop[19 : 15];
  assign _zz_CsrAccessPlugin_logic_fsm_writeLogic_alu_mask = {27'd0, _zz_CsrAccessPlugin_logic_fsm_writeLogic_alu_mask_1};
  assign _zz_CsrRamPlugin_logic_writeLogic_hits_ohFirst_masked = (CsrRamPlugin_logic_writeLogic_hits_ohFirst_input - 3'b001);
  assign _zz_CsrRamPlugin_logic_readLogic_hits_ohFirst_masked = (CsrRamPlugin_logic_readLogic_hits_ohFirst_input - 2'b01);
  assign _zz_CsrRamPlugin_logic_flush_counter_1 = (! CsrRamPlugin_logic_flush_done);
  assign _zz_CsrRamPlugin_logic_flush_counter = {3'd0, _zz_CsrRamPlugin_logic_flush_counter_1};
  assign _zz_toplevel_execute_ctrl1_down_early0_IntAluPlugin_SEL_lane0 = _zz_toplevel_execute_ctrl1_down_early0_IntAluPlugin_SEL_lane0_1[0];
  assign _zz_toplevel_execute_ctrl1_down_early0_IntAluPlugin_SEL_lane0_1 = (|{_zz_toplevel_execute_ctrl1_down_execute_lane0_logic_completions_onCtrl_0_ENABLE_lane0_3,{_zz_toplevel_execute_ctrl1_down_execute_lane0_logic_completions_onCtrl_0_ENABLE_lane0_2,{_zz_toplevel_execute_ctrl1_down_execute_lane0_logic_completions_onCtrl_0_ENABLE_lane0_1,{_zz_toplevel_execute_ctrl1_down_execute_lane0_logic_completions_onCtrl_0_ENABLE_lane0,((execute_lane0_logic_decoding_decodingBits & 33'h102001050) == 33'h100000010)}}}});
  assign _zz_toplevel_execute_ctrl1_down_early0_BarrelShifterPlugin_SEL_lane0 = _zz_toplevel_execute_ctrl1_down_early0_BarrelShifterPlugin_SEL_lane0_1[0];
  assign _zz_toplevel_execute_ctrl1_down_early0_BarrelShifterPlugin_SEL_lane0_1 = (|{_zz_toplevel_execute_ctrl1_down_execute_lane0_logic_completions_onCtrl_1_ENABLE_lane0,((execute_lane0_logic_decoding_decodingBits & 33'h102003054) == 33'h100001010)});
  assign _zz_toplevel_execute_ctrl1_down_early0_BranchPlugin_SEL_lane0 = _zz_toplevel_execute_ctrl1_down_early0_BranchPlugin_SEL_lane0_1[0];
  assign _zz_toplevel_execute_ctrl1_down_early0_BranchPlugin_SEL_lane0_1 = (|_zz_toplevel_execute_ctrl1_down_execute_lane0_logic_completions_onCtrl_1_ENABLE_lane0_1);
  assign _zz_toplevel_execute_ctrl1_down_early0_MulPlugin_SEL_lane0 = _zz_toplevel_execute_ctrl1_down_early0_MulPlugin_SEL_lane0_1[0];
  assign _zz_toplevel_execute_ctrl1_down_early0_MulPlugin_SEL_lane0_1 = (|((execute_lane0_logic_decoding_decodingBits & 33'h002004074) == 33'h002000030));
  assign _zz_toplevel_execute_ctrl1_down_early0_DivPlugin_SEL_lane0 = _zz_toplevel_execute_ctrl1_down_early0_DivPlugin_SEL_lane0_1[0];
  assign _zz_toplevel_execute_ctrl1_down_early0_DivPlugin_SEL_lane0_1 = (|_zz_toplevel_execute_ctrl1_down_execute_lane0_logic_completions_onCtrl_1_ENABLE_lane0_2);
  assign _zz_toplevel_execute_ctrl1_down_early0_EnvPlugin_SEL_lane0 = _zz_toplevel_execute_ctrl1_down_early0_EnvPlugin_SEL_lane0_1[0];
  assign _zz_toplevel_execute_ctrl1_down_early0_EnvPlugin_SEL_lane0_1 = (|{_zz_toplevel_execute_ctrl1_down_execute_lane0_logic_completions_onCtrl_0_ENABLE_lane0_4,((execute_lane0_logic_decoding_decodingBits & 33'h000003050) == 33'h000000050)});
  assign _zz_toplevel_execute_ctrl1_down_late0_IntAluPlugin_SEL_lane0 = _zz_toplevel_execute_ctrl1_down_late0_IntAluPlugin_SEL_lane0_1[0];
  assign _zz_toplevel_execute_ctrl1_down_late0_IntAluPlugin_SEL_lane0_1 = (|{((execute_lane0_logic_decoding_decodingBits & 33'h100000044) == 33'h000000004),{((execute_lane0_logic_decoding_decodingBits & 33'h100002040) == 33'h000002000),((execute_lane0_logic_decoding_decodingBits & 33'h100001040) == 33'h0)}});
  assign _zz_toplevel_execute_ctrl1_down_late0_BarrelShifterPlugin_SEL_lane0 = _zz_toplevel_execute_ctrl1_down_late0_BarrelShifterPlugin_SEL_lane0_1[0];
  assign _zz_toplevel_execute_ctrl1_down_late0_BarrelShifterPlugin_SEL_lane0_1 = (|((execute_lane0_logic_decoding_decodingBits & 33'h100003044) == 33'h000001000));
  assign _zz_toplevel_execute_ctrl1_down_late0_BranchPlugin_SEL_lane0_1 = _zz_toplevel_execute_ctrl1_down_late0_BranchPlugin_SEL_lane0_2[0];
  assign _zz_toplevel_execute_ctrl1_down_late0_BranchPlugin_SEL_lane0_2 = (|_zz_toplevel_execute_ctrl1_down_late0_BranchPlugin_SEL_lane0);
  assign _zz_toplevel_execute_ctrl1_down_MulPlugin_HIGH_lane0 = _zz_toplevel_execute_ctrl1_down_MulPlugin_HIGH_lane0_1[0];
  assign _zz_toplevel_execute_ctrl1_down_MulPlugin_HIGH_lane0_1 = (|{((execute_lane0_logic_decoding_decodingBits & 33'h002006074) == 33'h002002030),((execute_lane0_logic_decoding_decodingBits & 33'h002005074) == 33'h002001030)});
  assign _zz_toplevel_execute_ctrl1_down_CsrAccessPlugin_SEL_lane0 = _zz_toplevel_execute_ctrl1_down_CsrAccessPlugin_SEL_lane0_1[0];
  assign _zz_toplevel_execute_ctrl1_down_CsrAccessPlugin_SEL_lane0_1 = (|{((execute_lane0_logic_decoding_decodingBits & 33'h000001050) == 33'h000001050),((execute_lane0_logic_decoding_decodingBits & 33'h000002050) == 33'h000002050)});
  assign _zz_toplevel_execute_ctrl1_down_AguPlugin_SEL_lane0 = _zz_toplevel_execute_ctrl1_down_AguPlugin_SEL_lane0_1[0];
  assign _zz_toplevel_execute_ctrl1_down_AguPlugin_SEL_lane0_1 = (|{_zz_toplevel_execute_ctrl1_down_execute_lane0_logic_completions_onCtrl_2_ENABLE_lane0_1,_zz_toplevel_execute_ctrl1_down_execute_lane0_logic_completions_onCtrl_2_ENABLE_lane0});
  assign _zz_toplevel_execute_ctrl1_down_LsuPlugin_logic_FENCE_lane0 = _zz_toplevel_execute_ctrl1_down_LsuPlugin_logic_FENCE_lane0_1[0];
  assign _zz_toplevel_execute_ctrl1_down_LsuPlugin_logic_FENCE_lane0_1 = (|((execute_lane0_logic_decoding_decodingBits & 33'h000003048) == 33'h000000008));
  assign _zz_toplevel_execute_ctrl1_down_lane0_integer_WriteBackPlugin_SEL_lane0_1 = _zz_toplevel_execute_ctrl1_down_lane0_integer_WriteBackPlugin_SEL_lane0_2[0];
  assign _zz_toplevel_execute_ctrl1_down_lane0_integer_WriteBackPlugin_SEL_lane0_2 = (|{((execute_lane0_logic_decoding_decodingBits & 33'h000000048) == 33'h000000048),{((execute_lane0_logic_decoding_decodingBits & 33'h000001010) == 33'h000001010),{((execute_lane0_logic_decoding_decodingBits & 33'h000002010) == 33'h000002010),{_zz_toplevel_execute_ctrl1_down_AguPlugin_ATOMIC_lane0,{(_zz_toplevel_execute_ctrl1_down_lane0_integer_WriteBackPlugin_SEL_lane0_3 == _zz_toplevel_execute_ctrl1_down_lane0_integer_WriteBackPlugin_SEL_lane0_4),{_zz_toplevel_execute_ctrl1_down_lane0_integer_WriteBackPlugin_SEL_lane0,_zz_toplevel_execute_ctrl1_down_AguPlugin_LOAD_lane0}}}}}});
  assign _zz_toplevel_execute_ctrl1_down_COMPLETION_AT_2_lane0 = _zz_toplevel_execute_ctrl1_down_COMPLETION_AT_2_lane0_1[0];
  assign _zz_toplevel_execute_ctrl1_down_COMPLETION_AT_2_lane0_1 = (|{_zz_toplevel_execute_ctrl1_down_execute_lane0_logic_completions_onCtrl_0_ENABLE_lane0_4,{_zz_toplevel_execute_ctrl1_down_execute_lane0_logic_completions_onCtrl_0_ENABLE_lane0_3,{_zz_toplevel_execute_ctrl1_down_execute_lane0_logic_completions_onCtrl_0_ENABLE_lane0_2,{_zz_toplevel_execute_ctrl1_down_execute_lane0_logic_completions_onCtrl_0_ENABLE_lane0_1,{_zz_toplevel_execute_ctrl1_down_execute_lane0_logic_completions_onCtrl_0_ENABLE_lane0_6,{_zz_toplevel_execute_ctrl1_down_execute_lane0_logic_completions_onCtrl_0_ENABLE_lane0,_zz_toplevel_execute_ctrl1_down_execute_lane0_logic_completions_onCtrl_0_ENABLE_lane0_5}}}}}});
  assign _zz_toplevel_execute_ctrl1_down_COMPLETION_AT_3_lane0 = _zz_toplevel_execute_ctrl1_down_COMPLETION_AT_3_lane0_1[0];
  assign _zz_toplevel_execute_ctrl1_down_COMPLETION_AT_3_lane0_1 = (|{_zz_toplevel_execute_ctrl1_down_execute_lane0_logic_completions_onCtrl_1_ENABLE_lane0_5,{_zz_toplevel_execute_ctrl1_down_execute_lane0_logic_completions_onCtrl_1_ENABLE_lane0_4,{_zz_toplevel_execute_ctrl1_down_execute_lane0_logic_completions_onCtrl_1_ENABLE_lane0_1,{_zz_toplevel_execute_ctrl1_down_execute_lane0_logic_completions_onCtrl_1_ENABLE_lane0_2,{_zz_toplevel_execute_ctrl1_down_execute_lane0_logic_completions_onCtrl_1_ENABLE_lane0,_zz_toplevel_execute_ctrl1_down_execute_lane0_logic_completions_onCtrl_1_ENABLE_lane0_3}}}}});
  assign _zz_toplevel_execute_ctrl1_down_COMPLETION_AT_4_lane0 = _zz_toplevel_execute_ctrl1_down_COMPLETION_AT_4_lane0_1[0];
  assign _zz_toplevel_execute_ctrl1_down_COMPLETION_AT_4_lane0_1 = (|{_zz_toplevel_execute_ctrl1_down_execute_lane0_logic_completions_onCtrl_2_ENABLE_lane0_3,{_zz_toplevel_execute_ctrl1_down_execute_lane0_logic_completions_onCtrl_2_ENABLE_lane0_1,{_zz_toplevel_execute_ctrl1_down_execute_lane0_logic_completions_onCtrl_2_ENABLE_lane0,_zz_toplevel_execute_ctrl1_down_execute_lane0_logic_completions_onCtrl_2_ENABLE_lane0_2}}});
  assign _zz_toplevel_execute_ctrl1_down_execute_lane0_logic_completions_onCtrl_0_ENABLE_lane0_7 = _zz_toplevel_execute_ctrl1_down_execute_lane0_logic_completions_onCtrl_0_ENABLE_lane0_8[0];
  assign _zz_toplevel_execute_ctrl1_down_execute_lane0_logic_completions_onCtrl_0_ENABLE_lane0_8 = (|{_zz_toplevel_execute_ctrl1_down_execute_lane0_logic_completions_onCtrl_0_ENABLE_lane0_4,{_zz_toplevel_execute_ctrl1_down_execute_lane0_logic_completions_onCtrl_0_ENABLE_lane0_3,{_zz_toplevel_execute_ctrl1_down_execute_lane0_logic_completions_onCtrl_0_ENABLE_lane0_2,{_zz_toplevel_execute_ctrl1_down_execute_lane0_logic_completions_onCtrl_0_ENABLE_lane0_1,{_zz_toplevel_execute_ctrl1_down_execute_lane0_logic_completions_onCtrl_0_ENABLE_lane0_6,{_zz_toplevel_execute_ctrl1_down_execute_lane0_logic_completions_onCtrl_0_ENABLE_lane0,_zz_toplevel_execute_ctrl1_down_execute_lane0_logic_completions_onCtrl_0_ENABLE_lane0_5}}}}}});
  assign _zz_toplevel_execute_ctrl1_down_execute_lane0_logic_completions_onCtrl_1_ENABLE_lane0_6 = _zz_toplevel_execute_ctrl1_down_execute_lane0_logic_completions_onCtrl_1_ENABLE_lane0_7[0];
  assign _zz_toplevel_execute_ctrl1_down_execute_lane0_logic_completions_onCtrl_1_ENABLE_lane0_7 = (|{_zz_toplevel_execute_ctrl1_down_execute_lane0_logic_completions_onCtrl_1_ENABLE_lane0_5,{_zz_toplevel_execute_ctrl1_down_execute_lane0_logic_completions_onCtrl_1_ENABLE_lane0_4,{_zz_toplevel_execute_ctrl1_down_execute_lane0_logic_completions_onCtrl_1_ENABLE_lane0_1,{_zz_toplevel_execute_ctrl1_down_execute_lane0_logic_completions_onCtrl_1_ENABLE_lane0_2,{_zz_toplevel_execute_ctrl1_down_execute_lane0_logic_completions_onCtrl_1_ENABLE_lane0,_zz_toplevel_execute_ctrl1_down_execute_lane0_logic_completions_onCtrl_1_ENABLE_lane0_3}}}}});
  assign _zz_toplevel_execute_ctrl1_down_execute_lane0_logic_completions_onCtrl_2_ENABLE_lane0_4 = _zz_toplevel_execute_ctrl1_down_execute_lane0_logic_completions_onCtrl_2_ENABLE_lane0_5[0];
  assign _zz_toplevel_execute_ctrl1_down_execute_lane0_logic_completions_onCtrl_2_ENABLE_lane0_5 = (|{_zz_toplevel_execute_ctrl1_down_execute_lane0_logic_completions_onCtrl_2_ENABLE_lane0_3,{_zz_toplevel_execute_ctrl1_down_execute_lane0_logic_completions_onCtrl_2_ENABLE_lane0_1,{_zz_toplevel_execute_ctrl1_down_execute_lane0_logic_completions_onCtrl_2_ENABLE_lane0,_zz_toplevel_execute_ctrl1_down_execute_lane0_logic_completions_onCtrl_2_ENABLE_lane0_2}}});
  assign _zz_toplevel_execute_ctrl1_down_early0_IntAluPlugin_ALU_ADD_SUB_lane0 = _zz_toplevel_execute_ctrl1_down_early0_IntAluPlugin_ALU_ADD_SUB_lane0_1[0];
  assign _zz_toplevel_execute_ctrl1_down_early0_IntAluPlugin_ALU_ADD_SUB_lane0_1 = (|{_zz_toplevel_execute_ctrl1_down_late0_SrcPlugin_logic_SRC2_CTRL_lane0,_zz_toplevel_execute_ctrl1_down_late0_IntAluPlugin_ALU_ADD_SUB_lane0});
  assign _zz_toplevel_execute_ctrl1_down_early0_IntAluPlugin_ALU_SLTX_lane0 = _zz_toplevel_execute_ctrl1_down_early0_IntAluPlugin_ALU_SLTX_lane0_1[0];
  assign _zz_toplevel_execute_ctrl1_down_early0_IntAluPlugin_ALU_SLTX_lane0_1 = (|_zz_toplevel_execute_ctrl1_down_late0_IntAluPlugin_ALU_SLTX_lane0);
  assign _zz_toplevel_execute_ctrl1_down_SrcStageables_REVERT_lane0 = _zz_toplevel_execute_ctrl1_down_SrcStageables_REVERT_lane0_1[0];
  assign _zz_toplevel_execute_ctrl1_down_SrcStageables_REVERT_lane0_1 = (|{((execute_lane0_logic_decoding_decodingBits & 33'h000000040) == 33'h000000040),{((execute_lane0_logic_decoding_decodingBits & 33'h000002014) == 33'h000002010),((execute_lane0_logic_decoding_decodingBits & 33'h040000034) == 33'h040000030)}});
  assign _zz_toplevel_execute_ctrl1_down_SrcStageables_ZERO_lane0 = _zz_toplevel_execute_ctrl1_down_SrcStageables_ZERO_lane0_1[0];
  assign _zz_toplevel_execute_ctrl1_down_SrcStageables_ZERO_lane0_1 = (|((execute_lane0_logic_decoding_decodingBits & 33'h000000024) == 33'h000000024));
  assign _zz_toplevel_execute_ctrl1_down_lane0_IntFormatPlugin_logic_SIGNED_lane0 = _zz_toplevel_execute_ctrl1_down_lane0_IntFormatPlugin_logic_SIGNED_lane0_1[0];
  assign _zz_toplevel_execute_ctrl1_down_lane0_IntFormatPlugin_logic_SIGNED_lane0_1 = (|((execute_lane0_logic_decoding_decodingBits & 33'h000004010) == 33'h0));
  assign _zz_toplevel_execute_ctrl1_down_BYPASSED_AT_2_lane0 = _zz_toplevel_execute_ctrl1_down_BYPASSED_AT_2_lane0_1[0];
  assign _zz_toplevel_execute_ctrl1_down_BYPASSED_AT_2_lane0_1 = (|{_zz_toplevel_execute_ctrl1_down_execute_lane0_logic_completions_onCtrl_1_ENABLE_lane0_1,{_zz_toplevel_execute_ctrl1_down_BYPASSED_AT_3_lane0,{_zz_toplevel_execute_ctrl1_down_execute_lane0_logic_completions_onCtrl_0_ENABLE_lane0_3,{_zz_toplevel_execute_ctrl1_down_execute_lane0_logic_completions_onCtrl_0_ENABLE_lane0_1,{((execute_lane0_logic_decoding_decodingBits & 33'h102003020) == 33'h100000020),((execute_lane0_logic_decoding_decodingBits & 33'h102002068) == 33'h100002020)}}}}});
  assign _zz_toplevel_execute_ctrl1_down_BYPASSED_AT_3_lane0_1 = _zz_toplevel_execute_ctrl1_down_BYPASSED_AT_3_lane0_2[0];
  assign _zz_toplevel_execute_ctrl1_down_BYPASSED_AT_3_lane0_2 = (|{((execute_lane0_logic_decoding_decodingBits & 33'h100000040) == 33'h100000040),{((execute_lane0_logic_decoding_decodingBits & 33'h100004010) == 33'h100004010),{((execute_lane0_logic_decoding_decodingBits & 33'h100000030) == 33'h100000010),{_zz_toplevel_execute_ctrl1_down_BYPASSED_AT_3_lane0,((execute_lane0_logic_decoding_decodingBits & 33'h102000028) == 33'h100000020)}}}});
  assign _zz_toplevel_execute_ctrl1_down_MAY_FLUSH_PRECISE_3_lane0 = _zz_toplevel_execute_ctrl1_down_MAY_FLUSH_PRECISE_3_lane0_1[0];
  assign _zz_toplevel_execute_ctrl1_down_MAY_FLUSH_PRECISE_3_lane0_1 = (|{((execute_lane0_logic_decoding_decodingBits & 33'h000000050) == 33'h000000040),{_zz_toplevel_execute_ctrl1_down_SrcStageables_UNSIGNED_lane0,((execute_lane0_logic_decoding_decodingBits & 33'h000000018) == 33'h0)}});
  assign _zz_toplevel_execute_ctrl1_down_MAY_FLUSH_PRECISE_4_lane0 = _zz_toplevel_execute_ctrl1_down_MAY_FLUSH_PRECISE_4_lane0_1[0];
  assign _zz_toplevel_execute_ctrl1_down_MAY_FLUSH_PRECISE_4_lane0_1 = (|{_zz_toplevel_execute_ctrl1_down_late0_BranchPlugin_SEL_lane0,{((execute_lane0_logic_decoding_decodingBits & 33'h000002050) == 33'h000002000),_zz_toplevel_execute_ctrl1_down_execute_lane0_logic_completions_onCtrl_2_ENABLE_lane0}});
  assign _zz_toplevel_execute_ctrl1_down_SrcStageables_UNSIGNED_lane0_1 = _zz_toplevel_execute_ctrl1_down_SrcStageables_UNSIGNED_lane0_2[0];
  assign _zz_toplevel_execute_ctrl1_down_SrcStageables_UNSIGNED_lane0_2 = (|{_zz_toplevel_execute_ctrl1_down_SrcStageables_UNSIGNED_lane0,((execute_lane0_logic_decoding_decodingBits & 33'h000005000) == 33'h000001000)});
  assign _zz_toplevel_execute_ctrl1_down_BarrelShifterPlugin_LEFT_lane0_1 = _zz_toplevel_execute_ctrl1_down_BarrelShifterPlugin_LEFT_lane0_2[0];
  assign _zz_toplevel_execute_ctrl1_down_BarrelShifterPlugin_LEFT_lane0_2 = (|_zz_toplevel_execute_ctrl1_down_BarrelShifterPlugin_LEFT_lane0);
  assign _zz_toplevel_execute_ctrl1_down_BarrelShifterPlugin_SIGNED_lane0 = _zz_toplevel_execute_ctrl1_down_BarrelShifterPlugin_SIGNED_lane0_1[0];
  assign _zz_toplevel_execute_ctrl1_down_BarrelShifterPlugin_SIGNED_lane0_1 = (|((execute_lane0_logic_decoding_decodingBits & 33'h040000000) == 33'h040000000));
  assign _zz_toplevel_execute_ctrl1_down_RsUnsignedPlugin_RS1_SIGNED_lane0 = _zz_toplevel_execute_ctrl1_down_RsUnsignedPlugin_RS1_SIGNED_lane0_1[0];
  assign _zz_toplevel_execute_ctrl1_down_RsUnsignedPlugin_RS1_SIGNED_lane0_1 = (|{((execute_lane0_logic_decoding_decodingBits & 33'h000001000) == 33'h0),_zz_toplevel_execute_ctrl1_down_late0_IntAluPlugin_ALU_ADD_SUB_lane0});
  assign _zz_toplevel_execute_ctrl1_down_RsUnsignedPlugin_RS2_SIGNED_lane0 = _zz_toplevel_execute_ctrl1_down_RsUnsignedPlugin_RS2_SIGNED_lane0_1[0];
  assign _zz_toplevel_execute_ctrl1_down_RsUnsignedPlugin_RS2_SIGNED_lane0_1 = (|{((execute_lane0_logic_decoding_decodingBits & 33'h000005000) == 33'h000004000),_zz_toplevel_execute_ctrl1_down_late0_IntAluPlugin_ALU_ADD_SUB_lane0});
  assign _zz_toplevel_execute_ctrl1_down_DivPlugin_REM_lane0 = _zz_toplevel_execute_ctrl1_down_DivPlugin_REM_lane0_1[0];
  assign _zz_toplevel_execute_ctrl1_down_DivPlugin_REM_lane0_1 = (|_zz_toplevel_execute_ctrl1_down_CsrAccessPlugin_CSR_MASK_lane0);
  assign _zz_toplevel_execute_ctrl1_down_CsrAccessPlugin_CSR_IMM_lane0 = _zz_toplevel_execute_ctrl1_down_CsrAccessPlugin_CSR_IMM_lane0_1[0];
  assign _zz_toplevel_execute_ctrl1_down_CsrAccessPlugin_CSR_IMM_lane0_1 = (|((execute_lane0_logic_decoding_decodingBits & 33'h000004000) == 33'h000004000));
  assign _zz_toplevel_execute_ctrl1_down_CsrAccessPlugin_CSR_MASK_lane0_1 = _zz_toplevel_execute_ctrl1_down_CsrAccessPlugin_CSR_MASK_lane0_2[0];
  assign _zz_toplevel_execute_ctrl1_down_CsrAccessPlugin_CSR_MASK_lane0_2 = (|_zz_toplevel_execute_ctrl1_down_CsrAccessPlugin_CSR_MASK_lane0);
  assign _zz_toplevel_execute_ctrl1_down_CsrAccessPlugin_CSR_CLEAR_lane0_1 = _zz_toplevel_execute_ctrl1_down_CsrAccessPlugin_CSR_CLEAR_lane0_2[0];
  assign _zz_toplevel_execute_ctrl1_down_CsrAccessPlugin_CSR_CLEAR_lane0_2 = (|_zz_toplevel_execute_ctrl1_down_CsrAccessPlugin_CSR_CLEAR_lane0);
  assign _zz_toplevel_execute_ctrl1_down_AguPlugin_LOAD_lane0_1 = _zz_toplevel_execute_ctrl1_down_AguPlugin_LOAD_lane0_2[0];
  assign _zz_toplevel_execute_ctrl1_down_AguPlugin_LOAD_lane0_2 = (|{_zz_toplevel_execute_ctrl1_down_AguPlugin_LOAD_lane0,{((execute_lane0_logic_decoding_decodingBits & 33'h008002008) == 33'h000002008),((execute_lane0_logic_decoding_decodingBits & 33'h010002008) == 33'h000002008)}});
  assign _zz_toplevel_execute_ctrl1_down_AguPlugin_STORE_lane0_1 = _zz_toplevel_execute_ctrl1_down_AguPlugin_STORE_lane0_2[0];
  assign _zz_toplevel_execute_ctrl1_down_AguPlugin_STORE_lane0_2 = (|{((execute_lane0_logic_decoding_decodingBits & 33'h008000020) == 33'h008000020),{_zz_toplevel_execute_ctrl1_down_AguPlugin_STORE_lane0,((execute_lane0_logic_decoding_decodingBits & 33'h000000028) == 33'h000000020)}});
  assign _zz_toplevel_execute_ctrl1_down_AguPlugin_ATOMIC_lane0_1 = _zz_toplevel_execute_ctrl1_down_AguPlugin_ATOMIC_lane0_2[0];
  assign _zz_toplevel_execute_ctrl1_down_AguPlugin_ATOMIC_lane0_2 = (|_zz_toplevel_execute_ctrl1_down_AguPlugin_ATOMIC_lane0);
  assign _zz_toplevel_execute_ctrl1_down_AguPlugin_FLOAT_lane0 = _zz_toplevel_execute_ctrl1_down_AguPlugin_FLOAT_lane0_1[0];
  assign _zz_toplevel_execute_ctrl1_down_AguPlugin_FLOAT_lane0_1 = 1'b0;
  assign _zz_toplevel_execute_ctrl1_down_LsuPlugin_logic_LSU_PREFETCH_lane0 = _zz_toplevel_execute_ctrl1_down_LsuPlugin_logic_LSU_PREFETCH_lane0_1[0];
  assign _zz_toplevel_execute_ctrl1_down_LsuPlugin_logic_LSU_PREFETCH_lane0_1 = 1'b0;
  assign _zz_toplevel_execute_ctrl1_down_late0_IntAluPlugin_ALU_ADD_SUB_lane0_1 = _zz_toplevel_execute_ctrl1_down_late0_IntAluPlugin_ALU_ADD_SUB_lane0_2[0];
  assign _zz_toplevel_execute_ctrl1_down_late0_IntAluPlugin_ALU_ADD_SUB_lane0_2 = (|{_zz_toplevel_execute_ctrl1_down_late0_SrcPlugin_logic_SRC2_CTRL_lane0,_zz_toplevel_execute_ctrl1_down_late0_IntAluPlugin_ALU_ADD_SUB_lane0});
  assign _zz_toplevel_execute_ctrl1_down_late0_IntAluPlugin_ALU_SLTX_lane0_1 = _zz_toplevel_execute_ctrl1_down_late0_IntAluPlugin_ALU_SLTX_lane0_2[0];
  assign _zz_toplevel_execute_ctrl1_down_late0_IntAluPlugin_ALU_SLTX_lane0_2 = (|_zz_toplevel_execute_ctrl1_down_late0_IntAluPlugin_ALU_SLTX_lane0);
  assign _zz_WhiteboxerPlugin_logic_csr_access_payload_address = CsrAccessPlugin_logic_fsm_regs_uop;
  assign _zz_toplevel_execute_ctrl1_down_early1_IntAluPlugin_SEL_lane1 = _zz_toplevel_execute_ctrl1_down_early1_IntAluPlugin_SEL_lane1_1[0];
  assign _zz_toplevel_execute_ctrl1_down_early1_IntAluPlugin_SEL_lane1_1 = (|{_zz_toplevel_execute_ctrl1_down_execute_lane1_logic_completions_onCtrl_0_ENABLE_lane1_2,{_zz_toplevel_execute_ctrl1_down_execute_lane1_logic_completions_onCtrl_0_ENABLE_lane1_1,_zz_toplevel_execute_ctrl1_down_execute_lane1_logic_completions_onCtrl_0_ENABLE_lane1}});
  assign _zz_toplevel_execute_ctrl1_down_early1_BarrelShifterPlugin_SEL_lane1 = _zz_toplevel_execute_ctrl1_down_early1_BarrelShifterPlugin_SEL_lane1_1[0];
  assign _zz_toplevel_execute_ctrl1_down_early1_BarrelShifterPlugin_SEL_lane1_1 = (|((execute_lane1_logic_decoding_decodingBits & 33'h100003044) == 33'h100001000));
  assign _zz_toplevel_execute_ctrl1_down_early1_BranchPlugin_SEL_lane1 = _zz_toplevel_execute_ctrl1_down_early1_BranchPlugin_SEL_lane1_1[0];
  assign _zz_toplevel_execute_ctrl1_down_early1_BranchPlugin_SEL_lane1_1 = (|_zz_toplevel_execute_ctrl1_down_execute_lane1_logic_completions_onCtrl_1_ENABLE_lane1);
  assign _zz_toplevel_execute_ctrl1_down_late1_IntAluPlugin_SEL_lane1 = _zz_toplevel_execute_ctrl1_down_late1_IntAluPlugin_SEL_lane1_1[0];
  assign _zz_toplevel_execute_ctrl1_down_late1_IntAluPlugin_SEL_lane1_1 = (|{((execute_lane1_logic_decoding_decodingBits & 33'h100000044) == 33'h000000004),{((execute_lane1_logic_decoding_decodingBits & 33'h100002040) == 33'h000002000),((execute_lane1_logic_decoding_decodingBits & 33'h100001040) == 33'h0)}});
  assign _zz_toplevel_execute_ctrl1_down_late1_BarrelShifterPlugin_SEL_lane1 = _zz_toplevel_execute_ctrl1_down_late1_BarrelShifterPlugin_SEL_lane1_1[0];
  assign _zz_toplevel_execute_ctrl1_down_late1_BarrelShifterPlugin_SEL_lane1_1 = (|((execute_lane1_logic_decoding_decodingBits & 33'h100003044) == 33'h000001000));
  assign _zz_toplevel_execute_ctrl1_down_late1_BranchPlugin_SEL_lane1_1 = _zz_toplevel_execute_ctrl1_down_late1_BranchPlugin_SEL_lane1_2[0];
  assign _zz_toplevel_execute_ctrl1_down_late1_BranchPlugin_SEL_lane1_2 = (|_zz_toplevel_execute_ctrl1_down_late1_BranchPlugin_SEL_lane1);
  assign _zz_toplevel_execute_ctrl1_down_lane1_integer_WriteBackPlugin_SEL_lane1 = _zz_toplevel_execute_ctrl1_down_lane1_integer_WriteBackPlugin_SEL_lane1_1[0];
  assign _zz_toplevel_execute_ctrl1_down_lane1_integer_WriteBackPlugin_SEL_lane1_1 = (|{_zz_toplevel_execute_ctrl1_down_late1_SrcPlugin_logic_SRC2_CTRL_lane1,((execute_lane1_logic_decoding_decodingBits & 33'h000000040) == 33'h0)});
  assign _zz_toplevel_execute_ctrl1_down_COMPLETION_AT_2_lane1 = _zz_toplevel_execute_ctrl1_down_COMPLETION_AT_2_lane1_1[0];
  assign _zz_toplevel_execute_ctrl1_down_COMPLETION_AT_2_lane1_1 = (|{_zz_toplevel_execute_ctrl1_down_execute_lane1_logic_completions_onCtrl_0_ENABLE_lane1_2,{_zz_toplevel_execute_ctrl1_down_execute_lane1_logic_completions_onCtrl_0_ENABLE_lane1_1,_zz_toplevel_execute_ctrl1_down_execute_lane1_logic_completions_onCtrl_0_ENABLE_lane1}});
  assign _zz_toplevel_execute_ctrl1_down_COMPLETION_AT_3_lane1 = _zz_toplevel_execute_ctrl1_down_COMPLETION_AT_3_lane1_1[0];
  assign _zz_toplevel_execute_ctrl1_down_COMPLETION_AT_3_lane1_1 = (|{_zz_toplevel_execute_ctrl1_down_execute_lane1_logic_completions_onCtrl_1_ENABLE_lane1,_zz_toplevel_execute_ctrl1_down_execute_lane1_logic_completions_onCtrl_1_ENABLE_lane1_1});
  assign _zz_toplevel_execute_ctrl1_down_COMPLETION_AT_4_lane1 = _zz_toplevel_execute_ctrl1_down_COMPLETION_AT_4_lane1_1[0];
  assign _zz_toplevel_execute_ctrl1_down_COMPLETION_AT_4_lane1_1 = (|_zz_toplevel_execute_ctrl1_down_execute_lane1_logic_completions_onCtrl_2_ENABLE_lane1);
  assign _zz_toplevel_execute_ctrl1_down_execute_lane1_logic_completions_onCtrl_0_ENABLE_lane1_3 = _zz_toplevel_execute_ctrl1_down_execute_lane1_logic_completions_onCtrl_0_ENABLE_lane1_4[0];
  assign _zz_toplevel_execute_ctrl1_down_execute_lane1_logic_completions_onCtrl_0_ENABLE_lane1_4 = (|{_zz_toplevel_execute_ctrl1_down_execute_lane1_logic_completions_onCtrl_0_ENABLE_lane1_2,{_zz_toplevel_execute_ctrl1_down_execute_lane1_logic_completions_onCtrl_0_ENABLE_lane1_1,_zz_toplevel_execute_ctrl1_down_execute_lane1_logic_completions_onCtrl_0_ENABLE_lane1}});
  assign _zz_toplevel_execute_ctrl1_down_execute_lane1_logic_completions_onCtrl_1_ENABLE_lane1_2 = _zz_toplevel_execute_ctrl1_down_execute_lane1_logic_completions_onCtrl_1_ENABLE_lane1_3[0];
  assign _zz_toplevel_execute_ctrl1_down_execute_lane1_logic_completions_onCtrl_1_ENABLE_lane1_3 = (|{_zz_toplevel_execute_ctrl1_down_execute_lane1_logic_completions_onCtrl_1_ENABLE_lane1,_zz_toplevel_execute_ctrl1_down_execute_lane1_logic_completions_onCtrl_1_ENABLE_lane1_1});
  assign _zz_toplevel_execute_ctrl1_down_execute_lane1_logic_completions_onCtrl_2_ENABLE_lane1_1 = _zz_toplevel_execute_ctrl1_down_execute_lane1_logic_completions_onCtrl_2_ENABLE_lane1_2[0];
  assign _zz_toplevel_execute_ctrl1_down_execute_lane1_logic_completions_onCtrl_2_ENABLE_lane1_2 = (|_zz_toplevel_execute_ctrl1_down_execute_lane1_logic_completions_onCtrl_2_ENABLE_lane1);
  assign _zz_toplevel_execute_ctrl1_down_early1_IntAluPlugin_ALU_ADD_SUB_lane1 = _zz_toplevel_execute_ctrl1_down_early1_IntAluPlugin_ALU_ADD_SUB_lane1_1[0];
  assign _zz_toplevel_execute_ctrl1_down_early1_IntAluPlugin_ALU_ADD_SUB_lane1_1 = (|{_zz_toplevel_execute_ctrl1_down_late1_SrcPlugin_logic_SRC2_CTRL_lane1,_zz_toplevel_execute_ctrl1_down_late1_IntAluPlugin_ALU_ADD_SUB_lane1});
  assign _zz_toplevel_execute_ctrl1_down_early1_IntAluPlugin_ALU_SLTX_lane1 = _zz_toplevel_execute_ctrl1_down_early1_IntAluPlugin_ALU_SLTX_lane1_1[0];
  assign _zz_toplevel_execute_ctrl1_down_early1_IntAluPlugin_ALU_SLTX_lane1_1 = (|_zz_toplevel_execute_ctrl1_down_late1_IntAluPlugin_ALU_SLTX_lane1);
  assign _zz_toplevel_execute_ctrl1_down_SrcStageables_REVERT_lane1_1 = _zz_toplevel_execute_ctrl1_down_SrcStageables_REVERT_lane1_2[0];
  assign _zz_toplevel_execute_ctrl1_down_SrcStageables_REVERT_lane1_2 = (|{_zz_toplevel_execute_ctrl1_down_SrcStageables_REVERT_lane1,{((execute_lane1_logic_decoding_decodingBits & 33'h000002004) == 33'h000002000),((execute_lane1_logic_decoding_decodingBits & 33'h040000024) == 33'h040000020)}});
  assign _zz_toplevel_execute_ctrl1_down_SrcStageables_ZERO_lane1 = _zz_toplevel_execute_ctrl1_down_SrcStageables_ZERO_lane1_1[0];
  assign _zz_toplevel_execute_ctrl1_down_SrcStageables_ZERO_lane1_1 = (|((execute_lane1_logic_decoding_decodingBits & 33'h000000024) == 33'h000000024));
  assign _zz_toplevel_execute_ctrl1_down_lane1_IntFormatPlugin_logic_SIGNED_lane1 = _zz_toplevel_execute_ctrl1_down_lane1_IntFormatPlugin_logic_SIGNED_lane1_1[0];
  assign _zz_toplevel_execute_ctrl1_down_lane1_IntFormatPlugin_logic_SIGNED_lane1_1 = 1'b0;
  assign _zz_toplevel_execute_ctrl1_down_BYPASSED_AT_2_lane1 = _zz_toplevel_execute_ctrl1_down_BYPASSED_AT_2_lane1_1[0];
  assign _zz_toplevel_execute_ctrl1_down_BYPASSED_AT_2_lane1_1 = (|{((execute_lane1_logic_decoding_decodingBits & 33'h100000004) == 33'h100000004),{((execute_lane1_logic_decoding_decodingBits & 33'h100002000) == 33'h100002000),((execute_lane1_logic_decoding_decodingBits & 33'h100001000) == 33'h100000000)}});
  assign _zz_toplevel_execute_ctrl1_down_BYPASSED_AT_3_lane1 = _zz_toplevel_execute_ctrl1_down_BYPASSED_AT_3_lane1_1[0];
  assign _zz_toplevel_execute_ctrl1_down_BYPASSED_AT_3_lane1_1 = (|((execute_lane1_logic_decoding_decodingBits & 33'h100000000) == 33'h100000000));
  assign _zz_toplevel_execute_ctrl1_down_MAY_FLUSH_PRECISE_3_lane1 = _zz_toplevel_execute_ctrl1_down_MAY_FLUSH_PRECISE_3_lane1_1[0];
  assign _zz_toplevel_execute_ctrl1_down_MAY_FLUSH_PRECISE_3_lane1_1 = (|_zz_toplevel_execute_ctrl1_down_SrcStageables_REVERT_lane1);
  assign _zz_toplevel_execute_ctrl1_down_MAY_FLUSH_PRECISE_4_lane1 = _zz_toplevel_execute_ctrl1_down_MAY_FLUSH_PRECISE_4_lane1_1[0];
  assign _zz_toplevel_execute_ctrl1_down_MAY_FLUSH_PRECISE_4_lane1_1 = (|_zz_toplevel_execute_ctrl1_down_late1_BranchPlugin_SEL_lane1);
  assign _zz_toplevel_execute_ctrl1_down_SrcStageables_UNSIGNED_lane1 = _zz_toplevel_execute_ctrl1_down_SrcStageables_UNSIGNED_lane1_1[0];
  assign _zz_toplevel_execute_ctrl1_down_SrcStageables_UNSIGNED_lane1_1 = (|{((execute_lane1_logic_decoding_decodingBits & 33'h000002010) == 33'h000002000),((execute_lane1_logic_decoding_decodingBits & 33'h000005000) == 33'h000001000)});
  assign _zz_toplevel_execute_ctrl1_down_BarrelShifterPlugin_LEFT_lane1_1 = _zz_toplevel_execute_ctrl1_down_BarrelShifterPlugin_LEFT_lane1_2[0];
  assign _zz_toplevel_execute_ctrl1_down_BarrelShifterPlugin_LEFT_lane1_2 = (|_zz_toplevel_execute_ctrl1_down_BarrelShifterPlugin_LEFT_lane1);
  assign _zz_toplevel_execute_ctrl1_down_BarrelShifterPlugin_SIGNED_lane1 = _zz_toplevel_execute_ctrl1_down_BarrelShifterPlugin_SIGNED_lane1_1[0];
  assign _zz_toplevel_execute_ctrl1_down_BarrelShifterPlugin_SIGNED_lane1_1 = (|((execute_lane1_logic_decoding_decodingBits & 33'h040000000) == 33'h040000000));
  assign _zz_toplevel_execute_ctrl1_down_late1_IntAluPlugin_ALU_ADD_SUB_lane1_1 = _zz_toplevel_execute_ctrl1_down_late1_IntAluPlugin_ALU_ADD_SUB_lane1_2[0];
  assign _zz_toplevel_execute_ctrl1_down_late1_IntAluPlugin_ALU_ADD_SUB_lane1_2 = (|{_zz_toplevel_execute_ctrl1_down_late1_SrcPlugin_logic_SRC2_CTRL_lane1,_zz_toplevel_execute_ctrl1_down_late1_IntAluPlugin_ALU_ADD_SUB_lane1});
  assign _zz_toplevel_execute_ctrl1_down_late1_IntAluPlugin_ALU_SLTX_lane1_1 = _zz_toplevel_execute_ctrl1_down_late1_IntAluPlugin_ALU_SLTX_lane1_2[0];
  assign _zz_toplevel_execute_ctrl1_down_late1_IntAluPlugin_ALU_SLTX_lane1_2 = (|_zz_toplevel_execute_ctrl1_down_late1_IntAluPlugin_ALU_SLTX_lane1);
  assign _zz_FetchL1Plugin_pmaBuilder_onTransfers_0_addressHit = (|_zz_FetchL1Plugin_logic_ctrl_pmaPort_rsp_io);
  assign _zz_FetchL1Plugin_logic_ctrl_pmaPort_rsp_io_1 = (|_zz_FetchL1Plugin_logic_ctrl_pmaPort_rsp_io);
  assign _zz_LsuPlugin_pmaBuilder_l1_onTransfers_0_addressHit = (|_zz_LsuPlugin_logic_onPma_cached_rsp_io);
  assign _zz_LsuPlugin_logic_onPma_cached_rsp_io_1 = (|_zz_LsuPlugin_logic_onPma_cached_rsp_io);
  assign _zz_LsuPlugin_pmaBuilder_io_onTransfers_0_addressHit = (|((LsuPlugin_pmaBuilder_io_addressBits & 32'hc0000000) == 32'h0));
  assign _zz_LsuPlugin_pmaBuilder_io_onTransfers_1_addressHit = (|{_zz_LsuPlugin_logic_onPma_io_rsp_io_1,_zz_LsuPlugin_logic_onPma_io_rsp_io});
  assign _zz_LsuPlugin_logic_onPma_io_rsp_io_2 = (|{_zz_LsuPlugin_logic_onPma_io_rsp_io_1,_zz_LsuPlugin_logic_onPma_io_rsp_io});
  assign _zz__zz_WhiteboxerPlugin_logic_perf_executeFreezedCounter_1_1 = _zz_WhiteboxerPlugin_logic_perf_executeFreezedCounter;
  assign _zz__zz_WhiteboxerPlugin_logic_perf_executeFreezedCounter_1 = {59'd0, _zz__zz_WhiteboxerPlugin_logic_perf_executeFreezedCounter_1_1};
  assign _zz__zz_WhiteboxerPlugin_logic_perf_dispatchHazardsCounter_1_1 = _zz_WhiteboxerPlugin_logic_perf_dispatchHazardsCounter;
  assign _zz__zz_WhiteboxerPlugin_logic_perf_dispatchHazardsCounter_1 = {59'd0, _zz__zz_WhiteboxerPlugin_logic_perf_dispatchHazardsCounter_1_1};
  assign _zz__zz_WhiteboxerPlugin_logic_perf_candidatesCountCounters_0_1_1 = _zz_WhiteboxerPlugin_logic_perf_candidatesCountCounters_0;
  assign _zz__zz_WhiteboxerPlugin_logic_perf_candidatesCountCounters_0_1 = {59'd0, _zz__zz_WhiteboxerPlugin_logic_perf_candidatesCountCounters_0_1_1};
  assign _zz__zz_WhiteboxerPlugin_logic_perf_candidatesCountCounters_1_1_1 = _zz_WhiteboxerPlugin_logic_perf_candidatesCountCounters_1;
  assign _zz__zz_WhiteboxerPlugin_logic_perf_candidatesCountCounters_1_1 = {59'd0, _zz__zz_WhiteboxerPlugin_logic_perf_candidatesCountCounters_1_1_1};
  assign _zz__zz_WhiteboxerPlugin_logic_perf_candidatesCountCounters_2_1_1 = _zz_WhiteboxerPlugin_logic_perf_candidatesCountCounters_2;
  assign _zz__zz_WhiteboxerPlugin_logic_perf_candidatesCountCounters_2_1 = {59'd0, _zz__zz_WhiteboxerPlugin_logic_perf_candidatesCountCounters_2_1_1};
  assign _zz__zz_WhiteboxerPlugin_logic_perf_candidatesCountCounters_3_1_1 = _zz_WhiteboxerPlugin_logic_perf_candidatesCountCounters_3;
  assign _zz__zz_WhiteboxerPlugin_logic_perf_candidatesCountCounters_3_1 = {59'd0, _zz__zz_WhiteboxerPlugin_logic_perf_candidatesCountCounters_3_1_1};
  assign _zz__zz_WhiteboxerPlugin_logic_perf_dispatchFeedCounters_0_1_1 = _zz_WhiteboxerPlugin_logic_perf_dispatchFeedCounters_0;
  assign _zz__zz_WhiteboxerPlugin_logic_perf_dispatchFeedCounters_0_1 = {59'd0, _zz__zz_WhiteboxerPlugin_logic_perf_dispatchFeedCounters_0_1_1};
  assign _zz__zz_WhiteboxerPlugin_logic_perf_dispatchFeedCounters_1_1_1 = _zz_WhiteboxerPlugin_logic_perf_dispatchFeedCounters_1;
  assign _zz__zz_WhiteboxerPlugin_logic_perf_dispatchFeedCounters_1_1 = {59'd0, _zz__zz_WhiteboxerPlugin_logic_perf_dispatchFeedCounters_1_1_1};
  assign _zz__zz_WhiteboxerPlugin_logic_perf_dispatchFeedCounters_2_1_1 = _zz_WhiteboxerPlugin_logic_perf_dispatchFeedCounters_2;
  assign _zz__zz_WhiteboxerPlugin_logic_perf_dispatchFeedCounters_2_1 = {59'd0, _zz__zz_WhiteboxerPlugin_logic_perf_dispatchFeedCounters_2_1_1};
  assign _zz_FetchL1Plugin_logic_translationStorage_logic_sl_0_write_mask = (2'b01 <<< FetchL1Plugin_logic_translationStorage_logic_sl_0_allocId_value);
  assign _zz_LsuPlugin_logic_translationStorage_logic_sl_0_write_mask = (2'b01 <<< LsuPlugin_logic_translationStorage_logic_sl_0_allocId_value);
  assign _zz_BtbPlugin_logic_ras_mem_stack_port = BtbPlugin_logic_ras_write_payload_data;
  assign _zz_FetchL1Plugin_logic_ways_0_mem_port = {FetchL1Plugin_logic_waysWrite_tag_address,{FetchL1Plugin_logic_waysWrite_tag_error,FetchL1Plugin_logic_waysWrite_tag_loaded}};
  assign _zz_FetchL1Plugin_logic_ways_0_mem_port_1 = FetchL1Plugin_logic_waysWrite_mask[0];
  assign _zz_FetchL1Plugin_logic_ways_1_mem_port = {FetchL1Plugin_logic_waysWrite_tag_address,{FetchL1Plugin_logic_waysWrite_tag_error,FetchL1Plugin_logic_waysWrite_tag_loaded}};
  assign _zz_FetchL1Plugin_logic_ways_1_mem_port_1 = FetchL1Plugin_logic_waysWrite_mask[1];
  assign _zz_GSharePlugin_logic_mem_counter_port = {GSharePlugin_logic_mem_write_payload_data_3,{GSharePlugin_logic_mem_write_payload_data_2,{GSharePlugin_logic_mem_write_payload_data_1,GSharePlugin_logic_mem_write_payload_data_0}}};
  assign _zz_BtbPlugin_logic_mem_port = {{BtbPlugin_logic_onLearn_port_payload_data_1_isPop,{BtbPlugin_logic_onLearn_port_payload_data_1_isPush,{BtbPlugin_logic_onLearn_port_payload_data_1_isBranch,{BtbPlugin_logic_onLearn_port_payload_data_1_pcTarget,{BtbPlugin_logic_onLearn_port_payload_data_1_sliceLow,BtbPlugin_logic_onLearn_port_payload_data_1_hash}}}}},{BtbPlugin_logic_onLearn_port_payload_data_0_isPop,{BtbPlugin_logic_onLearn_port_payload_data_0_isPush,{BtbPlugin_logic_onLearn_port_payload_data_0_isBranch,{BtbPlugin_logic_onLearn_port_payload_data_0_pcTarget,{BtbPlugin_logic_onLearn_port_payload_data_0_sliceLow,BtbPlugin_logic_onLearn_port_payload_data_0_hash}}}}}};
  assign _zz_LsuL1Plugin_logic_ways_0_mem_port = {LsuL1Plugin_logic_waysWrite_tag_fault,{LsuL1Plugin_logic_waysWrite_tag_address,LsuL1Plugin_logic_waysWrite_tag_loaded}};
  assign _zz_LsuL1Plugin_logic_ways_0_mem_port_1 = LsuL1Plugin_logic_waysWrite_mask[0];
  assign _zz_LsuL1Plugin_logic_ways_1_mem_port = {LsuL1Plugin_logic_waysWrite_tag_fault,{LsuL1Plugin_logic_waysWrite_tag_address,LsuL1Plugin_logic_waysWrite_tag_loaded}};
  assign _zz_LsuL1Plugin_logic_ways_1_mem_port_1 = LsuL1Plugin_logic_waysWrite_mask[1];
  assign _zz_LsuL1Plugin_logic_shared_mem_port = {LsuL1Plugin_logic_shared_write_payload_data_dirty,LsuL1Plugin_logic_shared_write_payload_data_plru_0};
  assign _zz_LsuL1Plugin_logic_writeback_victimBuffer_port = LsuL1Plugin_logic_writeback_read_slotReadLast_payload_wordIndex;
  assign _zz_FetchL1Plugin_logic_translationStorage_logic_sl_0_ways_0_port = {FetchL1Plugin_logic_translationStorage_logic_sl_0_write_data_allowUser,{FetchL1Plugin_logic_translationStorage_logic_sl_0_write_data_allowExecute,{FetchL1Plugin_logic_translationStorage_logic_sl_0_write_data_allowWrite,{FetchL1Plugin_logic_translationStorage_logic_sl_0_write_data_allowRead,{FetchL1Plugin_logic_translationStorage_logic_sl_0_write_data_physicalAddress,{FetchL1Plugin_logic_translationStorage_logic_sl_0_write_data_virtualAddress,FetchL1Plugin_logic_translationStorage_logic_sl_0_write_data_valid}}}}}};
  assign _zz_FetchL1Plugin_logic_translationStorage_logic_sl_0_ways_0_port_1 = FetchL1Plugin_logic_translationStorage_logic_sl_0_write_mask[0];
  assign _zz_FetchL1Plugin_logic_translationStorage_logic_sl_0_ways_1_port = {FetchL1Plugin_logic_translationStorage_logic_sl_0_write_data_allowUser,{FetchL1Plugin_logic_translationStorage_logic_sl_0_write_data_allowExecute,{FetchL1Plugin_logic_translationStorage_logic_sl_0_write_data_allowWrite,{FetchL1Plugin_logic_translationStorage_logic_sl_0_write_data_allowRead,{FetchL1Plugin_logic_translationStorage_logic_sl_0_write_data_physicalAddress,{FetchL1Plugin_logic_translationStorage_logic_sl_0_write_data_virtualAddress,FetchL1Plugin_logic_translationStorage_logic_sl_0_write_data_valid}}}}}};
  assign _zz_FetchL1Plugin_logic_translationStorage_logic_sl_0_ways_1_port_1 = FetchL1Plugin_logic_translationStorage_logic_sl_0_write_mask[1];
  assign _zz_FetchL1Plugin_logic_translationStorage_logic_sl_1_ways_0_port = {FetchL1Plugin_logic_translationStorage_logic_sl_1_write_data_allowUser,{FetchL1Plugin_logic_translationStorage_logic_sl_1_write_data_allowExecute,{FetchL1Plugin_logic_translationStorage_logic_sl_1_write_data_allowWrite,{FetchL1Plugin_logic_translationStorage_logic_sl_1_write_data_allowRead,{FetchL1Plugin_logic_translationStorage_logic_sl_1_write_data_physicalAddress,{FetchL1Plugin_logic_translationStorage_logic_sl_1_write_data_virtualAddress,FetchL1Plugin_logic_translationStorage_logic_sl_1_write_data_valid}}}}}};
  assign _zz_FetchL1Plugin_logic_translationStorage_logic_sl_1_ways_0_port_1 = FetchL1Plugin_logic_translationStorage_logic_sl_1_write_mask[0];
  assign _zz_LsuPlugin_logic_translationStorage_logic_sl_0_ways_0_port = {LsuPlugin_logic_translationStorage_logic_sl_0_write_data_allowUser,{LsuPlugin_logic_translationStorage_logic_sl_0_write_data_allowExecute,{LsuPlugin_logic_translationStorage_logic_sl_0_write_data_allowWrite,{LsuPlugin_logic_translationStorage_logic_sl_0_write_data_allowRead,{LsuPlugin_logic_translationStorage_logic_sl_0_write_data_physicalAddress,{LsuPlugin_logic_translationStorage_logic_sl_0_write_data_virtualAddress,LsuPlugin_logic_translationStorage_logic_sl_0_write_data_valid}}}}}};
  assign _zz_LsuPlugin_logic_translationStorage_logic_sl_0_ways_0_port_1 = LsuPlugin_logic_translationStorage_logic_sl_0_write_mask[0];
  assign _zz_LsuPlugin_logic_translationStorage_logic_sl_0_ways_1_port = {LsuPlugin_logic_translationStorage_logic_sl_0_write_data_allowUser,{LsuPlugin_logic_translationStorage_logic_sl_0_write_data_allowExecute,{LsuPlugin_logic_translationStorage_logic_sl_0_write_data_allowWrite,{LsuPlugin_logic_translationStorage_logic_sl_0_write_data_allowRead,{LsuPlugin_logic_translationStorage_logic_sl_0_write_data_physicalAddress,{LsuPlugin_logic_translationStorage_logic_sl_0_write_data_virtualAddress,LsuPlugin_logic_translationStorage_logic_sl_0_write_data_valid}}}}}};
  assign _zz_LsuPlugin_logic_translationStorage_logic_sl_0_ways_1_port_1 = LsuPlugin_logic_translationStorage_logic_sl_0_write_mask[1];
  assign _zz_LsuPlugin_logic_translationStorage_logic_sl_1_ways_0_port = {LsuPlugin_logic_translationStorage_logic_sl_1_write_data_allowUser,{LsuPlugin_logic_translationStorage_logic_sl_1_write_data_allowExecute,{LsuPlugin_logic_translationStorage_logic_sl_1_write_data_allowWrite,{LsuPlugin_logic_translationStorage_logic_sl_1_write_data_allowRead,{LsuPlugin_logic_translationStorage_logic_sl_1_write_data_physicalAddress,{LsuPlugin_logic_translationStorage_logic_sl_1_write_data_virtualAddress,LsuPlugin_logic_translationStorage_logic_sl_1_write_data_valid}}}}}};
  assign _zz_LsuPlugin_logic_translationStorage_logic_sl_1_ways_0_port_1 = LsuPlugin_logic_translationStorage_logic_sl_1_write_mask[0];
  assign _zz_fetch_logic_ctrls_2_down_AlignerPlugin_logic_FETCH_MASK_1 = fetch_logic_ctrls_2_down_Fetch_WORD_PC[2 : 1];
  assign _zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_28 = AlignerPlugin_logic_extractors_0_ctx_instruction[11 : 10];
  assign _zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_30 = {AlignerPlugin_logic_extractors_0_ctx_instruction[12],AlignerPlugin_logic_extractors_0_ctx_instruction[6 : 5]};
  assign _zz_AlignerPlugin_logic_feeder_lanes_1_withRvc_dec_inst_28 = AlignerPlugin_logic_extractors_1_ctx_instruction[11 : 10];
  assign _zz_AlignerPlugin_logic_feeder_lanes_1_withRvc_dec_inst_30 = {AlignerPlugin_logic_extractors_1_ctx_instruction[12],AlignerPlugin_logic_extractors_1_ctx_instruction[6 : 5]};
  assign _zz_DispatchPlugin_logic_candidates_1_age_1 = (DispatchPlugin_logic_candidates_0_ctx_valid && 1'b1);
  assign _zz_DispatchPlugin_logic_candidates_2_age_1 = {(DispatchPlugin_logic_candidates_1_ctx_valid && 1'b1),(DispatchPlugin_logic_candidates_0_ctx_valid && 1'b1)};
  assign _zz_DispatchPlugin_logic_slotsFeeds_fit_1 = {(! DispatchPlugin_logic_candidates_2_moving),(! DispatchPlugin_logic_candidates_1_moving)};
  assign _zz_toplevel_execute_ctrl3_down_LsuL1Plugin_logic_BANKS_MUXES_lane0_0_1 = toplevel_execute_ctrl3_down_LsuL1_MIXED_ADDRESS_lane0[2 : 2];
  assign _zz_toplevel_execute_ctrl3_down_LsuL1Plugin_logic_BANKS_MUXES_lane0_1_1 = toplevel_execute_ctrl3_down_LsuL1_MIXED_ADDRESS_lane0[2 : 2];
  assign _zz_56 = {_zz_toplevel_execute_ctrl4_down_LsuL1Plugin_logic_MUXED_DATA_lane0_1,_zz_toplevel_execute_ctrl4_down_LsuL1Plugin_logic_MUXED_DATA_lane0};
  assign _zz_58 = {_zz_38[2],{_zz_38[1],_zz_38[0]}};
  assign _zz_LsuPlugin_logic_onCtrl_loadData_shited_1 = toplevel_execute_ctrl4_down_LsuL1_MIXED_ADDRESS_lane0[1 : 0];
  assign _zz_LsuPlugin_logic_onCtrl_loadData_shited_3 = toplevel_execute_ctrl4_down_LsuL1_MIXED_ADDRESS_lane0[1 : 1];
  assign _zz_WhiteboxerPlugin_logic_perf_candidatesCount_1 = {DispatchPlugin_logic_candidates_2_ctx_valid,{DispatchPlugin_logic_candidates_1_ctx_valid,DispatchPlugin_logic_candidates_0_ctx_valid}};
  assign _zz_WhiteboxerPlugin_logic_perf_dispatchFeedCount_1 = {toplevel_decode_ctrls_1_up_LANE_SEL_1,toplevel_decode_ctrls_1_up_LANE_SEL_0};
  assign _zz_early0_BarrelShifterPlugin_logic_shift_reversed_1 = toplevel_execute_ctrl2_down_early0_SrcPlugin_SRC1_lane0[9];
  assign _zz_early0_BarrelShifterPlugin_logic_shift_reversed_2 = toplevel_execute_ctrl2_down_early0_SrcPlugin_SRC1_lane0[10];
  assign _zz_early0_BarrelShifterPlugin_logic_shift_reversed_3 = {toplevel_execute_ctrl2_down_early0_SrcPlugin_SRC1_lane0[11],{toplevel_execute_ctrl2_down_early0_SrcPlugin_SRC1_lane0[12],{toplevel_execute_ctrl2_down_early0_SrcPlugin_SRC1_lane0[13],{toplevel_execute_ctrl2_down_early0_SrcPlugin_SRC1_lane0[14],{toplevel_execute_ctrl2_down_early0_SrcPlugin_SRC1_lane0[15],{toplevel_execute_ctrl2_down_early0_SrcPlugin_SRC1_lane0[16],{toplevel_execute_ctrl2_down_early0_SrcPlugin_SRC1_lane0[17],{toplevel_execute_ctrl2_down_early0_SrcPlugin_SRC1_lane0[18],{toplevel_execute_ctrl2_down_early0_SrcPlugin_SRC1_lane0[19],{_zz_early0_BarrelShifterPlugin_logic_shift_reversed_4,{_zz_early0_BarrelShifterPlugin_logic_shift_reversed_5,_zz_early0_BarrelShifterPlugin_logic_shift_reversed_6}}}}}}}}}}};
  assign _zz_early0_BarrelShifterPlugin_logic_shift_reversed_4 = toplevel_execute_ctrl2_down_early0_SrcPlugin_SRC1_lane0[20];
  assign _zz_early0_BarrelShifterPlugin_logic_shift_reversed_5 = toplevel_execute_ctrl2_down_early0_SrcPlugin_SRC1_lane0[21];
  assign _zz_early0_BarrelShifterPlugin_logic_shift_reversed_6 = {toplevel_execute_ctrl2_down_early0_SrcPlugin_SRC1_lane0[22],{toplevel_execute_ctrl2_down_early0_SrcPlugin_SRC1_lane0[23],{toplevel_execute_ctrl2_down_early0_SrcPlugin_SRC1_lane0[24],{toplevel_execute_ctrl2_down_early0_SrcPlugin_SRC1_lane0[25],{toplevel_execute_ctrl2_down_early0_SrcPlugin_SRC1_lane0[26],{toplevel_execute_ctrl2_down_early0_SrcPlugin_SRC1_lane0[27],{toplevel_execute_ctrl2_down_early0_SrcPlugin_SRC1_lane0[28],{toplevel_execute_ctrl2_down_early0_SrcPlugin_SRC1_lane0[29],{toplevel_execute_ctrl2_down_early0_SrcPlugin_SRC1_lane0[30],toplevel_execute_ctrl2_down_early0_SrcPlugin_SRC1_lane0[31]}}}}}}}}};
  assign _zz_early0_BarrelShifterPlugin_logic_shift_patched_1 = early0_BarrelShifterPlugin_logic_shift_shifted[9];
  assign _zz_early0_BarrelShifterPlugin_logic_shift_patched_2 = early0_BarrelShifterPlugin_logic_shift_shifted[10];
  assign _zz_early0_BarrelShifterPlugin_logic_shift_patched_3 = {early0_BarrelShifterPlugin_logic_shift_shifted[11],{early0_BarrelShifterPlugin_logic_shift_shifted[12],{early0_BarrelShifterPlugin_logic_shift_shifted[13],{early0_BarrelShifterPlugin_logic_shift_shifted[14],{early0_BarrelShifterPlugin_logic_shift_shifted[15],{early0_BarrelShifterPlugin_logic_shift_shifted[16],{early0_BarrelShifterPlugin_logic_shift_shifted[17],{early0_BarrelShifterPlugin_logic_shift_shifted[18],{early0_BarrelShifterPlugin_logic_shift_shifted[19],{_zz_early0_BarrelShifterPlugin_logic_shift_patched_4,{_zz_early0_BarrelShifterPlugin_logic_shift_patched_5,_zz_early0_BarrelShifterPlugin_logic_shift_patched_6}}}}}}}}}}};
  assign _zz_early0_BarrelShifterPlugin_logic_shift_patched_4 = early0_BarrelShifterPlugin_logic_shift_shifted[20];
  assign _zz_early0_BarrelShifterPlugin_logic_shift_patched_5 = early0_BarrelShifterPlugin_logic_shift_shifted[21];
  assign _zz_early0_BarrelShifterPlugin_logic_shift_patched_6 = {early0_BarrelShifterPlugin_logic_shift_shifted[22],{early0_BarrelShifterPlugin_logic_shift_shifted[23],{early0_BarrelShifterPlugin_logic_shift_shifted[24],{early0_BarrelShifterPlugin_logic_shift_shifted[25],{early0_BarrelShifterPlugin_logic_shift_shifted[26],{early0_BarrelShifterPlugin_logic_shift_shifted[27],{early0_BarrelShifterPlugin_logic_shift_shifted[28],{early0_BarrelShifterPlugin_logic_shift_shifted[29],{early0_BarrelShifterPlugin_logic_shift_shifted[30],early0_BarrelShifterPlugin_logic_shift_shifted[31]}}}}}}}}};
  assign _zz_late0_BarrelShifterPlugin_logic_shift_reversed_1 = toplevel_execute_ctrl4_down_late0_SrcPlugin_SRC1_lane0[9];
  assign _zz_late0_BarrelShifterPlugin_logic_shift_reversed_2 = toplevel_execute_ctrl4_down_late0_SrcPlugin_SRC1_lane0[10];
  assign _zz_late0_BarrelShifterPlugin_logic_shift_reversed_3 = {toplevel_execute_ctrl4_down_late0_SrcPlugin_SRC1_lane0[11],{toplevel_execute_ctrl4_down_late0_SrcPlugin_SRC1_lane0[12],{toplevel_execute_ctrl4_down_late0_SrcPlugin_SRC1_lane0[13],{toplevel_execute_ctrl4_down_late0_SrcPlugin_SRC1_lane0[14],{toplevel_execute_ctrl4_down_late0_SrcPlugin_SRC1_lane0[15],{toplevel_execute_ctrl4_down_late0_SrcPlugin_SRC1_lane0[16],{toplevel_execute_ctrl4_down_late0_SrcPlugin_SRC1_lane0[17],{toplevel_execute_ctrl4_down_late0_SrcPlugin_SRC1_lane0[18],{toplevel_execute_ctrl4_down_late0_SrcPlugin_SRC1_lane0[19],{_zz_late0_BarrelShifterPlugin_logic_shift_reversed_4,{_zz_late0_BarrelShifterPlugin_logic_shift_reversed_5,_zz_late0_BarrelShifterPlugin_logic_shift_reversed_6}}}}}}}}}}};
  assign _zz_late0_BarrelShifterPlugin_logic_shift_reversed_4 = toplevel_execute_ctrl4_down_late0_SrcPlugin_SRC1_lane0[20];
  assign _zz_late0_BarrelShifterPlugin_logic_shift_reversed_5 = toplevel_execute_ctrl4_down_late0_SrcPlugin_SRC1_lane0[21];
  assign _zz_late0_BarrelShifterPlugin_logic_shift_reversed_6 = {toplevel_execute_ctrl4_down_late0_SrcPlugin_SRC1_lane0[22],{toplevel_execute_ctrl4_down_late0_SrcPlugin_SRC1_lane0[23],{toplevel_execute_ctrl4_down_late0_SrcPlugin_SRC1_lane0[24],{toplevel_execute_ctrl4_down_late0_SrcPlugin_SRC1_lane0[25],{toplevel_execute_ctrl4_down_late0_SrcPlugin_SRC1_lane0[26],{toplevel_execute_ctrl4_down_late0_SrcPlugin_SRC1_lane0[27],{toplevel_execute_ctrl4_down_late0_SrcPlugin_SRC1_lane0[28],{toplevel_execute_ctrl4_down_late0_SrcPlugin_SRC1_lane0[29],{toplevel_execute_ctrl4_down_late0_SrcPlugin_SRC1_lane0[30],toplevel_execute_ctrl4_down_late0_SrcPlugin_SRC1_lane0[31]}}}}}}}}};
  assign _zz_late0_BarrelShifterPlugin_logic_shift_patched_1 = late0_BarrelShifterPlugin_logic_shift_shifted[9];
  assign _zz_late0_BarrelShifterPlugin_logic_shift_patched_2 = late0_BarrelShifterPlugin_logic_shift_shifted[10];
  assign _zz_late0_BarrelShifterPlugin_logic_shift_patched_3 = {late0_BarrelShifterPlugin_logic_shift_shifted[11],{late0_BarrelShifterPlugin_logic_shift_shifted[12],{late0_BarrelShifterPlugin_logic_shift_shifted[13],{late0_BarrelShifterPlugin_logic_shift_shifted[14],{late0_BarrelShifterPlugin_logic_shift_shifted[15],{late0_BarrelShifterPlugin_logic_shift_shifted[16],{late0_BarrelShifterPlugin_logic_shift_shifted[17],{late0_BarrelShifterPlugin_logic_shift_shifted[18],{late0_BarrelShifterPlugin_logic_shift_shifted[19],{_zz_late0_BarrelShifterPlugin_logic_shift_patched_4,{_zz_late0_BarrelShifterPlugin_logic_shift_patched_5,_zz_late0_BarrelShifterPlugin_logic_shift_patched_6}}}}}}}}}}};
  assign _zz_late0_BarrelShifterPlugin_logic_shift_patched_4 = late0_BarrelShifterPlugin_logic_shift_shifted[20];
  assign _zz_late0_BarrelShifterPlugin_logic_shift_patched_5 = late0_BarrelShifterPlugin_logic_shift_shifted[21];
  assign _zz_late0_BarrelShifterPlugin_logic_shift_patched_6 = {late0_BarrelShifterPlugin_logic_shift_shifted[22],{late0_BarrelShifterPlugin_logic_shift_shifted[23],{late0_BarrelShifterPlugin_logic_shift_shifted[24],{late0_BarrelShifterPlugin_logic_shift_shifted[25],{late0_BarrelShifterPlugin_logic_shift_shifted[26],{late0_BarrelShifterPlugin_logic_shift_shifted[27],{late0_BarrelShifterPlugin_logic_shift_shifted[28],{late0_BarrelShifterPlugin_logic_shift_shifted[29],{late0_BarrelShifterPlugin_logic_shift_shifted[30],late0_BarrelShifterPlugin_logic_shift_shifted[31]}}}}}}}}};
  assign _zz_early1_BarrelShifterPlugin_logic_shift_reversed_1 = toplevel_execute_ctrl2_down_early1_SrcPlugin_SRC1_lane1[9];
  assign _zz_early1_BarrelShifterPlugin_logic_shift_reversed_2 = toplevel_execute_ctrl2_down_early1_SrcPlugin_SRC1_lane1[10];
  assign _zz_early1_BarrelShifterPlugin_logic_shift_reversed_3 = {toplevel_execute_ctrl2_down_early1_SrcPlugin_SRC1_lane1[11],{toplevel_execute_ctrl2_down_early1_SrcPlugin_SRC1_lane1[12],{toplevel_execute_ctrl2_down_early1_SrcPlugin_SRC1_lane1[13],{toplevel_execute_ctrl2_down_early1_SrcPlugin_SRC1_lane1[14],{toplevel_execute_ctrl2_down_early1_SrcPlugin_SRC1_lane1[15],{toplevel_execute_ctrl2_down_early1_SrcPlugin_SRC1_lane1[16],{toplevel_execute_ctrl2_down_early1_SrcPlugin_SRC1_lane1[17],{toplevel_execute_ctrl2_down_early1_SrcPlugin_SRC1_lane1[18],{toplevel_execute_ctrl2_down_early1_SrcPlugin_SRC1_lane1[19],{_zz_early1_BarrelShifterPlugin_logic_shift_reversed_4,{_zz_early1_BarrelShifterPlugin_logic_shift_reversed_5,_zz_early1_BarrelShifterPlugin_logic_shift_reversed_6}}}}}}}}}}};
  assign _zz_early1_BarrelShifterPlugin_logic_shift_reversed_4 = toplevel_execute_ctrl2_down_early1_SrcPlugin_SRC1_lane1[20];
  assign _zz_early1_BarrelShifterPlugin_logic_shift_reversed_5 = toplevel_execute_ctrl2_down_early1_SrcPlugin_SRC1_lane1[21];
  assign _zz_early1_BarrelShifterPlugin_logic_shift_reversed_6 = {toplevel_execute_ctrl2_down_early1_SrcPlugin_SRC1_lane1[22],{toplevel_execute_ctrl2_down_early1_SrcPlugin_SRC1_lane1[23],{toplevel_execute_ctrl2_down_early1_SrcPlugin_SRC1_lane1[24],{toplevel_execute_ctrl2_down_early1_SrcPlugin_SRC1_lane1[25],{toplevel_execute_ctrl2_down_early1_SrcPlugin_SRC1_lane1[26],{toplevel_execute_ctrl2_down_early1_SrcPlugin_SRC1_lane1[27],{toplevel_execute_ctrl2_down_early1_SrcPlugin_SRC1_lane1[28],{toplevel_execute_ctrl2_down_early1_SrcPlugin_SRC1_lane1[29],{toplevel_execute_ctrl2_down_early1_SrcPlugin_SRC1_lane1[30],toplevel_execute_ctrl2_down_early1_SrcPlugin_SRC1_lane1[31]}}}}}}}}};
  assign _zz_early1_BarrelShifterPlugin_logic_shift_patched_1 = early1_BarrelShifterPlugin_logic_shift_shifted[9];
  assign _zz_early1_BarrelShifterPlugin_logic_shift_patched_2 = early1_BarrelShifterPlugin_logic_shift_shifted[10];
  assign _zz_early1_BarrelShifterPlugin_logic_shift_patched_3 = {early1_BarrelShifterPlugin_logic_shift_shifted[11],{early1_BarrelShifterPlugin_logic_shift_shifted[12],{early1_BarrelShifterPlugin_logic_shift_shifted[13],{early1_BarrelShifterPlugin_logic_shift_shifted[14],{early1_BarrelShifterPlugin_logic_shift_shifted[15],{early1_BarrelShifterPlugin_logic_shift_shifted[16],{early1_BarrelShifterPlugin_logic_shift_shifted[17],{early1_BarrelShifterPlugin_logic_shift_shifted[18],{early1_BarrelShifterPlugin_logic_shift_shifted[19],{_zz_early1_BarrelShifterPlugin_logic_shift_patched_4,{_zz_early1_BarrelShifterPlugin_logic_shift_patched_5,_zz_early1_BarrelShifterPlugin_logic_shift_patched_6}}}}}}}}}}};
  assign _zz_early1_BarrelShifterPlugin_logic_shift_patched_4 = early1_BarrelShifterPlugin_logic_shift_shifted[20];
  assign _zz_early1_BarrelShifterPlugin_logic_shift_patched_5 = early1_BarrelShifterPlugin_logic_shift_shifted[21];
  assign _zz_early1_BarrelShifterPlugin_logic_shift_patched_6 = {early1_BarrelShifterPlugin_logic_shift_shifted[22],{early1_BarrelShifterPlugin_logic_shift_shifted[23],{early1_BarrelShifterPlugin_logic_shift_shifted[24],{early1_BarrelShifterPlugin_logic_shift_shifted[25],{early1_BarrelShifterPlugin_logic_shift_shifted[26],{early1_BarrelShifterPlugin_logic_shift_shifted[27],{early1_BarrelShifterPlugin_logic_shift_shifted[28],{early1_BarrelShifterPlugin_logic_shift_shifted[29],{early1_BarrelShifterPlugin_logic_shift_shifted[30],early1_BarrelShifterPlugin_logic_shift_shifted[31]}}}}}}}}};
  assign _zz_late1_BarrelShifterPlugin_logic_shift_reversed_1 = toplevel_execute_ctrl4_down_late1_SrcPlugin_SRC1_lane1[9];
  assign _zz_late1_BarrelShifterPlugin_logic_shift_reversed_2 = toplevel_execute_ctrl4_down_late1_SrcPlugin_SRC1_lane1[10];
  assign _zz_late1_BarrelShifterPlugin_logic_shift_reversed_3 = {toplevel_execute_ctrl4_down_late1_SrcPlugin_SRC1_lane1[11],{toplevel_execute_ctrl4_down_late1_SrcPlugin_SRC1_lane1[12],{toplevel_execute_ctrl4_down_late1_SrcPlugin_SRC1_lane1[13],{toplevel_execute_ctrl4_down_late1_SrcPlugin_SRC1_lane1[14],{toplevel_execute_ctrl4_down_late1_SrcPlugin_SRC1_lane1[15],{toplevel_execute_ctrl4_down_late1_SrcPlugin_SRC1_lane1[16],{toplevel_execute_ctrl4_down_late1_SrcPlugin_SRC1_lane1[17],{toplevel_execute_ctrl4_down_late1_SrcPlugin_SRC1_lane1[18],{toplevel_execute_ctrl4_down_late1_SrcPlugin_SRC1_lane1[19],{_zz_late1_BarrelShifterPlugin_logic_shift_reversed_4,{_zz_late1_BarrelShifterPlugin_logic_shift_reversed_5,_zz_late1_BarrelShifterPlugin_logic_shift_reversed_6}}}}}}}}}}};
  assign _zz_late1_BarrelShifterPlugin_logic_shift_reversed_4 = toplevel_execute_ctrl4_down_late1_SrcPlugin_SRC1_lane1[20];
  assign _zz_late1_BarrelShifterPlugin_logic_shift_reversed_5 = toplevel_execute_ctrl4_down_late1_SrcPlugin_SRC1_lane1[21];
  assign _zz_late1_BarrelShifterPlugin_logic_shift_reversed_6 = {toplevel_execute_ctrl4_down_late1_SrcPlugin_SRC1_lane1[22],{toplevel_execute_ctrl4_down_late1_SrcPlugin_SRC1_lane1[23],{toplevel_execute_ctrl4_down_late1_SrcPlugin_SRC1_lane1[24],{toplevel_execute_ctrl4_down_late1_SrcPlugin_SRC1_lane1[25],{toplevel_execute_ctrl4_down_late1_SrcPlugin_SRC1_lane1[26],{toplevel_execute_ctrl4_down_late1_SrcPlugin_SRC1_lane1[27],{toplevel_execute_ctrl4_down_late1_SrcPlugin_SRC1_lane1[28],{toplevel_execute_ctrl4_down_late1_SrcPlugin_SRC1_lane1[29],{toplevel_execute_ctrl4_down_late1_SrcPlugin_SRC1_lane1[30],toplevel_execute_ctrl4_down_late1_SrcPlugin_SRC1_lane1[31]}}}}}}}}};
  assign _zz_late1_BarrelShifterPlugin_logic_shift_patched_1 = late1_BarrelShifterPlugin_logic_shift_shifted[9];
  assign _zz_late1_BarrelShifterPlugin_logic_shift_patched_2 = late1_BarrelShifterPlugin_logic_shift_shifted[10];
  assign _zz_late1_BarrelShifterPlugin_logic_shift_patched_3 = {late1_BarrelShifterPlugin_logic_shift_shifted[11],{late1_BarrelShifterPlugin_logic_shift_shifted[12],{late1_BarrelShifterPlugin_logic_shift_shifted[13],{late1_BarrelShifterPlugin_logic_shift_shifted[14],{late1_BarrelShifterPlugin_logic_shift_shifted[15],{late1_BarrelShifterPlugin_logic_shift_shifted[16],{late1_BarrelShifterPlugin_logic_shift_shifted[17],{late1_BarrelShifterPlugin_logic_shift_shifted[18],{late1_BarrelShifterPlugin_logic_shift_shifted[19],{_zz_late1_BarrelShifterPlugin_logic_shift_patched_4,{_zz_late1_BarrelShifterPlugin_logic_shift_patched_5,_zz_late1_BarrelShifterPlugin_logic_shift_patched_6}}}}}}}}}}};
  assign _zz_late1_BarrelShifterPlugin_logic_shift_patched_4 = late1_BarrelShifterPlugin_logic_shift_shifted[20];
  assign _zz_late1_BarrelShifterPlugin_logic_shift_patched_5 = late1_BarrelShifterPlugin_logic_shift_shifted[21];
  assign _zz_late1_BarrelShifterPlugin_logic_shift_patched_6 = {late1_BarrelShifterPlugin_logic_shift_shifted[22],{late1_BarrelShifterPlugin_logic_shift_shifted[23],{late1_BarrelShifterPlugin_logic_shift_shifted[24],{late1_BarrelShifterPlugin_logic_shift_shifted[25],{late1_BarrelShifterPlugin_logic_shift_shifted[26],{late1_BarrelShifterPlugin_logic_shift_shifted[27],{late1_BarrelShifterPlugin_logic_shift_shifted[28],{late1_BarrelShifterPlugin_logic_shift_shifted[29],{late1_BarrelShifterPlugin_logic_shift_shifted[30],late1_BarrelShifterPlugin_logic_shift_shifted[31]}}}}}}}}};
  assign _zz_AlignerPlugin_logic_extractors_0_usableMask = AlignerPlugin_logic_usedMask_0[4];
  assign _zz_AlignerPlugin_logic_extractors_0_usableMask_1 = (! AlignerPlugin_logic_usedMask_0[3]);
  assign _zz_AlignerPlugin_logic_extractors_0_usableMask_2 = (AlignerPlugin_logic_scanners_2_valid && (! AlignerPlugin_logic_usedMask_0[2]));
  assign _zz_AlignerPlugin_logic_extractors_0_usableMask_3 = (AlignerPlugin_logic_scanners_1_valid && (! AlignerPlugin_logic_usedMask_0[1]));
  assign _zz_AlignerPlugin_logic_extractors_0_usableMask_4 = (AlignerPlugin_logic_scanners_0_valid && (! AlignerPlugin_logic_usedMask_0[0]));
  assign _zz_AlignerPlugin_logic_extractors_0_redo_9 = AlignerPlugin_logic_scanners_0_redo;
  assign _zz_AlignerPlugin_logic_extractors_0_redo_10 = 1'b0;
  assign _zz_AlignerPlugin_logic_extractors_0_redo_11 = AlignerPlugin_logic_scanners_1_redo;
  assign _zz_AlignerPlugin_logic_extractors_0_redo_12 = 1'b0;
  assign _zz_AlignerPlugin_logic_extractors_0_redo_13 = AlignerPlugin_logic_scanners_2_redo;
  assign _zz_AlignerPlugin_logic_extractors_0_redo_14 = 1'b0;
  assign _zz_AlignerPlugin_logic_extractors_0_redo_15 = AlignerPlugin_logic_scanners_3_redo;
  assign _zz_AlignerPlugin_logic_extractors_0_redo_16 = 1'b0;
  assign _zz_AlignerPlugin_logic_extractors_0_redo_17 = AlignerPlugin_logic_scanners_4_redo;
  assign _zz_AlignerPlugin_logic_extractors_0_redo_18 = 1'b0;
  assign _zz_AlignerPlugin_logic_extractors_0_redo_19 = AlignerPlugin_logic_scanners_5_redo;
  assign _zz_AlignerPlugin_logic_extractors_0_redo_20 = 1'b0;
  assign _zz_AlignerPlugin_logic_extractors_0_redo_21 = AlignerPlugin_logic_scanners_6_redo;
  assign _zz_AlignerPlugin_logic_extractors_0_redo_22 = 1'b0;
  assign _zz_AlignerPlugin_logic_extractors_0_redo_23 = AlignerPlugin_logic_scanners_7_redo;
  assign _zz_AlignerPlugin_logic_extractors_0_redo_24 = 1'b0;
  assign _zz_AlignerPlugin_logic_extractors_0_localMask = AlignerPlugin_logic_scanners_0_checker_1_required;
  assign _zz_AlignerPlugin_logic_extractors_0_localMask_1 = AlignerPlugin_logic_scanners_0_checker_0_required;
  assign _zz_AlignerPlugin_logic_extractors_0_localMask_2 = AlignerPlugin_logic_scanners_1_checker_1_required;
  assign _zz_AlignerPlugin_logic_extractors_0_localMask_3 = AlignerPlugin_logic_scanners_1_checker_0_required;
  assign _zz_AlignerPlugin_logic_extractors_0_localMask_4 = AlignerPlugin_logic_scanners_2_checker_1_required;
  assign _zz_AlignerPlugin_logic_extractors_0_localMask_5 = AlignerPlugin_logic_scanners_2_checker_0_required;
  assign _zz_AlignerPlugin_logic_extractors_0_localMask_6 = AlignerPlugin_logic_scanners_3_checker_1_required;
  assign _zz_AlignerPlugin_logic_extractors_0_localMask_7 = AlignerPlugin_logic_scanners_3_checker_0_required;
  assign _zz_AlignerPlugin_logic_extractors_0_localMask_8 = AlignerPlugin_logic_scanners_4_checker_1_required;
  assign _zz_AlignerPlugin_logic_extractors_0_localMask_9 = AlignerPlugin_logic_scanners_4_checker_0_required;
  assign _zz_AlignerPlugin_logic_extractors_0_localMask_10 = AlignerPlugin_logic_scanners_5_checker_1_required;
  assign _zz_AlignerPlugin_logic_extractors_0_localMask_11 = AlignerPlugin_logic_scanners_5_checker_0_required;
  assign _zz_AlignerPlugin_logic_extractors_0_localMask_12 = AlignerPlugin_logic_scanners_6_checker_1_required;
  assign _zz_AlignerPlugin_logic_extractors_0_localMask_13 = AlignerPlugin_logic_scanners_6_checker_0_required;
  assign _zz_AlignerPlugin_logic_extractors_0_localMask_14 = AlignerPlugin_logic_scanners_7_checker_1_required;
  assign _zz_AlignerPlugin_logic_extractors_0_localMask_15 = AlignerPlugin_logic_scanners_7_checker_0_required;
  assign _zz_AlignerPlugin_logic_extractors_1_usableMask = AlignerPlugin_logic_usedMask_1[4];
  assign _zz_AlignerPlugin_logic_extractors_1_usableMask_1 = (! AlignerPlugin_logic_usedMask_1[3]);
  assign _zz_AlignerPlugin_logic_extractors_1_usableMask_2 = (AlignerPlugin_logic_scanners_2_valid && (! AlignerPlugin_logic_usedMask_1[2]));
  assign _zz_AlignerPlugin_logic_extractors_1_usableMask_3 = (AlignerPlugin_logic_scanners_1_valid && (! AlignerPlugin_logic_usedMask_1[1]));
  assign _zz_AlignerPlugin_logic_extractors_1_redo_8 = AlignerPlugin_logic_scanners_1_redo;
  assign _zz_AlignerPlugin_logic_extractors_1_redo_9 = 1'b0;
  assign _zz_AlignerPlugin_logic_extractors_1_redo_10 = AlignerPlugin_logic_scanners_2_redo;
  assign _zz_AlignerPlugin_logic_extractors_1_redo_11 = 1'b0;
  assign _zz_AlignerPlugin_logic_extractors_1_redo_12 = AlignerPlugin_logic_scanners_3_redo;
  assign _zz_AlignerPlugin_logic_extractors_1_redo_13 = 1'b0;
  assign _zz_AlignerPlugin_logic_extractors_1_redo_14 = AlignerPlugin_logic_scanners_4_redo;
  assign _zz_AlignerPlugin_logic_extractors_1_redo_15 = 1'b0;
  assign _zz_AlignerPlugin_logic_extractors_1_redo_16 = AlignerPlugin_logic_scanners_5_redo;
  assign _zz_AlignerPlugin_logic_extractors_1_redo_17 = 1'b0;
  assign _zz_AlignerPlugin_logic_extractors_1_redo_18 = AlignerPlugin_logic_scanners_6_redo;
  assign _zz_AlignerPlugin_logic_extractors_1_redo_19 = 1'b0;
  assign _zz_AlignerPlugin_logic_extractors_1_localMask = AlignerPlugin_logic_scanners_1_checker_1_required;
  assign _zz_AlignerPlugin_logic_extractors_1_localMask_1 = AlignerPlugin_logic_scanners_1_checker_0_required;
  assign _zz_AlignerPlugin_logic_extractors_1_localMask_2 = AlignerPlugin_logic_scanners_2_checker_1_required;
  assign _zz_AlignerPlugin_logic_extractors_1_localMask_3 = AlignerPlugin_logic_scanners_2_checker_0_required;
  assign _zz_AlignerPlugin_logic_extractors_1_localMask_4 = AlignerPlugin_logic_scanners_3_checker_1_required;
  assign _zz_AlignerPlugin_logic_extractors_1_localMask_5 = AlignerPlugin_logic_scanners_3_checker_0_required;
  assign _zz_AlignerPlugin_logic_extractors_1_localMask_6 = AlignerPlugin_logic_scanners_4_checker_1_required;
  assign _zz_AlignerPlugin_logic_extractors_1_localMask_7 = AlignerPlugin_logic_scanners_4_checker_0_required;
  assign _zz_AlignerPlugin_logic_extractors_1_localMask_8 = AlignerPlugin_logic_scanners_5_checker_1_required;
  assign _zz_AlignerPlugin_logic_extractors_1_localMask_9 = AlignerPlugin_logic_scanners_5_checker_0_required;
  assign _zz_AlignerPlugin_logic_extractors_1_localMask_10 = AlignerPlugin_logic_scanners_6_checker_1_required;
  assign _zz_AlignerPlugin_logic_extractors_1_localMask_11 = AlignerPlugin_logic_scanners_6_checker_0_required;
  assign _zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_23 = {_zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_12,AlignerPlugin_logic_extractors_0_ctx_instruction[4 : 3]};
  assign _zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_24 = AlignerPlugin_logic_extractors_0_ctx_instruction[5];
  assign _zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_25 = AlignerPlugin_logic_extractors_0_ctx_instruction[2];
  assign _zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_31 = 7'h0;
  assign _zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_32 = AlignerPlugin_logic_extractors_0_ctx_instruction[6 : 2];
  assign _zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_33 = AlignerPlugin_logic_extractors_0_ctx_instruction[12];
  assign _zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_34 = AlignerPlugin_logic_extractors_0_ctx_instruction[11 : 7];
  assign _zz_AlignerPlugin_logic_feeder_lanes_1_withRvc_dec_inst_23 = {_zz_AlignerPlugin_logic_feeder_lanes_1_withRvc_dec_inst_12,AlignerPlugin_logic_extractors_1_ctx_instruction[4 : 3]};
  assign _zz_AlignerPlugin_logic_feeder_lanes_1_withRvc_dec_inst_24 = AlignerPlugin_logic_extractors_1_ctx_instruction[5];
  assign _zz_AlignerPlugin_logic_feeder_lanes_1_withRvc_dec_inst_25 = AlignerPlugin_logic_extractors_1_ctx_instruction[2];
  assign _zz_AlignerPlugin_logic_feeder_lanes_1_withRvc_dec_inst_31 = 7'h0;
  assign _zz_AlignerPlugin_logic_feeder_lanes_1_withRvc_dec_inst_32 = AlignerPlugin_logic_extractors_1_ctx_instruction[6 : 2];
  assign _zz_AlignerPlugin_logic_feeder_lanes_1_withRvc_dec_inst_33 = AlignerPlugin_logic_extractors_1_ctx_instruction[12];
  assign _zz_AlignerPlugin_logic_feeder_lanes_1_withRvc_dec_inst_34 = AlignerPlugin_logic_extractors_1_ctx_instruction[11 : 7];
  assign _zz_fetch_logic_ctrls_0_down_GSharePlugin_logic_HASH_1 = _zz_fetch_logic_ctrls_0_down_GSharePlugin_logic_HASH[6];
  assign _zz_fetch_logic_ctrls_0_down_GSharePlugin_logic_HASH_2 = _zz_fetch_logic_ctrls_0_down_GSharePlugin_logic_HASH[7];
  assign _zz_fetch_logic_ctrls_0_down_GSharePlugin_logic_HASH_3 = {_zz_fetch_logic_ctrls_0_down_GSharePlugin_logic_HASH[8],{_zz_fetch_logic_ctrls_0_down_GSharePlugin_logic_HASH[9],{_zz_fetch_logic_ctrls_0_down_GSharePlugin_logic_HASH[10],_zz_fetch_logic_ctrls_0_down_GSharePlugin_logic_HASH[11]}}};
  assign _zz_GSharePlugin_logic_onLearn_hash_1 = _zz_GSharePlugin_logic_onLearn_hash[6];
  assign _zz_GSharePlugin_logic_onLearn_hash_2 = _zz_GSharePlugin_logic_onLearn_hash[7];
  assign _zz_GSharePlugin_logic_onLearn_hash_3 = {_zz_GSharePlugin_logic_onLearn_hash[8],{_zz_GSharePlugin_logic_onLearn_hash[9],{_zz_GSharePlugin_logic_onLearn_hash[10],_zz_GSharePlugin_logic_onLearn_hash[11]}}};
  assign _zz_toplevel_decode_ctrls_1_down_RD_ENABLE_0_1 = 32'h00002008;
  assign _zz_toplevel_decode_ctrls_1_down_RD_ENABLE_0_2 = (toplevel_decode_ctrls_1_down_Decode_INSTRUCTION_0 & 32'h00000050);
  assign _zz_toplevel_decode_ctrls_1_down_RD_ENABLE_0_3 = 32'h00000010;
  assign _zz_toplevel_decode_ctrls_1_down_RD_ENABLE_0_4 = ((toplevel_decode_ctrls_1_down_Decode_INSTRUCTION_0 & 32'h00000028) == 32'h0);
  assign _zz_toplevel_decode_ctrls_1_down_Decode_LEGAL_0 = 32'h0000107f;
  assign _zz_toplevel_decode_ctrls_1_down_Decode_LEGAL_0_1 = (toplevel_decode_ctrls_1_down_Decode_INSTRUCTION_0 & 32'h0000207f);
  assign _zz_toplevel_decode_ctrls_1_down_Decode_LEGAL_0_2 = 32'h00002073;
  assign _zz_toplevel_decode_ctrls_1_down_Decode_LEGAL_0_3 = ((toplevel_decode_ctrls_1_down_Decode_INSTRUCTION_0 & 32'h0000407f) == 32'h00004063);
  assign _zz_toplevel_decode_ctrls_1_down_Decode_LEGAL_0_4 = ((toplevel_decode_ctrls_1_down_Decode_INSTRUCTION_0 & 32'h0000207f) == 32'h00002013);
  assign _zz_toplevel_decode_ctrls_1_down_Decode_LEGAL_0_5 = {((toplevel_decode_ctrls_1_down_Decode_INSTRUCTION_0 & 32'h0000107f) == 32'h00000013),{((toplevel_decode_ctrls_1_down_Decode_INSTRUCTION_0 & 32'h0000603f) == 32'h00000023),{((toplevel_decode_ctrls_1_down_Decode_INSTRUCTION_0 & _zz_toplevel_decode_ctrls_1_down_Decode_LEGAL_0_6) == 32'h00000003),{(_zz_toplevel_decode_ctrls_1_down_Decode_LEGAL_0_7 == _zz_toplevel_decode_ctrls_1_down_Decode_LEGAL_0_8),{_zz_toplevel_decode_ctrls_1_down_Decode_LEGAL_0_9,{_zz_toplevel_decode_ctrls_1_down_Decode_LEGAL_0_10,_zz_toplevel_decode_ctrls_1_down_Decode_LEGAL_0_11}}}}}};
  assign _zz_toplevel_decode_ctrls_1_down_Decode_LEGAL_0_6 = 32'h0000207f;
  assign _zz_toplevel_decode_ctrls_1_down_Decode_LEGAL_0_7 = (toplevel_decode_ctrls_1_down_Decode_INSTRUCTION_0 & 32'h0000505f);
  assign _zz_toplevel_decode_ctrls_1_down_Decode_LEGAL_0_8 = 32'h00000003;
  assign _zz_toplevel_decode_ctrls_1_down_Decode_LEGAL_0_9 = ((toplevel_decode_ctrls_1_down_Decode_INSTRUCTION_0 & 32'h0000707b) == 32'h00000063);
  assign _zz_toplevel_decode_ctrls_1_down_Decode_LEGAL_0_10 = ((toplevel_decode_ctrls_1_down_Decode_INSTRUCTION_0 & 32'h0000607f) == 32'h0000000f);
  assign _zz_toplevel_decode_ctrls_1_down_Decode_LEGAL_0_11 = {((toplevel_decode_ctrls_1_down_Decode_INSTRUCTION_0 & 32'h1800707f) == 32'h0000202f),{((toplevel_decode_ctrls_1_down_Decode_INSTRUCTION_0 & 32'hfc00007f) == 32'h00000033),{((toplevel_decode_ctrls_1_down_Decode_INSTRUCTION_0 & _zz_toplevel_decode_ctrls_1_down_Decode_LEGAL_0_12) == 32'h0800202f),{(_zz_toplevel_decode_ctrls_1_down_Decode_LEGAL_0_13 == _zz_toplevel_decode_ctrls_1_down_Decode_LEGAL_0_14),{_zz_toplevel_decode_ctrls_1_down_Decode_LEGAL_0_15,{_zz_toplevel_decode_ctrls_1_down_Decode_LEGAL_0_16,_zz_toplevel_decode_ctrls_1_down_Decode_LEGAL_0_17}}}}}};
  assign _zz_toplevel_decode_ctrls_1_down_Decode_LEGAL_0_12 = 32'he800707f;
  assign _zz_toplevel_decode_ctrls_1_down_Decode_LEGAL_0_13 = (toplevel_decode_ctrls_1_down_Decode_INSTRUCTION_0 & 32'hfc00305f);
  assign _zz_toplevel_decode_ctrls_1_down_Decode_LEGAL_0_14 = 32'h00001013;
  assign _zz_toplevel_decode_ctrls_1_down_Decode_LEGAL_0_15 = ((toplevel_decode_ctrls_1_down_Decode_INSTRUCTION_0 & 32'hbc00707f) == 32'h00005013);
  assign _zz_toplevel_decode_ctrls_1_down_Decode_LEGAL_0_16 = ((toplevel_decode_ctrls_1_down_Decode_INSTRUCTION_0 & 32'hbe00707f) == 32'h00005033);
  assign _zz_toplevel_decode_ctrls_1_down_Decode_LEGAL_0_17 = {((toplevel_decode_ctrls_1_down_Decode_INSTRUCTION_0 & 32'hbe00707f) == 32'h00000033),{((toplevel_decode_ctrls_1_down_Decode_INSTRUCTION_0 & 32'hf9f0707f) == 32'h1000202f),{((toplevel_decode_ctrls_1_down_Decode_INSTRUCTION_0 & _zz_toplevel_decode_ctrls_1_down_Decode_LEGAL_0_18) == 32'h12000073),{(_zz_toplevel_decode_ctrls_1_down_Decode_LEGAL_0_19 == _zz_toplevel_decode_ctrls_1_down_Decode_LEGAL_0_20),{_zz_toplevel_decode_ctrls_1_down_Decode_LEGAL_0_21,_zz_toplevel_decode_ctrls_1_down_Decode_LEGAL_0_22}}}}};
  assign _zz_toplevel_decode_ctrls_1_down_Decode_LEGAL_0_18 = 32'hfe007fff;
  assign _zz_toplevel_decode_ctrls_1_down_Decode_LEGAL_0_19 = (toplevel_decode_ctrls_1_down_Decode_INSTRUCTION_0 & 32'hdfffffff);
  assign _zz_toplevel_decode_ctrls_1_down_Decode_LEGAL_0_20 = 32'h10200073;
  assign _zz_toplevel_decode_ctrls_1_down_Decode_LEGAL_0_21 = ((toplevel_decode_ctrls_1_down_Decode_INSTRUCTION_0 & 32'hffefffff) == 32'h00000073);
  assign _zz_toplevel_decode_ctrls_1_down_Decode_LEGAL_0_22 = ((toplevel_decode_ctrls_1_down_Decode_INSTRUCTION_0 & 32'hffffffff) == 32'h10500073);
  assign _zz_toplevel_decode_ctrls_1_down_RD_ENABLE_1_1 = 32'h00002008;
  assign _zz_toplevel_decode_ctrls_1_down_RD_ENABLE_1_2 = (toplevel_decode_ctrls_1_down_Decode_INSTRUCTION_1 & 32'h00000050);
  assign _zz_toplevel_decode_ctrls_1_down_RD_ENABLE_1_3 = 32'h00000010;
  assign _zz_toplevel_decode_ctrls_1_down_RD_ENABLE_1_4 = ((toplevel_decode_ctrls_1_down_Decode_INSTRUCTION_1 & 32'h00000028) == 32'h0);
  assign _zz_toplevel_decode_ctrls_1_down_Decode_LEGAL_1 = 32'h0000107f;
  assign _zz_toplevel_decode_ctrls_1_down_Decode_LEGAL_1_1 = (toplevel_decode_ctrls_1_down_Decode_INSTRUCTION_1 & 32'h0000207f);
  assign _zz_toplevel_decode_ctrls_1_down_Decode_LEGAL_1_2 = 32'h00002073;
  assign _zz_toplevel_decode_ctrls_1_down_Decode_LEGAL_1_3 = ((toplevel_decode_ctrls_1_down_Decode_INSTRUCTION_1 & 32'h0000407f) == 32'h00004063);
  assign _zz_toplevel_decode_ctrls_1_down_Decode_LEGAL_1_4 = ((toplevel_decode_ctrls_1_down_Decode_INSTRUCTION_1 & 32'h0000207f) == 32'h00002013);
  assign _zz_toplevel_decode_ctrls_1_down_Decode_LEGAL_1_5 = {((toplevel_decode_ctrls_1_down_Decode_INSTRUCTION_1 & 32'h0000107f) == 32'h00000013),{((toplevel_decode_ctrls_1_down_Decode_INSTRUCTION_1 & 32'h0000603f) == 32'h00000023),{((toplevel_decode_ctrls_1_down_Decode_INSTRUCTION_1 & _zz_toplevel_decode_ctrls_1_down_Decode_LEGAL_1_6) == 32'h00000003),{(_zz_toplevel_decode_ctrls_1_down_Decode_LEGAL_1_7 == _zz_toplevel_decode_ctrls_1_down_Decode_LEGAL_1_8),{_zz_toplevel_decode_ctrls_1_down_Decode_LEGAL_1_9,{_zz_toplevel_decode_ctrls_1_down_Decode_LEGAL_1_10,_zz_toplevel_decode_ctrls_1_down_Decode_LEGAL_1_11}}}}}};
  assign _zz_toplevel_decode_ctrls_1_down_Decode_LEGAL_1_6 = 32'h0000207f;
  assign _zz_toplevel_decode_ctrls_1_down_Decode_LEGAL_1_7 = (toplevel_decode_ctrls_1_down_Decode_INSTRUCTION_1 & 32'h0000505f);
  assign _zz_toplevel_decode_ctrls_1_down_Decode_LEGAL_1_8 = 32'h00000003;
  assign _zz_toplevel_decode_ctrls_1_down_Decode_LEGAL_1_9 = ((toplevel_decode_ctrls_1_down_Decode_INSTRUCTION_1 & 32'h0000707b) == 32'h00000063);
  assign _zz_toplevel_decode_ctrls_1_down_Decode_LEGAL_1_10 = ((toplevel_decode_ctrls_1_down_Decode_INSTRUCTION_1 & 32'h0000607f) == 32'h0000000f);
  assign _zz_toplevel_decode_ctrls_1_down_Decode_LEGAL_1_11 = {((toplevel_decode_ctrls_1_down_Decode_INSTRUCTION_1 & 32'h1800707f) == 32'h0000202f),{((toplevel_decode_ctrls_1_down_Decode_INSTRUCTION_1 & 32'hfc00007f) == 32'h00000033),{((toplevel_decode_ctrls_1_down_Decode_INSTRUCTION_1 & _zz_toplevel_decode_ctrls_1_down_Decode_LEGAL_1_12) == 32'h0800202f),{(_zz_toplevel_decode_ctrls_1_down_Decode_LEGAL_1_13 == _zz_toplevel_decode_ctrls_1_down_Decode_LEGAL_1_14),{_zz_toplevel_decode_ctrls_1_down_Decode_LEGAL_1_15,{_zz_toplevel_decode_ctrls_1_down_Decode_LEGAL_1_16,_zz_toplevel_decode_ctrls_1_down_Decode_LEGAL_1_17}}}}}};
  assign _zz_toplevel_decode_ctrls_1_down_Decode_LEGAL_1_12 = 32'he800707f;
  assign _zz_toplevel_decode_ctrls_1_down_Decode_LEGAL_1_13 = (toplevel_decode_ctrls_1_down_Decode_INSTRUCTION_1 & 32'hfc00305f);
  assign _zz_toplevel_decode_ctrls_1_down_Decode_LEGAL_1_14 = 32'h00001013;
  assign _zz_toplevel_decode_ctrls_1_down_Decode_LEGAL_1_15 = ((toplevel_decode_ctrls_1_down_Decode_INSTRUCTION_1 & 32'hbc00707f) == 32'h00005013);
  assign _zz_toplevel_decode_ctrls_1_down_Decode_LEGAL_1_16 = ((toplevel_decode_ctrls_1_down_Decode_INSTRUCTION_1 & 32'hbe00707f) == 32'h00005033);
  assign _zz_toplevel_decode_ctrls_1_down_Decode_LEGAL_1_17 = {((toplevel_decode_ctrls_1_down_Decode_INSTRUCTION_1 & 32'hbe00707f) == 32'h00000033),{((toplevel_decode_ctrls_1_down_Decode_INSTRUCTION_1 & 32'hf9f0707f) == 32'h1000202f),{((toplevel_decode_ctrls_1_down_Decode_INSTRUCTION_1 & _zz_toplevel_decode_ctrls_1_down_Decode_LEGAL_1_18) == 32'h12000073),{(_zz_toplevel_decode_ctrls_1_down_Decode_LEGAL_1_19 == _zz_toplevel_decode_ctrls_1_down_Decode_LEGAL_1_20),{_zz_toplevel_decode_ctrls_1_down_Decode_LEGAL_1_21,_zz_toplevel_decode_ctrls_1_down_Decode_LEGAL_1_22}}}}};
  assign _zz_toplevel_decode_ctrls_1_down_Decode_LEGAL_1_18 = 32'hfe007fff;
  assign _zz_toplevel_decode_ctrls_1_down_Decode_LEGAL_1_19 = (toplevel_decode_ctrls_1_down_Decode_INSTRUCTION_1 & 32'hdfffffff);
  assign _zz_toplevel_decode_ctrls_1_down_Decode_LEGAL_1_20 = 32'h10200073;
  assign _zz_toplevel_decode_ctrls_1_down_Decode_LEGAL_1_21 = ((toplevel_decode_ctrls_1_down_Decode_INSTRUCTION_1 & 32'hffefffff) == 32'h00000073);
  assign _zz_toplevel_decode_ctrls_1_down_Decode_LEGAL_1_22 = ((toplevel_decode_ctrls_1_down_Decode_INSTRUCTION_1 & 32'hffffffff) == 32'h10500073);
  assign _zz_CsrRamPlugin_csrMapper_ramAddress_1 = 12'h002;
  assign _zz_CsrRamPlugin_csrMapper_ramAddress_2 = 12'h040;
  assign _zz_DispatchPlugin_logic_rsHazardChecker_0_onLl_0_onRs_0_hazard = (DispatchPlugin_logic_candidates_0_ctx_hm_DispatchPlugin_logic_hcs_0_onRs_0_ENABLES_0 && toplevel_execute_ctrl1_up_RD_ENABLE_lane1);
  assign _zz_DispatchPlugin_logic_rsHazardChecker_0_onLl_0_onRs_0_hazard_1 = (toplevel_execute_ctrl1_up_RD_PHYS_lane1 == DispatchPlugin_logic_candidates_0_ctx_hm_RS1_PHYS);
  assign _zz_DispatchPlugin_logic_rsHazardChecker_0_onLl_0_onRs_0_hazard_2 = ((DispatchPlugin_logic_candidates_0_ctx_hm_DispatchPlugin_logic_hcs_0_onRs_0_ENABLES_0 && toplevel_execute_ctrl2_up_RD_ENABLE_lane0) && (toplevel_execute_ctrl2_up_RD_PHYS_lane0 == DispatchPlugin_logic_candidates_0_ctx_hm_RS1_PHYS));
  assign _zz_DispatchPlugin_logic_rsHazardChecker_0_onLl_0_onRs_0_hazard_3 = 1'b1;
  assign _zz_DispatchPlugin_logic_rsHazardChecker_0_onLl_0_onRs_0_hazard_4 = ((DispatchPlugin_logic_candidates_0_ctx_hm_DispatchPlugin_logic_hcs_0_onRs_0_ENABLES_0 && toplevel_execute_ctrl1_up_RD_ENABLE_lane0) && (toplevel_execute_ctrl1_up_RD_PHYS_lane0 == DispatchPlugin_logic_candidates_0_ctx_hm_RS1_PHYS));
  assign _zz_DispatchPlugin_logic_rsHazardChecker_0_onLl_0_onRs_0_hazard_5 = 1'b1;
  assign _zz_DispatchPlugin_logic_rsHazardChecker_0_onLl_0_onRs_1_hazard = (DispatchPlugin_logic_candidates_0_ctx_hm_DispatchPlugin_logic_hcs_0_onRs_1_ENABLES_0 && toplevel_execute_ctrl1_up_RD_ENABLE_lane1);
  assign _zz_DispatchPlugin_logic_rsHazardChecker_0_onLl_0_onRs_1_hazard_1 = (toplevel_execute_ctrl1_up_RD_PHYS_lane1 == DispatchPlugin_logic_candidates_0_ctx_hm_RS2_PHYS);
  assign _zz_DispatchPlugin_logic_rsHazardChecker_0_onLl_0_onRs_1_hazard_2 = ((DispatchPlugin_logic_candidates_0_ctx_hm_DispatchPlugin_logic_hcs_0_onRs_1_ENABLES_0 && toplevel_execute_ctrl2_up_RD_ENABLE_lane0) && (toplevel_execute_ctrl2_up_RD_PHYS_lane0 == DispatchPlugin_logic_candidates_0_ctx_hm_RS2_PHYS));
  assign _zz_DispatchPlugin_logic_rsHazardChecker_0_onLl_0_onRs_1_hazard_3 = 1'b1;
  assign _zz_DispatchPlugin_logic_rsHazardChecker_0_onLl_0_onRs_1_hazard_4 = ((DispatchPlugin_logic_candidates_0_ctx_hm_DispatchPlugin_logic_hcs_0_onRs_1_ENABLES_0 && toplevel_execute_ctrl1_up_RD_ENABLE_lane0) && (toplevel_execute_ctrl1_up_RD_PHYS_lane0 == DispatchPlugin_logic_candidates_0_ctx_hm_RS2_PHYS));
  assign _zz_DispatchPlugin_logic_rsHazardChecker_0_onLl_0_onRs_1_hazard_5 = 1'b1;
  assign _zz_DispatchPlugin_logic_rsHazardChecker_0_onLl_1_onRs_0_hazard = (DispatchPlugin_logic_candidates_0_ctx_hm_DispatchPlugin_logic_hcs_1_onRs_0_ENABLES_0 && toplevel_execute_ctrl1_up_RD_ENABLE_lane1);
  assign _zz_DispatchPlugin_logic_rsHazardChecker_0_onLl_1_onRs_0_hazard_1 = (toplevel_execute_ctrl1_up_RD_PHYS_lane1 == DispatchPlugin_logic_candidates_0_ctx_hm_RS1_PHYS);
  assign _zz_DispatchPlugin_logic_rsHazardChecker_0_onLl_1_onRs_0_hazard_2 = ((DispatchPlugin_logic_candidates_0_ctx_hm_DispatchPlugin_logic_hcs_1_onRs_0_ENABLES_0 && toplevel_execute_ctrl2_up_RD_ENABLE_lane0) && (toplevel_execute_ctrl2_up_RD_PHYS_lane0 == DispatchPlugin_logic_candidates_0_ctx_hm_RS1_PHYS));
  assign _zz_DispatchPlugin_logic_rsHazardChecker_0_onLl_1_onRs_0_hazard_3 = 1'b1;
  assign _zz_DispatchPlugin_logic_rsHazardChecker_0_onLl_1_onRs_0_hazard_4 = ((DispatchPlugin_logic_candidates_0_ctx_hm_DispatchPlugin_logic_hcs_1_onRs_0_ENABLES_0 && toplevel_execute_ctrl1_up_RD_ENABLE_lane0) && (toplevel_execute_ctrl1_up_RD_PHYS_lane0 == DispatchPlugin_logic_candidates_0_ctx_hm_RS1_PHYS));
  assign _zz_DispatchPlugin_logic_rsHazardChecker_0_onLl_1_onRs_0_hazard_5 = 1'b1;
  assign _zz_DispatchPlugin_logic_rsHazardChecker_0_onLl_1_onRs_1_hazard = (DispatchPlugin_logic_candidates_0_ctx_hm_DispatchPlugin_logic_hcs_1_onRs_1_ENABLES_0 && toplevel_execute_ctrl1_up_RD_ENABLE_lane1);
  assign _zz_DispatchPlugin_logic_rsHazardChecker_0_onLl_1_onRs_1_hazard_1 = (toplevel_execute_ctrl1_up_RD_PHYS_lane1 == DispatchPlugin_logic_candidates_0_ctx_hm_RS2_PHYS);
  assign _zz_DispatchPlugin_logic_rsHazardChecker_0_onLl_1_onRs_1_hazard_2 = ((DispatchPlugin_logic_candidates_0_ctx_hm_DispatchPlugin_logic_hcs_1_onRs_1_ENABLES_0 && toplevel_execute_ctrl2_up_RD_ENABLE_lane0) && (toplevel_execute_ctrl2_up_RD_PHYS_lane0 == DispatchPlugin_logic_candidates_0_ctx_hm_RS2_PHYS));
  assign _zz_DispatchPlugin_logic_rsHazardChecker_0_onLl_1_onRs_1_hazard_3 = 1'b1;
  assign _zz_DispatchPlugin_logic_rsHazardChecker_0_onLl_1_onRs_1_hazard_4 = ((DispatchPlugin_logic_candidates_0_ctx_hm_DispatchPlugin_logic_hcs_1_onRs_1_ENABLES_0 && toplevel_execute_ctrl1_up_RD_ENABLE_lane0) && (toplevel_execute_ctrl1_up_RD_PHYS_lane0 == DispatchPlugin_logic_candidates_0_ctx_hm_RS2_PHYS));
  assign _zz_DispatchPlugin_logic_rsHazardChecker_0_onLl_1_onRs_1_hazard_5 = 1'b1;
  assign _zz_DispatchPlugin_logic_rsHazardChecker_1_onLl_0_onRs_0_hazard = (DispatchPlugin_logic_candidates_1_ctx_hm_DispatchPlugin_logic_hcs_0_onRs_0_ENABLES_0 && toplevel_execute_ctrl1_up_RD_ENABLE_lane1);
  assign _zz_DispatchPlugin_logic_rsHazardChecker_1_onLl_0_onRs_0_hazard_1 = (toplevel_execute_ctrl1_up_RD_PHYS_lane1 == DispatchPlugin_logic_candidates_1_ctx_hm_RS1_PHYS);
  assign _zz_DispatchPlugin_logic_rsHazardChecker_1_onLl_0_onRs_0_hazard_2 = ((DispatchPlugin_logic_candidates_1_ctx_hm_DispatchPlugin_logic_hcs_0_onRs_0_ENABLES_0 && toplevel_execute_ctrl2_up_RD_ENABLE_lane0) && (toplevel_execute_ctrl2_up_RD_PHYS_lane0 == DispatchPlugin_logic_candidates_1_ctx_hm_RS1_PHYS));
  assign _zz_DispatchPlugin_logic_rsHazardChecker_1_onLl_0_onRs_0_hazard_3 = 1'b1;
  assign _zz_DispatchPlugin_logic_rsHazardChecker_1_onLl_0_onRs_0_hazard_4 = ((DispatchPlugin_logic_candidates_1_ctx_hm_DispatchPlugin_logic_hcs_0_onRs_0_ENABLES_0 && toplevel_execute_ctrl1_up_RD_ENABLE_lane0) && (toplevel_execute_ctrl1_up_RD_PHYS_lane0 == DispatchPlugin_logic_candidates_1_ctx_hm_RS1_PHYS));
  assign _zz_DispatchPlugin_logic_rsHazardChecker_1_onLl_0_onRs_0_hazard_5 = 1'b1;
  assign _zz_DispatchPlugin_logic_rsHazardChecker_1_onLl_0_onRs_1_hazard = (DispatchPlugin_logic_candidates_1_ctx_hm_DispatchPlugin_logic_hcs_0_onRs_1_ENABLES_0 && toplevel_execute_ctrl1_up_RD_ENABLE_lane1);
  assign _zz_DispatchPlugin_logic_rsHazardChecker_1_onLl_0_onRs_1_hazard_1 = (toplevel_execute_ctrl1_up_RD_PHYS_lane1 == DispatchPlugin_logic_candidates_1_ctx_hm_RS2_PHYS);
  assign _zz_DispatchPlugin_logic_rsHazardChecker_1_onLl_0_onRs_1_hazard_2 = ((DispatchPlugin_logic_candidates_1_ctx_hm_DispatchPlugin_logic_hcs_0_onRs_1_ENABLES_0 && toplevel_execute_ctrl2_up_RD_ENABLE_lane0) && (toplevel_execute_ctrl2_up_RD_PHYS_lane0 == DispatchPlugin_logic_candidates_1_ctx_hm_RS2_PHYS));
  assign _zz_DispatchPlugin_logic_rsHazardChecker_1_onLl_0_onRs_1_hazard_3 = 1'b1;
  assign _zz_DispatchPlugin_logic_rsHazardChecker_1_onLl_0_onRs_1_hazard_4 = ((DispatchPlugin_logic_candidates_1_ctx_hm_DispatchPlugin_logic_hcs_0_onRs_1_ENABLES_0 && toplevel_execute_ctrl1_up_RD_ENABLE_lane0) && (toplevel_execute_ctrl1_up_RD_PHYS_lane0 == DispatchPlugin_logic_candidates_1_ctx_hm_RS2_PHYS));
  assign _zz_DispatchPlugin_logic_rsHazardChecker_1_onLl_0_onRs_1_hazard_5 = 1'b1;
  assign _zz_DispatchPlugin_logic_rsHazardChecker_1_onLl_1_onRs_0_hazard = (DispatchPlugin_logic_candidates_1_ctx_hm_DispatchPlugin_logic_hcs_1_onRs_0_ENABLES_0 && toplevel_execute_ctrl1_up_RD_ENABLE_lane1);
  assign _zz_DispatchPlugin_logic_rsHazardChecker_1_onLl_1_onRs_0_hazard_1 = (toplevel_execute_ctrl1_up_RD_PHYS_lane1 == DispatchPlugin_logic_candidates_1_ctx_hm_RS1_PHYS);
  assign _zz_DispatchPlugin_logic_rsHazardChecker_1_onLl_1_onRs_0_hazard_2 = ((DispatchPlugin_logic_candidates_1_ctx_hm_DispatchPlugin_logic_hcs_1_onRs_0_ENABLES_0 && toplevel_execute_ctrl2_up_RD_ENABLE_lane0) && (toplevel_execute_ctrl2_up_RD_PHYS_lane0 == DispatchPlugin_logic_candidates_1_ctx_hm_RS1_PHYS));
  assign _zz_DispatchPlugin_logic_rsHazardChecker_1_onLl_1_onRs_0_hazard_3 = 1'b1;
  assign _zz_DispatchPlugin_logic_rsHazardChecker_1_onLl_1_onRs_0_hazard_4 = ((DispatchPlugin_logic_candidates_1_ctx_hm_DispatchPlugin_logic_hcs_1_onRs_0_ENABLES_0 && toplevel_execute_ctrl1_up_RD_ENABLE_lane0) && (toplevel_execute_ctrl1_up_RD_PHYS_lane0 == DispatchPlugin_logic_candidates_1_ctx_hm_RS1_PHYS));
  assign _zz_DispatchPlugin_logic_rsHazardChecker_1_onLl_1_onRs_0_hazard_5 = 1'b1;
  assign _zz_DispatchPlugin_logic_rsHazardChecker_1_onLl_1_onRs_1_hazard = (DispatchPlugin_logic_candidates_1_ctx_hm_DispatchPlugin_logic_hcs_1_onRs_1_ENABLES_0 && toplevel_execute_ctrl1_up_RD_ENABLE_lane1);
  assign _zz_DispatchPlugin_logic_rsHazardChecker_1_onLl_1_onRs_1_hazard_1 = (toplevel_execute_ctrl1_up_RD_PHYS_lane1 == DispatchPlugin_logic_candidates_1_ctx_hm_RS2_PHYS);
  assign _zz_DispatchPlugin_logic_rsHazardChecker_1_onLl_1_onRs_1_hazard_2 = ((DispatchPlugin_logic_candidates_1_ctx_hm_DispatchPlugin_logic_hcs_1_onRs_1_ENABLES_0 && toplevel_execute_ctrl2_up_RD_ENABLE_lane0) && (toplevel_execute_ctrl2_up_RD_PHYS_lane0 == DispatchPlugin_logic_candidates_1_ctx_hm_RS2_PHYS));
  assign _zz_DispatchPlugin_logic_rsHazardChecker_1_onLl_1_onRs_1_hazard_3 = 1'b1;
  assign _zz_DispatchPlugin_logic_rsHazardChecker_1_onLl_1_onRs_1_hazard_4 = ((DispatchPlugin_logic_candidates_1_ctx_hm_DispatchPlugin_logic_hcs_1_onRs_1_ENABLES_0 && toplevel_execute_ctrl1_up_RD_ENABLE_lane0) && (toplevel_execute_ctrl1_up_RD_PHYS_lane0 == DispatchPlugin_logic_candidates_1_ctx_hm_RS2_PHYS));
  assign _zz_DispatchPlugin_logic_rsHazardChecker_1_onLl_1_onRs_1_hazard_5 = 1'b1;
  assign _zz_DispatchPlugin_logic_rsHazardChecker_2_onLl_0_onRs_0_hazard = (DispatchPlugin_logic_candidates_2_ctx_hm_DispatchPlugin_logic_hcs_0_onRs_0_ENABLES_0 && toplevel_execute_ctrl1_up_RD_ENABLE_lane1);
  assign _zz_DispatchPlugin_logic_rsHazardChecker_2_onLl_0_onRs_0_hazard_1 = (toplevel_execute_ctrl1_up_RD_PHYS_lane1 == DispatchPlugin_logic_candidates_2_ctx_hm_RS1_PHYS);
  assign _zz_DispatchPlugin_logic_rsHazardChecker_2_onLl_0_onRs_0_hazard_2 = ((DispatchPlugin_logic_candidates_2_ctx_hm_DispatchPlugin_logic_hcs_0_onRs_0_ENABLES_0 && toplevel_execute_ctrl2_up_RD_ENABLE_lane0) && (toplevel_execute_ctrl2_up_RD_PHYS_lane0 == DispatchPlugin_logic_candidates_2_ctx_hm_RS1_PHYS));
  assign _zz_DispatchPlugin_logic_rsHazardChecker_2_onLl_0_onRs_0_hazard_3 = 1'b1;
  assign _zz_DispatchPlugin_logic_rsHazardChecker_2_onLl_0_onRs_0_hazard_4 = ((DispatchPlugin_logic_candidates_2_ctx_hm_DispatchPlugin_logic_hcs_0_onRs_0_ENABLES_0 && toplevel_execute_ctrl1_up_RD_ENABLE_lane0) && (toplevel_execute_ctrl1_up_RD_PHYS_lane0 == DispatchPlugin_logic_candidates_2_ctx_hm_RS1_PHYS));
  assign _zz_DispatchPlugin_logic_rsHazardChecker_2_onLl_0_onRs_0_hazard_5 = 1'b1;
  assign _zz_DispatchPlugin_logic_rsHazardChecker_2_onLl_0_onRs_1_hazard = (DispatchPlugin_logic_candidates_2_ctx_hm_DispatchPlugin_logic_hcs_0_onRs_1_ENABLES_0 && toplevel_execute_ctrl1_up_RD_ENABLE_lane1);
  assign _zz_DispatchPlugin_logic_rsHazardChecker_2_onLl_0_onRs_1_hazard_1 = (toplevel_execute_ctrl1_up_RD_PHYS_lane1 == DispatchPlugin_logic_candidates_2_ctx_hm_RS2_PHYS);
  assign _zz_DispatchPlugin_logic_rsHazardChecker_2_onLl_0_onRs_1_hazard_2 = ((DispatchPlugin_logic_candidates_2_ctx_hm_DispatchPlugin_logic_hcs_0_onRs_1_ENABLES_0 && toplevel_execute_ctrl2_up_RD_ENABLE_lane0) && (toplevel_execute_ctrl2_up_RD_PHYS_lane0 == DispatchPlugin_logic_candidates_2_ctx_hm_RS2_PHYS));
  assign _zz_DispatchPlugin_logic_rsHazardChecker_2_onLl_0_onRs_1_hazard_3 = 1'b1;
  assign _zz_DispatchPlugin_logic_rsHazardChecker_2_onLl_0_onRs_1_hazard_4 = ((DispatchPlugin_logic_candidates_2_ctx_hm_DispatchPlugin_logic_hcs_0_onRs_1_ENABLES_0 && toplevel_execute_ctrl1_up_RD_ENABLE_lane0) && (toplevel_execute_ctrl1_up_RD_PHYS_lane0 == DispatchPlugin_logic_candidates_2_ctx_hm_RS2_PHYS));
  assign _zz_DispatchPlugin_logic_rsHazardChecker_2_onLl_0_onRs_1_hazard_5 = 1'b1;
  assign _zz_DispatchPlugin_logic_rsHazardChecker_2_onLl_1_onRs_0_hazard = (DispatchPlugin_logic_candidates_2_ctx_hm_DispatchPlugin_logic_hcs_1_onRs_0_ENABLES_0 && toplevel_execute_ctrl1_up_RD_ENABLE_lane1);
  assign _zz_DispatchPlugin_logic_rsHazardChecker_2_onLl_1_onRs_0_hazard_1 = (toplevel_execute_ctrl1_up_RD_PHYS_lane1 == DispatchPlugin_logic_candidates_2_ctx_hm_RS1_PHYS);
  assign _zz_DispatchPlugin_logic_rsHazardChecker_2_onLl_1_onRs_0_hazard_2 = ((DispatchPlugin_logic_candidates_2_ctx_hm_DispatchPlugin_logic_hcs_1_onRs_0_ENABLES_0 && toplevel_execute_ctrl2_up_RD_ENABLE_lane0) && (toplevel_execute_ctrl2_up_RD_PHYS_lane0 == DispatchPlugin_logic_candidates_2_ctx_hm_RS1_PHYS));
  assign _zz_DispatchPlugin_logic_rsHazardChecker_2_onLl_1_onRs_0_hazard_3 = 1'b1;
  assign _zz_DispatchPlugin_logic_rsHazardChecker_2_onLl_1_onRs_0_hazard_4 = ((DispatchPlugin_logic_candidates_2_ctx_hm_DispatchPlugin_logic_hcs_1_onRs_0_ENABLES_0 && toplevel_execute_ctrl1_up_RD_ENABLE_lane0) && (toplevel_execute_ctrl1_up_RD_PHYS_lane0 == DispatchPlugin_logic_candidates_2_ctx_hm_RS1_PHYS));
  assign _zz_DispatchPlugin_logic_rsHazardChecker_2_onLl_1_onRs_0_hazard_5 = 1'b1;
  assign _zz_DispatchPlugin_logic_rsHazardChecker_2_onLl_1_onRs_1_hazard = (DispatchPlugin_logic_candidates_2_ctx_hm_DispatchPlugin_logic_hcs_1_onRs_1_ENABLES_0 && toplevel_execute_ctrl1_up_RD_ENABLE_lane1);
  assign _zz_DispatchPlugin_logic_rsHazardChecker_2_onLl_1_onRs_1_hazard_1 = (toplevel_execute_ctrl1_up_RD_PHYS_lane1 == DispatchPlugin_logic_candidates_2_ctx_hm_RS2_PHYS);
  assign _zz_DispatchPlugin_logic_rsHazardChecker_2_onLl_1_onRs_1_hazard_2 = ((DispatchPlugin_logic_candidates_2_ctx_hm_DispatchPlugin_logic_hcs_1_onRs_1_ENABLES_0 && toplevel_execute_ctrl2_up_RD_ENABLE_lane0) && (toplevel_execute_ctrl2_up_RD_PHYS_lane0 == DispatchPlugin_logic_candidates_2_ctx_hm_RS2_PHYS));
  assign _zz_DispatchPlugin_logic_rsHazardChecker_2_onLl_1_onRs_1_hazard_3 = 1'b1;
  assign _zz_DispatchPlugin_logic_rsHazardChecker_2_onLl_1_onRs_1_hazard_4 = ((DispatchPlugin_logic_candidates_2_ctx_hm_DispatchPlugin_logic_hcs_1_onRs_1_ENABLES_0 && toplevel_execute_ctrl1_up_RD_ENABLE_lane0) && (toplevel_execute_ctrl1_up_RD_PHYS_lane0 == DispatchPlugin_logic_candidates_2_ctx_hm_RS2_PHYS));
  assign _zz_DispatchPlugin_logic_rsHazardChecker_2_onLl_1_onRs_1_hazard_5 = 1'b1;
  assign _zz__zz_BtbPlugin_logic_applyIt_entry_hash = fetch_logic_ctrls_2_down_BtbPlugin_logic_chunksLogic_0_readRsp_ENTRY_pcTarget;
  assign _zz__zz_BtbPlugin_logic_applyIt_entry_hash_1 = {fetch_logic_ctrls_2_down_BtbPlugin_logic_chunksLogic_0_readRsp_ENTRY_sliceLow,fetch_logic_ctrls_2_down_BtbPlugin_logic_chunksLogic_0_readRsp_ENTRY_hash};
  assign _zz__zz_BtbPlugin_logic_applyIt_entry_hash_2 = fetch_logic_ctrls_2_down_BtbPlugin_logic_chunksLogic_1_readRsp_ENTRY_pcTarget;
  assign _zz__zz_BtbPlugin_logic_applyIt_entry_hash_3 = {fetch_logic_ctrls_2_down_BtbPlugin_logic_chunksLogic_1_readRsp_ENTRY_sliceLow,fetch_logic_ctrls_2_down_BtbPlugin_logic_chunksLogic_1_readRsp_ENTRY_hash};
  assign _zz_AlignerPlugin_logic_buffer_flushIt = 1'b1;
  assign _zz_AlignerPlugin_logic_buffer_flushIt_1 = (early0_EnvPlugin_logic_flushPort_valid && 1'b1);
  assign _zz_AlignerPlugin_logic_buffer_flushIt_2 = (CsrAccessPlugin_logic_flushPort_valid && 1'b1);
  assign _zz_AlignerPlugin_logic_buffer_flushIt_3 = {(early0_BranchPlugin_logic_flushPort_valid && 1'b1),(LsuPlugin_logic_flushPort_valid && 1'b1)};
  assign _zz_AlignerPlugin_logic_extractors_0_ctx_instruction_1 = _zz_AlignerPlugin_logic_extractors_0_ctx_instruction[0];
  assign _zz_AlignerPlugin_logic_extractors_0_ctx_instruction_2 = 32'h0;
  assign _zz_AlignerPlugin_logic_extractors_0_ctx_instruction_3 = _zz_AlignerPlugin_logic_extractors_0_ctx_instruction[1];
  assign _zz_AlignerPlugin_logic_extractors_0_ctx_instruction_4 = 32'h0;
  assign _zz_AlignerPlugin_logic_extractors_0_ctx_instruction_5 = _zz_AlignerPlugin_logic_extractors_0_ctx_instruction[2];
  assign _zz_AlignerPlugin_logic_extractors_0_ctx_instruction_6 = 32'h0;
  assign _zz_AlignerPlugin_logic_extractors_0_ctx_instruction_7 = _zz_AlignerPlugin_logic_extractors_0_ctx_instruction[3];
  assign _zz_AlignerPlugin_logic_extractors_0_ctx_instruction_8 = 32'h0;
  assign _zz_AlignerPlugin_logic_extractors_0_ctx_instruction_9 = _zz_AlignerPlugin_logic_extractors_0_ctx_instruction[4];
  assign _zz_AlignerPlugin_logic_extractors_0_ctx_instruction_10 = 32'h0;
  assign _zz_AlignerPlugin_logic_extractors_0_ctx_instruction_11 = _zz_AlignerPlugin_logic_extractors_0_ctx_instruction[5];
  assign _zz_AlignerPlugin_logic_extractors_0_ctx_instruction_12 = 32'h0;
  assign _zz_AlignerPlugin_logic_extractors_0_ctx_instruction_13 = _zz_AlignerPlugin_logic_extractors_0_ctx_instruction[6];
  assign _zz_AlignerPlugin_logic_extractors_0_ctx_instruction_14 = 32'h0;
  assign _zz_AlignerPlugin_logic_extractors_0_ctx_instruction_15 = _zz_AlignerPlugin_logic_extractors_0_ctx_instruction[7];
  assign _zz_AlignerPlugin_logic_extractors_0_ctx_instruction_16 = 32'h0;
  assign _zz_DispatchPlugin_logic_candidates_0_cancel = 1'b1;
  assign _zz_DispatchPlugin_logic_candidates_0_cancel_1 = 1'b1;
  assign _zz__zz_DispatchPlugin_logic_slots_0_ctx_valid_4 = DispatchPlugin_logic_candidates_1_ctx_hm_DispatchPlugin_logic_hcs_3_onRs_0_ENABLES_0;
  assign _zz__zz_DispatchPlugin_logic_slots_0_ctx_valid_4_1 = {DispatchPlugin_logic_candidates_1_ctx_hm_DispatchPlugin_logic_hcs_2_onRs_1_ENABLES_0,{DispatchPlugin_logic_candidates_1_ctx_hm_DispatchPlugin_logic_hcs_2_onRs_0_ENABLES_0,{DispatchPlugin_logic_candidates_1_ctx_hm_DispatchPlugin_logic_hcs_1_onRs_1_ENABLES_1,{DispatchPlugin_logic_candidates_1_ctx_hm_DispatchPlugin_logic_hcs_1_onRs_1_ENABLES_0,{DispatchPlugin_logic_candidates_1_ctx_hm_DispatchPlugin_logic_hcs_1_onRs_0_ENABLES_0,{_zz__zz_DispatchPlugin_logic_slots_0_ctx_valid_4_2,_zz__zz_DispatchPlugin_logic_slots_0_ctx_valid_4_3}}}}}};
  assign _zz__zz_DispatchPlugin_logic_slots_0_ctx_valid_4_10 = DispatchPlugin_logic_candidates_1_ctx_valid;
  assign _zz__zz_DispatchPlugin_logic_slots_0_ctx_valid_4_11 = DispatchPlugin_logic_candidates_2_ctx_hm_DispatchPlugin_logic_hcs_3_onRs_0_ENABLES_0;
  assign _zz__zz_DispatchPlugin_logic_slots_0_ctx_valid_4_12 = {DispatchPlugin_logic_candidates_2_ctx_hm_DispatchPlugin_logic_hcs_2_onRs_1_ENABLES_0,{DispatchPlugin_logic_candidates_2_ctx_hm_DispatchPlugin_logic_hcs_2_onRs_0_ENABLES_0,{DispatchPlugin_logic_candidates_2_ctx_hm_DispatchPlugin_logic_hcs_1_onRs_1_ENABLES_1,{DispatchPlugin_logic_candidates_2_ctx_hm_DispatchPlugin_logic_hcs_1_onRs_1_ENABLES_0,{DispatchPlugin_logic_candidates_2_ctx_hm_DispatchPlugin_logic_hcs_1_onRs_0_ENABLES_0,{_zz__zz_DispatchPlugin_logic_slots_0_ctx_valid_4_13,_zz__zz_DispatchPlugin_logic_slots_0_ctx_valid_4_14}}}}}};
  assign _zz__zz_DispatchPlugin_logic_slots_0_ctx_valid_4_21 = DispatchPlugin_logic_candidates_2_ctx_valid;
  assign _zz__zz_DispatchPlugin_logic_slots_0_ctx_valid_4_2 = DispatchPlugin_logic_candidates_1_ctx_hm_DispatchPlugin_logic_hcs_0_onRs_1_ENABLES_0;
  assign _zz__zz_DispatchPlugin_logic_slots_0_ctx_valid_4_3 = {DispatchPlugin_logic_candidates_1_ctx_hm_DispatchPlugin_logic_hcs_0_onRs_0_ENABLES_0,{DispatchPlugin_logic_candidates_1_ctx_hm_RD_PHYS,{DispatchPlugin_logic_candidates_1_ctx_hm_RD_ENABLE,{DispatchPlugin_logic_candidates_1_ctx_hm_RS2_PHYS,{DispatchPlugin_logic_candidates_1_ctx_hm_RS2_ENABLE,{DispatchPlugin_logic_candidates_1_ctx_hm_RS1_PHYS,{_zz__zz_DispatchPlugin_logic_slots_0_ctx_valid_4_4,_zz__zz_DispatchPlugin_logic_slots_0_ctx_valid_4_5}}}}}}};
  assign _zz__zz_DispatchPlugin_logic_slots_0_ctx_valid_4_13 = DispatchPlugin_logic_candidates_2_ctx_hm_DispatchPlugin_logic_hcs_0_onRs_1_ENABLES_0;
  assign _zz__zz_DispatchPlugin_logic_slots_0_ctx_valid_4_14 = {DispatchPlugin_logic_candidates_2_ctx_hm_DispatchPlugin_logic_hcs_0_onRs_0_ENABLES_0,{DispatchPlugin_logic_candidates_2_ctx_hm_RD_PHYS,{DispatchPlugin_logic_candidates_2_ctx_hm_RD_ENABLE,{DispatchPlugin_logic_candidates_2_ctx_hm_RS2_PHYS,{DispatchPlugin_logic_candidates_2_ctx_hm_RS2_ENABLE,{DispatchPlugin_logic_candidates_2_ctx_hm_RS1_PHYS,{_zz__zz_DispatchPlugin_logic_slots_0_ctx_valid_4_15,_zz__zz_DispatchPlugin_logic_slots_0_ctx_valid_4_16}}}}}}};
  assign _zz__zz_DispatchPlugin_logic_slots_0_ctx_valid_4_4 = DispatchPlugin_logic_candidates_1_ctx_hm_RS1_ENABLE;
  assign _zz__zz_DispatchPlugin_logic_slots_0_ctx_valid_4_5 = {DispatchPlugin_logic_candidates_1_ctx_hm_Decode_UOP_ID,{DispatchPlugin_logic_candidates_1_ctx_hm_TRAP,{DispatchPlugin_logic_candidates_1_ctx_hm_PC,{DispatchPlugin_logic_candidates_1_ctx_hm_DONT_FLUSH_PRECISE_4,{DispatchPlugin_logic_candidates_1_ctx_hm_DONT_FLUSH_PRECISE_3,{_zz__zz_DispatchPlugin_logic_slots_0_ctx_valid_4_6,_zz__zz_DispatchPlugin_logic_slots_0_ctx_valid_4_7}}}}}};
  assign _zz__zz_DispatchPlugin_logic_slots_0_ctx_valid_4_15 = DispatchPlugin_logic_candidates_2_ctx_hm_RS1_ENABLE;
  assign _zz__zz_DispatchPlugin_logic_slots_0_ctx_valid_4_16 = {DispatchPlugin_logic_candidates_2_ctx_hm_Decode_UOP_ID,{DispatchPlugin_logic_candidates_2_ctx_hm_TRAP,{DispatchPlugin_logic_candidates_2_ctx_hm_PC,{DispatchPlugin_logic_candidates_2_ctx_hm_DONT_FLUSH_PRECISE_4,{DispatchPlugin_logic_candidates_2_ctx_hm_DONT_FLUSH_PRECISE_3,{_zz__zz_DispatchPlugin_logic_slots_0_ctx_valid_4_17,_zz__zz_DispatchPlugin_logic_slots_0_ctx_valid_4_18}}}}}};
  assign _zz__zz_DispatchPlugin_logic_slots_0_ctx_valid_4_6 = DispatchPlugin_logic_candidates_1_ctx_hm_Decode_INSTRUCTION_SLICE_COUNT;
  assign _zz__zz_DispatchPlugin_logic_slots_0_ctx_valid_4_7 = {DispatchPlugin_logic_candidates_1_ctx_hm_DispatchPlugin_DONT_FLUSH_FROM_LANES,{DispatchPlugin_logic_candidates_1_ctx_hm_DispatchPlugin_DONT_FLUSH,{DispatchPlugin_logic_candidates_1_ctx_hm_DispatchPlugin_MAY_FLUSH,{DispatchPlugin_logic_candidates_1_ctx_hm_DispatchPlugin_FENCE_OLDER,{DispatchPlugin_logic_candidates_1_ctx_hm_Prediction_BRANCH_HISTORY,{_zz__zz_DispatchPlugin_logic_slots_0_ctx_valid_4_8,_zz__zz_DispatchPlugin_logic_slots_0_ctx_valid_4_9}}}}}};
  assign _zz__zz_DispatchPlugin_logic_slots_0_ctx_valid_4_17 = DispatchPlugin_logic_candidates_2_ctx_hm_Decode_INSTRUCTION_SLICE_COUNT;
  assign _zz__zz_DispatchPlugin_logic_slots_0_ctx_valid_4_18 = {DispatchPlugin_logic_candidates_2_ctx_hm_DispatchPlugin_DONT_FLUSH_FROM_LANES,{DispatchPlugin_logic_candidates_2_ctx_hm_DispatchPlugin_DONT_FLUSH,{DispatchPlugin_logic_candidates_2_ctx_hm_DispatchPlugin_MAY_FLUSH,{DispatchPlugin_logic_candidates_2_ctx_hm_DispatchPlugin_FENCE_OLDER,{DispatchPlugin_logic_candidates_2_ctx_hm_Prediction_BRANCH_HISTORY,{_zz__zz_DispatchPlugin_logic_slots_0_ctx_valid_4_19,_zz__zz_DispatchPlugin_logic_slots_0_ctx_valid_4_20}}}}}};
  assign _zz__zz_DispatchPlugin_logic_slots_0_ctx_valid_4_8 = {DispatchPlugin_logic_candidates_1_ctx_hm_GSharePlugin_GSHARE_COUNTER_3,{DispatchPlugin_logic_candidates_1_ctx_hm_GSharePlugin_GSHARE_COUNTER_2,{DispatchPlugin_logic_candidates_1_ctx_hm_GSharePlugin_GSHARE_COUNTER_1,DispatchPlugin_logic_candidates_1_ctx_hm_GSharePlugin_GSHARE_COUNTER_0}}};
  assign _zz__zz_DispatchPlugin_logic_slots_0_ctx_valid_4_9 = {DispatchPlugin_logic_candidates_1_ctx_hm_Prediction_ALIGNED_SLICES_BRANCH,{DispatchPlugin_logic_candidates_1_ctx_hm_Prediction_ALIGNED_SLICES_TAKEN,{DispatchPlugin_logic_candidates_1_ctx_hm_Prediction_ALIGNED_JUMPED_PC,DispatchPlugin_logic_candidates_1_ctx_hm_Prediction_ALIGNED_JUMPED}}};
  assign _zz__zz_DispatchPlugin_logic_slots_0_ctx_valid_4_19 = {DispatchPlugin_logic_candidates_2_ctx_hm_GSharePlugin_GSHARE_COUNTER_3,{DispatchPlugin_logic_candidates_2_ctx_hm_GSharePlugin_GSHARE_COUNTER_2,{DispatchPlugin_logic_candidates_2_ctx_hm_GSharePlugin_GSHARE_COUNTER_1,DispatchPlugin_logic_candidates_2_ctx_hm_GSharePlugin_GSHARE_COUNTER_0}}};
  assign _zz__zz_DispatchPlugin_logic_slots_0_ctx_valid_4_20 = {DispatchPlugin_logic_candidates_2_ctx_hm_Prediction_ALIGNED_SLICES_BRANCH,{DispatchPlugin_logic_candidates_2_ctx_hm_Prediction_ALIGNED_SLICES_TAKEN,{DispatchPlugin_logic_candidates_2_ctx_hm_Prediction_ALIGNED_JUMPED_PC,DispatchPlugin_logic_candidates_2_ctx_hm_Prediction_ALIGNED_JUMPED}}};
  assign _zz__zz_toplevel_execute_ctrl0_up_GSharePlugin_GSHARE_COUNTER_lane0_0 = DispatchPlugin_logic_candidates_0_ctx_hm_GSharePlugin_GSHARE_COUNTER_2;
  assign _zz__zz_toplevel_execute_ctrl0_up_GSharePlugin_GSHARE_COUNTER_lane0_0_1 = {DispatchPlugin_logic_candidates_0_ctx_hm_GSharePlugin_GSHARE_COUNTER_1,DispatchPlugin_logic_candidates_0_ctx_hm_GSharePlugin_GSHARE_COUNTER_0};
  assign _zz__zz_toplevel_execute_ctrl0_up_GSharePlugin_GSHARE_COUNTER_lane0_0_2 = DispatchPlugin_logic_candidates_1_ctx_hm_GSharePlugin_GSHARE_COUNTER_2;
  assign _zz__zz_toplevel_execute_ctrl0_up_GSharePlugin_GSHARE_COUNTER_lane0_0_3 = {DispatchPlugin_logic_candidates_1_ctx_hm_GSharePlugin_GSHARE_COUNTER_1,DispatchPlugin_logic_candidates_1_ctx_hm_GSharePlugin_GSHARE_COUNTER_0};
  assign _zz__zz_toplevel_execute_ctrl0_up_GSharePlugin_GSHARE_COUNTER_lane0_0_4 = DispatchPlugin_logic_candidates_2_ctx_hm_GSharePlugin_GSHARE_COUNTER_1;
  assign _zz__zz_toplevel_execute_ctrl0_up_GSharePlugin_GSHARE_COUNTER_lane0_0_5 = DispatchPlugin_logic_candidates_2_ctx_hm_GSharePlugin_GSHARE_COUNTER_0;
  assign _zz__zz_toplevel_execute_ctrl0_up_GSharePlugin_GSHARE_COUNTER_lane1_0 = DispatchPlugin_logic_candidates_0_ctx_hm_GSharePlugin_GSHARE_COUNTER_1;
  assign _zz__zz_toplevel_execute_ctrl0_up_GSharePlugin_GSHARE_COUNTER_lane1_0_1 = DispatchPlugin_logic_candidates_0_ctx_hm_GSharePlugin_GSHARE_COUNTER_0;
  assign _zz__zz_toplevel_execute_ctrl0_up_GSharePlugin_GSHARE_COUNTER_lane1_0_2 = DispatchPlugin_logic_candidates_1_ctx_hm_GSharePlugin_GSHARE_COUNTER_1;
  assign _zz__zz_toplevel_execute_ctrl0_up_GSharePlugin_GSHARE_COUNTER_lane1_0_3 = DispatchPlugin_logic_candidates_1_ctx_hm_GSharePlugin_GSHARE_COUNTER_0;
  assign _zz_decode_logic_flushes_0_onLanes_0_doIt = 1'b1;
  assign _zz_decode_logic_flushes_0_onLanes_0_doIt_1 = (CsrAccessPlugin_logic_flushPort_valid && 1'b1);
  assign _zz_decode_logic_flushes_0_onLanes_0_doIt_2 = (early0_BranchPlugin_logic_flushPort_valid && 1'b1);
  assign _zz_decode_logic_flushes_0_onLanes_0_doIt_3 = (LsuPlugin_logic_flushPort_valid && 1'b1);
  assign _zz_decode_logic_flushes_0_onLanes_1_doIt = 1'b1;
  assign _zz_decode_logic_flushes_0_onLanes_1_doIt_1 = (CsrAccessPlugin_logic_flushPort_valid && 1'b1);
  assign _zz_decode_logic_flushes_0_onLanes_1_doIt_2 = (early0_BranchPlugin_logic_flushPort_valid && 1'b1);
  assign _zz_decode_logic_flushes_0_onLanes_1_doIt_3 = (LsuPlugin_logic_flushPort_valid && 1'b1);
  assign _zz_decode_logic_flushes_1_onLanes_0_doIt = 1'b0;
  assign _zz_decode_logic_flushes_1_onLanes_0_doIt_1 = (DecoderPlugin_logic_laneLogic_1_flushPort_payload_laneAge == 1'b0);
  assign _zz_decode_logic_flushes_1_onLanes_0_doIt_2 = 1'b1;
  assign _zz_decode_logic_flushes_1_onLanes_0_doIt_3 = (DecoderPlugin_logic_laneLogic_0_flushPort_payload_laneAge < 1'b0);
  assign _zz_decode_logic_flushes_1_onLanes_0_doIt_4 = ((DecoderPlugin_logic_laneLogic_0_flushPort_payload_laneAge == 1'b0) && DecoderPlugin_logic_laneLogic_0_flushPort_payload_self);
  assign _zz_decode_logic_flushes_1_onLanes_0_doIt_5 = 1'b1;
  assign _zz_decode_logic_flushes_1_onLanes_0_doIt_6 = (early1_BranchPlugin_logic_flushPort_valid && 1'b1);
  assign _zz_decode_logic_flushes_1_onLanes_0_doIt_7 = (late0_BranchPlugin_logic_flushPort_valid && 1'b1);
  assign _zz_decode_logic_flushes_1_onLanes_0_doIt_8 = {(early0_EnvPlugin_logic_flushPort_valid && 1'b1),{(CsrAccessPlugin_logic_flushPort_valid && 1'b1),{(early0_BranchPlugin_logic_flushPort_valid && 1'b1),(LsuPlugin_logic_flushPort_valid && 1'b1)}}};
  assign _zz_decode_logic_flushes_1_onLanes_1_doIt_1 = (DecoderPlugin_logic_laneLogic_0_flushPort_payload_laneAge == _zz_decode_logic_flushes_1_onLanes_1_doIt);
  assign _zz_decode_logic_flushes_1_onLanes_1_doIt_2 = 1'b1;
  assign _zz_decode_logic_flushes_1_onLanes_1_doIt_3 = (late0_BranchPlugin_logic_flushPort_valid && 1'b1);
  assign _zz_decode_logic_flushes_1_onLanes_1_doIt_4 = (early0_EnvPlugin_logic_flushPort_valid && 1'b1);
  assign _zz_decode_logic_flushes_1_onLanes_1_doIt_5 = {(CsrAccessPlugin_logic_flushPort_valid && 1'b1),{(early0_BranchPlugin_logic_flushPort_valid && 1'b1),(LsuPlugin_logic_flushPort_valid && 1'b1)}};
  assign _zz__zz_TrapPlugin_logic_harts_0_trap_pending_arbiter_down_payload_exception = {TrapPlugin_logic_harts_0_trap_pending_arbiter_ports_0_payload_tval,TrapPlugin_logic_harts_0_trap_pending_arbiter_ports_0_payload_exception};
  assign _zz__zz_TrapPlugin_logic_harts_0_trap_pending_arbiter_down_payload_exception_1 = {TrapPlugin_logic_harts_0_trap_pending_arbiter_ports_1_payload_tval,TrapPlugin_logic_harts_0_trap_pending_arbiter_ports_1_payload_exception};
  assign _zz__zz_TrapPlugin_logic_harts_0_trap_pending_arbiter_down_payload_exception_2 = {TrapPlugin_logic_harts_0_trap_pending_arbiter_ports_2_payload_tval,TrapPlugin_logic_harts_0_trap_pending_arbiter_ports_2_payload_exception};
  assign _zz__zz_TrapPlugin_logic_harts_0_trap_pending_arbiter_down_payload_exception_3 = {TrapPlugin_logic_harts_0_trap_pending_arbiter_ports_3_payload_tval,TrapPlugin_logic_harts_0_trap_pending_arbiter_ports_3_payload_exception};
  assign _zz_LsuPlugin_logic_onAddress0_translationPort_logic_ctrl_lineTranslated = toplevel_execute_ctrl3_down_LsuL1_MIXED_ADDRESS_lane0[11 : 0];
  assign _zz_LsuPlugin_logic_onAddress0_translationPort_logic_ctrl_lineTranslated_1 = toplevel_execute_ctrl3_down_LsuL1_MIXED_ADDRESS_lane0[11 : 0];
  assign _zz_FetchL1Plugin_logic_translationPort_logic_ctrl_lineTranslated = fetch_logic_ctrls_1_down_Fetch_WORD_PC[11 : 0];
  assign _zz_FetchL1Plugin_logic_translationPort_logic_ctrl_lineTranslated_1 = fetch_logic_ctrls_1_down_Fetch_WORD_PC[11 : 0];
  assign _zz_PcPlugin_logic_harts_0_aggregator_target_7 = TrapPlugin_logic_harts_0_trap_pcPort_payload_pc;
  assign _zz_PcPlugin_logic_harts_0_aggregator_target_8 = 32'h0;
  assign _zz_PcPlugin_logic_harts_0_aggregator_target_9 = late0_BranchPlugin_logic_pcPort_payload_pc;
  assign _zz_PcPlugin_logic_harts_0_aggregator_target_10 = 32'h0;
  assign _zz_PcPlugin_logic_harts_0_aggregator_target_11 = late1_BranchPlugin_logic_pcPort_payload_pc;
  assign _zz_PcPlugin_logic_harts_0_aggregator_target_12 = 32'h0;
  assign _zz_PcPlugin_logic_harts_0_aggregator_target_13 = early0_BranchPlugin_logic_pcPort_payload_pc;
  assign _zz_PcPlugin_logic_harts_0_aggregator_target_14 = 32'h0;
  assign _zz_PcPlugin_logic_harts_0_aggregator_target_15 = early1_BranchPlugin_logic_pcPort_payload_pc;
  assign _zz_PcPlugin_logic_harts_0_aggregator_target_16 = 32'h0;
  assign _zz_PcPlugin_logic_harts_0_aggregator_target_17 = BtbPlugin_logic_pcPort_payload_pc;
  assign _zz_PcPlugin_logic_harts_0_aggregator_target_18 = 32'h0;
  assign _zz_COMB_CSR_CsrRamPlugin_csrMapper_selFilter = 12'h340;
  assign _zz_COMB_CSR_CsrRamPlugin_csrMapper_selFilter_1 = (CsrAccessPlugin_logic_fsm_inject_csrAddress == 12'h341);
  assign _zz_COMB_CSR_CsrRamPlugin_csrMapper_selFilter_2 = (CsrAccessPlugin_logic_fsm_inject_csrAddress == 12'h343);
  assign _zz_COMB_CSR_CsrRamPlugin_csrMapper_selFilter_3 = (CsrAccessPlugin_logic_fsm_inject_csrAddress == 12'h305);
  assign _zz_CsrAccessPlugin_logic_fsm_inject_implemented = COMB_CSR_322;
  assign _zz_CsrAccessPlugin_logic_fsm_inject_implemented_1 = {COMB_CSR_771,{COMB_CSR_770,{COMB_CSR_772,{COMB_CSR_836,{COMB_CSR_834,{COMB_CSR_768,{COMB_CSR_769,{COMB_CSR_3860,{COMB_CSR_3859,{COMB_CSR_3858,{_zz_CsrAccessPlugin_logic_fsm_inject_implemented_2,_zz_CsrAccessPlugin_logic_fsm_inject_implemented_3}}}}}}}}}}};
  assign _zz_CsrAccessPlugin_logic_fsm_inject_implemented_2 = COMB_CSR_3857;
  assign _zz_CsrAccessPlugin_logic_fsm_inject_implemented_3 = {COMB_CSR_1954,{COMB_CSR_1953,COMB_CSR_1952}};
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_13 = (32'h0 | _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_14);
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_16 = (32'h0 | 32'h0);
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_17 = (((when_CsrService_l188 && REG_CSR_769) ? 32'h40141105 : 32'h0) | _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_18);
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_20 = (_zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_21 | _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_23);
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_25 = (_zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_26 | _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_27);
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_29 = (_zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_30 | _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_32);
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_34 = (_zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_35 | _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_37);
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_38 = (_zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_39 | _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_41);
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_43 = (_zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_44 | _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_46);
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_48 = (_zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_49 | _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_51);
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_53 = (_zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_54 | _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_56);
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_58 = (_zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_59 | _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_61);
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_63 = (_zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_64 | _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_66);
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_68 = (_zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_69 | _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_71);
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_73 = (_zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_74 | _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_76);
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_78 = (_zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_79 | _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_81);
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_82 = (_zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_83 | _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_85);
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_86 = (_zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_87 | _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_89);
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_91 = (_zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_92 | _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_94);
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_96 = (_zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_97 | _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_99);
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_101 = (_zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_102 | _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_104);
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_106 = (_zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_107 | _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_109);
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_111 = (_zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_112 | _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_114);
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_116 = (_zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_117 | _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_119);
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_121 = (_zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_122 | _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_124);
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_126 = (_zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_127 | _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_129);
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_131 = (_zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_132 | ((when_CsrService_l188 && REG_CSR_3073) ? PrivilegedPlugin_logic_rdtime[31 : 0] : 32'h0));
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_134 = (((when_CsrService_l188 && REG_CSR_3201) ? PrivilegedPlugin_logic_rdtime[63 : 32] : 32'h0) | _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_135);
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_137 = (_zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_138 | _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_140);
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_142 = (_zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_143 | _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_145);
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_147 = (_zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_148 | _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_149);
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_151 = (CsrRamPlugin_csrMapper_withRead ? CsrRamPlugin_csrMapper_read_data : 32'h0);
  assign _zz__zz_toplevel_execute_ctrl1_down_integer_RS1_lane0_1 = _zz_toplevel_execute_ctrl1_down_integer_RS1_lane0[0];
  assign _zz__zz_toplevel_execute_ctrl1_down_integer_RS1_lane0_1_1 = 32'h0;
  assign _zz__zz_toplevel_execute_ctrl1_down_integer_RS1_lane0_1_2 = _zz_toplevel_execute_ctrl1_down_integer_RS1_lane0[1];
  assign _zz__zz_toplevel_execute_ctrl1_down_integer_RS1_lane0_1_3 = 32'h0;
  assign _zz__zz_toplevel_execute_ctrl1_down_integer_RS1_lane0_1_4 = _zz_toplevel_execute_ctrl1_down_integer_RS1_lane0[2];
  assign _zz__zz_toplevel_execute_ctrl1_down_integer_RS1_lane0_1_5 = 32'h0;
  assign _zz__zz_toplevel_execute_ctrl1_down_integer_RS1_lane0_1_6 = _zz_toplevel_execute_ctrl1_down_integer_RS1_lane0[3];
  assign _zz__zz_toplevel_execute_ctrl1_down_integer_RS1_lane0_1_7 = 32'h0;
  assign _zz__zz_toplevel_execute_ctrl1_down_integer_RS1_lane0_1_8 = _zz_toplevel_execute_ctrl1_down_integer_RS1_lane0[4];
  assign _zz__zz_toplevel_execute_ctrl1_down_integer_RS1_lane0_1_9 = 32'h0;
  assign _zz__zz_toplevel_execute_ctrl1_down_integer_RS1_lane0_1_10 = _zz_toplevel_execute_ctrl1_down_integer_RS1_lane0[5];
  assign _zz__zz_toplevel_execute_ctrl1_down_integer_RS1_lane0_1_11 = 32'h0;
  assign _zz__zz_toplevel_execute_ctrl1_down_integer_RS1_lane0_1_12 = _zz_toplevel_execute_ctrl1_down_integer_RS1_lane0[6];
  assign _zz__zz_toplevel_execute_ctrl1_down_integer_RS1_lane0_1_13 = 32'h0;
  assign _zz__zz_toplevel_execute_ctrl1_down_integer_RS1_lane0_1_14 = _zz_toplevel_execute_ctrl1_down_integer_RS1_lane0[7];
  assign _zz__zz_toplevel_execute_ctrl1_down_integer_RS1_lane0_1_15 = 32'h0;
  assign _zz__zz_toplevel_execute_ctrl1_down_integer_RS2_lane0_1 = _zz_toplevel_execute_ctrl1_down_integer_RS2_lane0[0];
  assign _zz__zz_toplevel_execute_ctrl1_down_integer_RS2_lane0_1_1 = 32'h0;
  assign _zz__zz_toplevel_execute_ctrl1_down_integer_RS2_lane0_1_2 = _zz_toplevel_execute_ctrl1_down_integer_RS2_lane0[1];
  assign _zz__zz_toplevel_execute_ctrl1_down_integer_RS2_lane0_1_3 = 32'h0;
  assign _zz__zz_toplevel_execute_ctrl1_down_integer_RS2_lane0_1_4 = _zz_toplevel_execute_ctrl1_down_integer_RS2_lane0[2];
  assign _zz__zz_toplevel_execute_ctrl1_down_integer_RS2_lane0_1_5 = 32'h0;
  assign _zz__zz_toplevel_execute_ctrl1_down_integer_RS2_lane0_1_6 = _zz_toplevel_execute_ctrl1_down_integer_RS2_lane0[3];
  assign _zz__zz_toplevel_execute_ctrl1_down_integer_RS2_lane0_1_7 = 32'h0;
  assign _zz__zz_toplevel_execute_ctrl1_down_integer_RS2_lane0_1_8 = _zz_toplevel_execute_ctrl1_down_integer_RS2_lane0[4];
  assign _zz__zz_toplevel_execute_ctrl1_down_integer_RS2_lane0_1_9 = 32'h0;
  assign _zz__zz_toplevel_execute_ctrl1_down_integer_RS2_lane0_1_10 = _zz_toplevel_execute_ctrl1_down_integer_RS2_lane0[5];
  assign _zz__zz_toplevel_execute_ctrl1_down_integer_RS2_lane0_1_11 = 32'h0;
  assign _zz__zz_toplevel_execute_ctrl1_down_integer_RS2_lane0_1_12 = _zz_toplevel_execute_ctrl1_down_integer_RS2_lane0[6];
  assign _zz__zz_toplevel_execute_ctrl1_down_integer_RS2_lane0_1_13 = 32'h0;
  assign _zz__zz_toplevel_execute_ctrl1_down_integer_RS2_lane0_1_14 = _zz_toplevel_execute_ctrl1_down_integer_RS2_lane0[7];
  assign _zz__zz_toplevel_execute_ctrl1_down_integer_RS2_lane0_1_15 = 32'h0;
  assign _zz_toplevel_execute_ctrl1_down_lane0_integer_WriteBackPlugin_SEL_lane0_3 = (execute_lane0_logic_decoding_decodingBits & 33'h000000050);
  assign _zz_toplevel_execute_ctrl1_down_lane0_integer_WriteBackPlugin_SEL_lane0_4 = 33'h000000010;
  assign _zz_toplevel_execute_ctrl1_down_lane0_IntFormatPlugin_logic_WIDTH_ID_lane0 = 33'h000002020;
  assign _zz_toplevel_execute_ctrl1_down_lane0_IntFormatPlugin_logic_WIDTH_ID_lane0_1 = (execute_lane0_logic_decoding_decodingBits & 33'h008002000);
  assign _zz_toplevel_execute_ctrl1_down_lane0_IntFormatPlugin_logic_WIDTH_ID_lane0_2 = 33'h000002000;
  assign _zz__zz_toplevel_execute_ctrl1_down_early0_EnvPlugin_OP_lane0_2 = 33'h002001000;
  assign _zz__zz_toplevel_execute_ctrl1_down_early0_EnvPlugin_OP_lane0_2_1 = 33'h010201000;
  assign _zz__zz_toplevel_execute_ctrl1_down_early0_EnvPlugin_OP_lane0_2_2 = (execute_lane0_logic_decoding_decodingBits & 33'h012400000);
  assign _zz__zz_toplevel_execute_ctrl1_down_early0_EnvPlugin_OP_lane0_2_3 = 33'h010000000;
  assign _zz__zz_toplevel_execute_ctrl1_down_early0_EnvPlugin_OP_lane0_2_4 = ((execute_lane0_logic_decoding_decodingBits & 33'h010100000) == 33'h000100000);
  assign _zz__zz_toplevel_execute_ctrl1_down_early0_EnvPlugin_OP_lane0_2_5 = ((execute_lane0_logic_decoding_decodingBits & 33'h012200000) == 33'h010000000);
  assign _zz_when_ExecuteLanePlugin_l300_2 = (early0_EnvPlugin_logic_flushPort_payload_laneAge == toplevel_execute_ctrl2_down_LANE_AGE_lane0);
  assign _zz_when_ExecuteLanePlugin_l300_2_1 = 1'b1;
  assign _zz_when_ExecuteLanePlugin_l300_2_2 = (CsrAccessPlugin_logic_flushPort_payload_laneAge < toplevel_execute_ctrl2_down_LANE_AGE_lane0);
  assign _zz_when_ExecuteLanePlugin_l300_2_3 = ((CsrAccessPlugin_logic_flushPort_payload_laneAge == toplevel_execute_ctrl2_down_LANE_AGE_lane0) && CsrAccessPlugin_logic_flushPort_payload_self);
  assign _zz_when_ExecuteLanePlugin_l300_2_4 = 1'b1;
  assign _zz_when_ExecuteLanePlugin_l300_2_5 = 1'b1;
  assign _zz_when_ExecuteLanePlugin_l300_3 = 1'b1;
  assign _zz_when_ExecuteLanePlugin_l300_3_1 = (early0_BranchPlugin_logic_flushPort_payload_laneAge < toplevel_execute_ctrl3_down_LANE_AGE_lane0);
  assign _zz_when_ExecuteLanePlugin_l300_3_2 = ((early0_BranchPlugin_logic_flushPort_payload_laneAge == toplevel_execute_ctrl3_down_LANE_AGE_lane0) && early0_BranchPlugin_logic_flushPort_payload_self);
  assign _zz_when_ExecuteLanePlugin_l300_4 = (late0_BranchPlugin_logic_flushPort_payload_laneAge == toplevel_execute_ctrl4_down_LANE_AGE_lane0);
  assign _zz_when_ExecuteLanePlugin_l300_4_1 = (LsuPlugin_logic_flushPort_payload_laneAge == toplevel_execute_ctrl4_down_LANE_AGE_lane0);
  assign _zz_fetch_logic_flushes_0_doIt = 1'b1;
  assign _zz_fetch_logic_flushes_0_doIt_1 = (CsrAccessPlugin_logic_flushPort_valid && 1'b1);
  assign _zz_fetch_logic_flushes_0_doIt_2 = (early0_BranchPlugin_logic_flushPort_valid && 1'b1);
  assign _zz_fetch_logic_flushes_0_doIt_3 = {(LsuPlugin_logic_flushPort_valid && 1'b1),(BtbPlugin_logic_flushPort_valid && 1'b1)};
  assign _zz_fetch_logic_flushes_1_doIt = 1'b1;
  assign _zz_fetch_logic_flushes_1_doIt_1 = (CsrAccessPlugin_logic_flushPort_valid && 1'b1);
  assign _zz_fetch_logic_flushes_1_doIt_2 = (early0_BranchPlugin_logic_flushPort_valid && 1'b1);
  assign _zz_fetch_logic_flushes_1_doIt_3 = {(LsuPlugin_logic_flushPort_valid && 1'b1),((BtbPlugin_logic_flushPort_valid && 1'b1) && (1'b0 || (1'b1 && BtbPlugin_logic_flushPort_payload_self)))};
  assign _zz__zz_toplevel_execute_ctrl1_down_integer_RS1_lane1_1 = _zz_toplevel_execute_ctrl1_down_integer_RS1_lane1[0];
  assign _zz__zz_toplevel_execute_ctrl1_down_integer_RS1_lane1_1_1 = 32'h0;
  assign _zz__zz_toplevel_execute_ctrl1_down_integer_RS1_lane1_1_2 = _zz_toplevel_execute_ctrl1_down_integer_RS1_lane1[1];
  assign _zz__zz_toplevel_execute_ctrl1_down_integer_RS1_lane1_1_3 = 32'h0;
  assign _zz__zz_toplevel_execute_ctrl1_down_integer_RS1_lane1_1_4 = _zz_toplevel_execute_ctrl1_down_integer_RS1_lane1[2];
  assign _zz__zz_toplevel_execute_ctrl1_down_integer_RS1_lane1_1_5 = 32'h0;
  assign _zz__zz_toplevel_execute_ctrl1_down_integer_RS1_lane1_1_6 = _zz_toplevel_execute_ctrl1_down_integer_RS1_lane1[3];
  assign _zz__zz_toplevel_execute_ctrl1_down_integer_RS1_lane1_1_7 = 32'h0;
  assign _zz__zz_toplevel_execute_ctrl1_down_integer_RS1_lane1_1_8 = _zz_toplevel_execute_ctrl1_down_integer_RS1_lane1[4];
  assign _zz__zz_toplevel_execute_ctrl1_down_integer_RS1_lane1_1_9 = 32'h0;
  assign _zz__zz_toplevel_execute_ctrl1_down_integer_RS1_lane1_1_10 = _zz_toplevel_execute_ctrl1_down_integer_RS1_lane1[5];
  assign _zz__zz_toplevel_execute_ctrl1_down_integer_RS1_lane1_1_11 = 32'h0;
  assign _zz__zz_toplevel_execute_ctrl1_down_integer_RS1_lane1_1_12 = _zz_toplevel_execute_ctrl1_down_integer_RS1_lane1[6];
  assign _zz__zz_toplevel_execute_ctrl1_down_integer_RS1_lane1_1_13 = 32'h0;
  assign _zz__zz_toplevel_execute_ctrl1_down_integer_RS1_lane1_1_14 = _zz_toplevel_execute_ctrl1_down_integer_RS1_lane1[7];
  assign _zz__zz_toplevel_execute_ctrl1_down_integer_RS1_lane1_1_15 = 32'h0;
  assign _zz__zz_toplevel_execute_ctrl1_down_integer_RS2_lane1_1 = _zz_toplevel_execute_ctrl1_down_integer_RS2_lane1[0];
  assign _zz__zz_toplevel_execute_ctrl1_down_integer_RS2_lane1_1_1 = 32'h0;
  assign _zz__zz_toplevel_execute_ctrl1_down_integer_RS2_lane1_1_2 = _zz_toplevel_execute_ctrl1_down_integer_RS2_lane1[1];
  assign _zz__zz_toplevel_execute_ctrl1_down_integer_RS2_lane1_1_3 = 32'h0;
  assign _zz__zz_toplevel_execute_ctrl1_down_integer_RS2_lane1_1_4 = _zz_toplevel_execute_ctrl1_down_integer_RS2_lane1[2];
  assign _zz__zz_toplevel_execute_ctrl1_down_integer_RS2_lane1_1_5 = 32'h0;
  assign _zz__zz_toplevel_execute_ctrl1_down_integer_RS2_lane1_1_6 = _zz_toplevel_execute_ctrl1_down_integer_RS2_lane1[3];
  assign _zz__zz_toplevel_execute_ctrl1_down_integer_RS2_lane1_1_7 = 32'h0;
  assign _zz__zz_toplevel_execute_ctrl1_down_integer_RS2_lane1_1_8 = _zz_toplevel_execute_ctrl1_down_integer_RS2_lane1[4];
  assign _zz__zz_toplevel_execute_ctrl1_down_integer_RS2_lane1_1_9 = 32'h0;
  assign _zz__zz_toplevel_execute_ctrl1_down_integer_RS2_lane1_1_10 = _zz_toplevel_execute_ctrl1_down_integer_RS2_lane1[5];
  assign _zz__zz_toplevel_execute_ctrl1_down_integer_RS2_lane1_1_11 = 32'h0;
  assign _zz__zz_toplevel_execute_ctrl1_down_integer_RS2_lane1_1_12 = _zz_toplevel_execute_ctrl1_down_integer_RS2_lane1[6];
  assign _zz__zz_toplevel_execute_ctrl1_down_integer_RS2_lane1_1_13 = 32'h0;
  assign _zz__zz_toplevel_execute_ctrl1_down_integer_RS2_lane1_1_14 = _zz_toplevel_execute_ctrl1_down_integer_RS2_lane1[7];
  assign _zz__zz_toplevel_execute_ctrl1_down_integer_RS2_lane1_1_15 = 32'h0;
  assign _zz_when_ExecuteLanePlugin_l300_7 = (early0_EnvPlugin_logic_flushPort_payload_laneAge == toplevel_execute_ctrl2_down_LANE_AGE_lane1);
  assign _zz_when_ExecuteLanePlugin_l300_7_1 = 1'b1;
  assign _zz_when_ExecuteLanePlugin_l300_7_2 = (CsrAccessPlugin_logic_flushPort_payload_laneAge < toplevel_execute_ctrl2_down_LANE_AGE_lane1);
  assign _zz_when_ExecuteLanePlugin_l300_7_3 = ((CsrAccessPlugin_logic_flushPort_payload_laneAge == toplevel_execute_ctrl2_down_LANE_AGE_lane1) && CsrAccessPlugin_logic_flushPort_payload_self);
  assign _zz_when_ExecuteLanePlugin_l300_7_4 = 1'b1;
  assign _zz_when_ExecuteLanePlugin_l300_7_5 = 1'b1;
  assign _zz_when_ExecuteLanePlugin_l300_8 = 1'b1;
  assign _zz_when_ExecuteLanePlugin_l300_8_1 = (early0_BranchPlugin_logic_flushPort_payload_laneAge < toplevel_execute_ctrl3_down_LANE_AGE_lane1);
  assign _zz_when_ExecuteLanePlugin_l300_8_2 = ((early0_BranchPlugin_logic_flushPort_payload_laneAge == toplevel_execute_ctrl3_down_LANE_AGE_lane1) && early0_BranchPlugin_logic_flushPort_payload_self);
  assign _zz_when_ExecuteLanePlugin_l300_9 = (late0_BranchPlugin_logic_flushPort_payload_laneAge == toplevel_execute_ctrl4_down_LANE_AGE_lane1);
  assign _zz_when_ExecuteLanePlugin_l300_9_1 = (LsuPlugin_logic_flushPort_payload_laneAge == toplevel_execute_ctrl4_down_LANE_AGE_lane1);
  assign BtbPlugin_logic_ras_mem_stack_spinal_port0 = BtbPlugin_logic_ras_mem_stack[BtbPlugin_logic_ras_ptr_pop_aheadValue];
  always @(posedge clk_cpu) begin
    if(_zz_5) begin
      BtbPlugin_logic_ras_mem_stack[BtbPlugin_logic_ras_write_payload_address] <= _zz_BtbPlugin_logic_ras_mem_stack_port;
    end
  end

integer verilogIndex;

initial begin
  for (verilogIndex = 0; verilogIndex < 512; verilogIndex = verilogIndex + 1)begin
FetchL1Plugin_logic_banks_0_mem[verilogIndex] = -1;
  end
end
  always @(posedge clk_cpu) begin
    if(_zz_9) begin
      FetchL1Plugin_logic_banks_0_mem[FetchL1Plugin_logic_banks_0_write_payload_address] <= FetchL1Plugin_logic_banks_0_write_payload_data;
    end
  end

  always @(posedge clk_cpu) begin
    if(FetchL1Plugin_logic_banks_0_read_cmd_valid) begin
      FetchL1Plugin_logic_banks_0_mem_spinal_port1 <= FetchL1Plugin_logic_banks_0_mem[FetchL1Plugin_logic_banks_0_read_cmd_payload];
    end
  end


initial begin
  for (verilogIndex = 0; verilogIndex < 512; verilogIndex = verilogIndex + 1)begin
FetchL1Plugin_logic_banks_1_mem[verilogIndex] = -1;
  end
end
  always @(posedge clk_cpu) begin
    if(_zz_8) begin
      FetchL1Plugin_logic_banks_1_mem[FetchL1Plugin_logic_banks_1_write_payload_address] <= FetchL1Plugin_logic_banks_1_write_payload_data;
    end
  end

  always @(posedge clk_cpu) begin
    if(FetchL1Plugin_logic_banks_1_read_cmd_valid) begin
      FetchL1Plugin_logic_banks_1_mem_spinal_port1 <= FetchL1Plugin_logic_banks_1_mem[FetchL1Plugin_logic_banks_1_read_cmd_payload];
    end
  end


initial begin
  for (verilogIndex = 0; verilogIndex < 64; verilogIndex = verilogIndex + 1)begin
FetchL1Plugin_logic_ways_0_mem[verilogIndex] = -1;
  end
end
  always @(posedge clk_cpu) begin
    if(_zz_FetchL1Plugin_logic_ways_0_mem_port_1) begin
      FetchL1Plugin_logic_ways_0_mem[FetchL1Plugin_logic_waysWrite_address] <= _zz_FetchL1Plugin_logic_ways_0_mem_port;
    end
  end

  always @(posedge clk_cpu) begin
    if(FetchL1Plugin_logic_ways_0_read_cmd_valid) begin
      FetchL1Plugin_logic_ways_0_mem_spinal_port1 <= FetchL1Plugin_logic_ways_0_mem[FetchL1Plugin_logic_ways_0_read_cmd_payload];
    end
  end


initial begin
  for (verilogIndex = 0; verilogIndex < 64; verilogIndex = verilogIndex + 1)begin
FetchL1Plugin_logic_ways_1_mem[verilogIndex] = -1;
  end
end
  always @(posedge clk_cpu) begin
    if(_zz_FetchL1Plugin_logic_ways_1_mem_port_1) begin
      FetchL1Plugin_logic_ways_1_mem[FetchL1Plugin_logic_waysWrite_address] <= _zz_FetchL1Plugin_logic_ways_1_mem_port;
    end
  end

  always @(posedge clk_cpu) begin
    if(FetchL1Plugin_logic_ways_1_read_cmd_valid) begin
      FetchL1Plugin_logic_ways_1_mem_spinal_port1 <= FetchL1Plugin_logic_ways_1_mem[FetchL1Plugin_logic_ways_1_read_cmd_payload];
    end
  end

  always @(posedge clk_cpu) begin
    if(_zz_7) begin
      FetchL1Plugin_logic_plru_mem[FetchL1Plugin_logic_plru_write_payload_address] <= FetchL1Plugin_logic_plru_write_payload_data_0;
    end
  end

  always @(posedge clk_cpu) begin
    if(FetchL1Plugin_logic_plru_read_cmd_valid) begin
      FetchL1Plugin_logic_plru_mem_spinal_port1 <= FetchL1Plugin_logic_plru_mem[FetchL1Plugin_logic_plru_read_cmd_payload];
    end
  end

  always @(posedge clk_cpu) begin
    if(_zz_6) begin
      GSharePlugin_logic_mem_counter[GSharePlugin_logic_mem_write_payload_address] <= _zz_GSharePlugin_logic_mem_counter_port;
    end
  end

  always @(posedge clk_cpu) begin
    if(fetch_logic_ctrls_0_down_isReady) begin
      GSharePlugin_logic_mem_counter_spinal_port1 <= GSharePlugin_logic_mem_counter[fetch_logic_ctrls_0_down_GSharePlugin_logic_HASH];
    end
  end

  always @(*) begin
    BtbPlugin_logic_mem_spinal_port1 = {_zz_BtbPlugin_logic_memsymbol_read_1, _zz_BtbPlugin_logic_memsymbol_read};
  end
  always @(posedge clk_cpu) begin
    if(BtbPlugin_logic_onLearn_port_payload_mask[0] && BtbPlugin_logic_onLearn_port_valid) begin
      BtbPlugin_logic_mem_symbol0[BtbPlugin_logic_onLearn_port_payload_address] <= _zz_BtbPlugin_logic_mem_port[50 : 0];
    end
    if(BtbPlugin_logic_onLearn_port_payload_mask[1] && BtbPlugin_logic_onLearn_port_valid) begin
      BtbPlugin_logic_mem_symbol1[BtbPlugin_logic_onLearn_port_payload_address] <= _zz_BtbPlugin_logic_mem_port[101 : 51];
    end
  end

  always @(posedge clk_cpu) begin
    if(BtbPlugin_logic_readPort_cmd_valid) begin
      _zz_BtbPlugin_logic_memsymbol_read <= BtbPlugin_logic_mem_symbol0[BtbPlugin_logic_readPort_cmd_payload];
      _zz_BtbPlugin_logic_memsymbol_read_1 <= BtbPlugin_logic_mem_symbol1[BtbPlugin_logic_readPort_cmd_payload];
    end
  end

  always @(*) begin
    LsuL1Plugin_logic_banks_0_mem_spinal_port1 = {_zz_LsuL1Plugin_logic_banks_0_memsymbol_read_7, _zz_LsuL1Plugin_logic_banks_0_memsymbol_read_6, _zz_LsuL1Plugin_logic_banks_0_memsymbol_read_5, _zz_LsuL1Plugin_logic_banks_0_memsymbol_read_4, _zz_LsuL1Plugin_logic_banks_0_memsymbol_read_3, _zz_LsuL1Plugin_logic_banks_0_memsymbol_read_2, _zz_LsuL1Plugin_logic_banks_0_memsymbol_read_1, _zz_LsuL1Plugin_logic_banks_0_memsymbol_read};
  end
  always @(posedge clk_cpu) begin
    if(LsuL1Plugin_logic_banks_0_write_payload_mask[0] && LsuL1Plugin_logic_banks_0_write_valid) begin
      LsuL1Plugin_logic_banks_0_mem_symbol0[LsuL1Plugin_logic_banks_0_write_payload_address] <= LsuL1Plugin_logic_banks_0_write_payload_data[7 : 0];
    end
    if(LsuL1Plugin_logic_banks_0_write_payload_mask[1] && LsuL1Plugin_logic_banks_0_write_valid) begin
      LsuL1Plugin_logic_banks_0_mem_symbol1[LsuL1Plugin_logic_banks_0_write_payload_address] <= LsuL1Plugin_logic_banks_0_write_payload_data[15 : 8];
    end
    if(LsuL1Plugin_logic_banks_0_write_payload_mask[2] && LsuL1Plugin_logic_banks_0_write_valid) begin
      LsuL1Plugin_logic_banks_0_mem_symbol2[LsuL1Plugin_logic_banks_0_write_payload_address] <= LsuL1Plugin_logic_banks_0_write_payload_data[23 : 16];
    end
    if(LsuL1Plugin_logic_banks_0_write_payload_mask[3] && LsuL1Plugin_logic_banks_0_write_valid) begin
      LsuL1Plugin_logic_banks_0_mem_symbol3[LsuL1Plugin_logic_banks_0_write_payload_address] <= LsuL1Plugin_logic_banks_0_write_payload_data[31 : 24];
    end
    if(LsuL1Plugin_logic_banks_0_write_payload_mask[4] && LsuL1Plugin_logic_banks_0_write_valid) begin
      LsuL1Plugin_logic_banks_0_mem_symbol4[LsuL1Plugin_logic_banks_0_write_payload_address] <= LsuL1Plugin_logic_banks_0_write_payload_data[39 : 32];
    end
    if(LsuL1Plugin_logic_banks_0_write_payload_mask[5] && LsuL1Plugin_logic_banks_0_write_valid) begin
      LsuL1Plugin_logic_banks_0_mem_symbol5[LsuL1Plugin_logic_banks_0_write_payload_address] <= LsuL1Plugin_logic_banks_0_write_payload_data[47 : 40];
    end
    if(LsuL1Plugin_logic_banks_0_write_payload_mask[6] && LsuL1Plugin_logic_banks_0_write_valid) begin
      LsuL1Plugin_logic_banks_0_mem_symbol6[LsuL1Plugin_logic_banks_0_write_payload_address] <= LsuL1Plugin_logic_banks_0_write_payload_data[55 : 48];
    end
    if(LsuL1Plugin_logic_banks_0_write_payload_mask[7] && LsuL1Plugin_logic_banks_0_write_valid) begin
      LsuL1Plugin_logic_banks_0_mem_symbol7[LsuL1Plugin_logic_banks_0_write_payload_address] <= LsuL1Plugin_logic_banks_0_write_payload_data[63 : 56];
    end
  end

  always @(posedge clk_cpu) begin
    if(LsuL1Plugin_logic_banks_0_read_cmd_valid) begin
      _zz_LsuL1Plugin_logic_banks_0_memsymbol_read <= LsuL1Plugin_logic_banks_0_mem_symbol0[LsuL1Plugin_logic_banks_0_read_cmd_payload];
      _zz_LsuL1Plugin_logic_banks_0_memsymbol_read_1 <= LsuL1Plugin_logic_banks_0_mem_symbol1[LsuL1Plugin_logic_banks_0_read_cmd_payload];
      _zz_LsuL1Plugin_logic_banks_0_memsymbol_read_2 <= LsuL1Plugin_logic_banks_0_mem_symbol2[LsuL1Plugin_logic_banks_0_read_cmd_payload];
      _zz_LsuL1Plugin_logic_banks_0_memsymbol_read_3 <= LsuL1Plugin_logic_banks_0_mem_symbol3[LsuL1Plugin_logic_banks_0_read_cmd_payload];
      _zz_LsuL1Plugin_logic_banks_0_memsymbol_read_4 <= LsuL1Plugin_logic_banks_0_mem_symbol4[LsuL1Plugin_logic_banks_0_read_cmd_payload];
      _zz_LsuL1Plugin_logic_banks_0_memsymbol_read_5 <= LsuL1Plugin_logic_banks_0_mem_symbol5[LsuL1Plugin_logic_banks_0_read_cmd_payload];
      _zz_LsuL1Plugin_logic_banks_0_memsymbol_read_6 <= LsuL1Plugin_logic_banks_0_mem_symbol6[LsuL1Plugin_logic_banks_0_read_cmd_payload];
      _zz_LsuL1Plugin_logic_banks_0_memsymbol_read_7 <= LsuL1Plugin_logic_banks_0_mem_symbol7[LsuL1Plugin_logic_banks_0_read_cmd_payload];
    end
  end

  always @(*) begin
    LsuL1Plugin_logic_banks_1_mem_spinal_port1 = {_zz_LsuL1Plugin_logic_banks_1_memsymbol_read_7, _zz_LsuL1Plugin_logic_banks_1_memsymbol_read_6, _zz_LsuL1Plugin_logic_banks_1_memsymbol_read_5, _zz_LsuL1Plugin_logic_banks_1_memsymbol_read_4, _zz_LsuL1Plugin_logic_banks_1_memsymbol_read_3, _zz_LsuL1Plugin_logic_banks_1_memsymbol_read_2, _zz_LsuL1Plugin_logic_banks_1_memsymbol_read_1, _zz_LsuL1Plugin_logic_banks_1_memsymbol_read};
  end
  always @(posedge clk_cpu) begin
    if(LsuL1Plugin_logic_banks_1_write_payload_mask[0] && LsuL1Plugin_logic_banks_1_write_valid) begin
      LsuL1Plugin_logic_banks_1_mem_symbol0[LsuL1Plugin_logic_banks_1_write_payload_address] <= LsuL1Plugin_logic_banks_1_write_payload_data[7 : 0];
    end
    if(LsuL1Plugin_logic_banks_1_write_payload_mask[1] && LsuL1Plugin_logic_banks_1_write_valid) begin
      LsuL1Plugin_logic_banks_1_mem_symbol1[LsuL1Plugin_logic_banks_1_write_payload_address] <= LsuL1Plugin_logic_banks_1_write_payload_data[15 : 8];
    end
    if(LsuL1Plugin_logic_banks_1_write_payload_mask[2] && LsuL1Plugin_logic_banks_1_write_valid) begin
      LsuL1Plugin_logic_banks_1_mem_symbol2[LsuL1Plugin_logic_banks_1_write_payload_address] <= LsuL1Plugin_logic_banks_1_write_payload_data[23 : 16];
    end
    if(LsuL1Plugin_logic_banks_1_write_payload_mask[3] && LsuL1Plugin_logic_banks_1_write_valid) begin
      LsuL1Plugin_logic_banks_1_mem_symbol3[LsuL1Plugin_logic_banks_1_write_payload_address] <= LsuL1Plugin_logic_banks_1_write_payload_data[31 : 24];
    end
    if(LsuL1Plugin_logic_banks_1_write_payload_mask[4] && LsuL1Plugin_logic_banks_1_write_valid) begin
      LsuL1Plugin_logic_banks_1_mem_symbol4[LsuL1Plugin_logic_banks_1_write_payload_address] <= LsuL1Plugin_logic_banks_1_write_payload_data[39 : 32];
    end
    if(LsuL1Plugin_logic_banks_1_write_payload_mask[5] && LsuL1Plugin_logic_banks_1_write_valid) begin
      LsuL1Plugin_logic_banks_1_mem_symbol5[LsuL1Plugin_logic_banks_1_write_payload_address] <= LsuL1Plugin_logic_banks_1_write_payload_data[47 : 40];
    end
    if(LsuL1Plugin_logic_banks_1_write_payload_mask[6] && LsuL1Plugin_logic_banks_1_write_valid) begin
      LsuL1Plugin_logic_banks_1_mem_symbol6[LsuL1Plugin_logic_banks_1_write_payload_address] <= LsuL1Plugin_logic_banks_1_write_payload_data[55 : 48];
    end
    if(LsuL1Plugin_logic_banks_1_write_payload_mask[7] && LsuL1Plugin_logic_banks_1_write_valid) begin
      LsuL1Plugin_logic_banks_1_mem_symbol7[LsuL1Plugin_logic_banks_1_write_payload_address] <= LsuL1Plugin_logic_banks_1_write_payload_data[63 : 56];
    end
  end

  always @(posedge clk_cpu) begin
    if(LsuL1Plugin_logic_banks_1_read_cmd_valid) begin
      _zz_LsuL1Plugin_logic_banks_1_memsymbol_read <= LsuL1Plugin_logic_banks_1_mem_symbol0[LsuL1Plugin_logic_banks_1_read_cmd_payload];
      _zz_LsuL1Plugin_logic_banks_1_memsymbol_read_1 <= LsuL1Plugin_logic_banks_1_mem_symbol1[LsuL1Plugin_logic_banks_1_read_cmd_payload];
      _zz_LsuL1Plugin_logic_banks_1_memsymbol_read_2 <= LsuL1Plugin_logic_banks_1_mem_symbol2[LsuL1Plugin_logic_banks_1_read_cmd_payload];
      _zz_LsuL1Plugin_logic_banks_1_memsymbol_read_3 <= LsuL1Plugin_logic_banks_1_mem_symbol3[LsuL1Plugin_logic_banks_1_read_cmd_payload];
      _zz_LsuL1Plugin_logic_banks_1_memsymbol_read_4 <= LsuL1Plugin_logic_banks_1_mem_symbol4[LsuL1Plugin_logic_banks_1_read_cmd_payload];
      _zz_LsuL1Plugin_logic_banks_1_memsymbol_read_5 <= LsuL1Plugin_logic_banks_1_mem_symbol5[LsuL1Plugin_logic_banks_1_read_cmd_payload];
      _zz_LsuL1Plugin_logic_banks_1_memsymbol_read_6 <= LsuL1Plugin_logic_banks_1_mem_symbol6[LsuL1Plugin_logic_banks_1_read_cmd_payload];
      _zz_LsuL1Plugin_logic_banks_1_memsymbol_read_7 <= LsuL1Plugin_logic_banks_1_mem_symbol7[LsuL1Plugin_logic_banks_1_read_cmd_payload];
    end
  end

  always @(posedge clk_cpu) begin
    if(_zz_LsuL1Plugin_logic_ways_0_mem_port_1) begin
      LsuL1Plugin_logic_ways_0_mem[LsuL1Plugin_logic_waysWrite_address] <= _zz_LsuL1Plugin_logic_ways_0_mem_port;
    end
  end

  always @(posedge clk_cpu) begin
    if(LsuL1Plugin_logic_ways_0_lsuRead_cmd_valid) begin
      LsuL1Plugin_logic_ways_0_mem_spinal_port1 <= LsuL1Plugin_logic_ways_0_mem[LsuL1Plugin_logic_ways_0_lsuRead_cmd_payload];
    end
  end

  always @(posedge clk_cpu) begin
    if(_zz_LsuL1Plugin_logic_ways_1_mem_port_1) begin
      LsuL1Plugin_logic_ways_1_mem[LsuL1Plugin_logic_waysWrite_address] <= _zz_LsuL1Plugin_logic_ways_1_mem_port;
    end
  end

  always @(posedge clk_cpu) begin
    if(LsuL1Plugin_logic_ways_1_lsuRead_cmd_valid) begin
      LsuL1Plugin_logic_ways_1_mem_spinal_port1 <= LsuL1Plugin_logic_ways_1_mem[LsuL1Plugin_logic_ways_1_lsuRead_cmd_payload];
    end
  end

  always @(posedge clk_cpu) begin
    if(_zz_4) begin
      LsuL1Plugin_logic_shared_mem[LsuL1Plugin_logic_shared_write_payload_address] <= _zz_LsuL1Plugin_logic_shared_mem_port;
    end
  end

  always @(posedge clk_cpu) begin
    if(LsuL1Plugin_logic_shared_lsuRead_cmd_valid) begin
      LsuL1Plugin_logic_shared_mem_spinal_port1 <= LsuL1Plugin_logic_shared_mem[LsuL1Plugin_logic_shared_lsuRead_cmd_payload];
    end
  end

  always @(posedge clk_cpu) begin
    if(_zz_3) begin
      LsuL1Plugin_logic_writeback_victimBuffer[_zz_LsuL1Plugin_logic_writeback_victimBuffer_port] <= LsuL1Plugin_logic_writeback_read_readedData;
    end
  end

  always @(posedge clk_cpu) begin
    if(LsuL1Plugin_logic_writeback_write_bufferRead_ready) begin
      LsuL1Plugin_logic_writeback_victimBuffer_spinal_port1 <= LsuL1Plugin_logic_writeback_victimBuffer[_zz_LsuL1Plugin_logic_writeback_write_word];
    end
  end

  always @(posedge clk_cpu) begin
    if(_zz_FetchL1Plugin_logic_translationStorage_logic_sl_0_ways_0_port_1) begin
      FetchL1Plugin_logic_translationStorage_logic_sl_0_ways_0[FetchL1Plugin_logic_translationStorage_logic_sl_0_write_address] <= _zz_FetchL1Plugin_logic_translationStorage_logic_sl_0_ways_0_port;
    end
  end

  assign FetchL1Plugin_logic_translationStorage_logic_sl_0_ways_0_spinal_port1 = FetchL1Plugin_logic_translationStorage_logic_sl_0_ways_0[FetchL1Plugin_logic_translationPort_logic_read_0_readAddress];
  always @(posedge clk_cpu) begin
    if(_zz_FetchL1Plugin_logic_translationStorage_logic_sl_0_ways_1_port_1) begin
      FetchL1Plugin_logic_translationStorage_logic_sl_0_ways_1[FetchL1Plugin_logic_translationStorage_logic_sl_0_write_address] <= _zz_FetchL1Plugin_logic_translationStorage_logic_sl_0_ways_1_port;
    end
  end

  assign FetchL1Plugin_logic_translationStorage_logic_sl_0_ways_1_spinal_port1 = FetchL1Plugin_logic_translationStorage_logic_sl_0_ways_1[FetchL1Plugin_logic_translationPort_logic_read_0_readAddress];
  always @(posedge clk_cpu) begin
    if(_zz_FetchL1Plugin_logic_translationStorage_logic_sl_1_ways_0_port_1) begin
      FetchL1Plugin_logic_translationStorage_logic_sl_1_ways_0[FetchL1Plugin_logic_translationStorage_logic_sl_1_write_address] <= _zz_FetchL1Plugin_logic_translationStorage_logic_sl_1_ways_0_port;
    end
  end

  assign FetchL1Plugin_logic_translationStorage_logic_sl_1_ways_0_spinal_port1 = FetchL1Plugin_logic_translationStorage_logic_sl_1_ways_0[FetchL1Plugin_logic_translationPort_logic_read_1_readAddress];
  always @(posedge clk_cpu) begin
    if(_zz_LsuPlugin_logic_translationStorage_logic_sl_0_ways_0_port_1) begin
      LsuPlugin_logic_translationStorage_logic_sl_0_ways_0[LsuPlugin_logic_translationStorage_logic_sl_0_write_address] <= _zz_LsuPlugin_logic_translationStorage_logic_sl_0_ways_0_port;
    end
  end

  assign LsuPlugin_logic_translationStorage_logic_sl_0_ways_0_spinal_port1 = LsuPlugin_logic_translationStorage_logic_sl_0_ways_0[LsuPlugin_logic_onAddress0_translationPort_logic_read_0_readAddress];
  always @(posedge clk_cpu) begin
    if(_zz_LsuPlugin_logic_translationStorage_logic_sl_0_ways_1_port_1) begin
      LsuPlugin_logic_translationStorage_logic_sl_0_ways_1[LsuPlugin_logic_translationStorage_logic_sl_0_write_address] <= _zz_LsuPlugin_logic_translationStorage_logic_sl_0_ways_1_port;
    end
  end

  assign LsuPlugin_logic_translationStorage_logic_sl_0_ways_1_spinal_port1 = LsuPlugin_logic_translationStorage_logic_sl_0_ways_1[LsuPlugin_logic_onAddress0_translationPort_logic_read_0_readAddress];
  always @(posedge clk_cpu) begin
    if(_zz_LsuPlugin_logic_translationStorage_logic_sl_1_ways_0_port_1) begin
      LsuPlugin_logic_translationStorage_logic_sl_1_ways_0[LsuPlugin_logic_translationStorage_logic_sl_1_write_address] <= _zz_LsuPlugin_logic_translationStorage_logic_sl_1_ways_0_port;
    end
  end

  assign LsuPlugin_logic_translationStorage_logic_sl_1_ways_0_spinal_port1 = LsuPlugin_logic_translationStorage_logic_sl_1_ways_0[LsuPlugin_logic_onAddress0_translationPort_logic_read_1_readAddress];
  always @(posedge clk_cpu) begin
    if(_zz_2) begin
      CsrRamPlugin_logic_mem[CsrRamPlugin_logic_writeLogic_port_payload_address] <= CsrRamPlugin_logic_writeLogic_port_payload_data;
    end
  end

  always @(posedge clk_cpu) begin
    if(CsrRamPlugin_logic_readLogic_port_cmd_valid) begin
      CsrRamPlugin_logic_mem_spinal_port1 <= CsrRamPlugin_logic_mem[CsrRamPlugin_logic_readLogic_port_cmd_payload];
    end
  end

  DivRadix early0_DivPlugin_logic_processing_div (
    .io_flush                  (toplevel_execute_ctrl2_down_isReady                              ), //i
    .io_cmd_valid              (early0_DivPlugin_logic_processing_div_io_cmd_valid               ), //i
    .io_cmd_ready              (early0_DivPlugin_logic_processing_div_io_cmd_ready               ), //o
    .io_cmd_payload_a          (early0_DivPlugin_logic_processing_a_delay_1[31:0]                ), //i
    .io_cmd_payload_b          (early0_DivPlugin_logic_processing_b_delay_1[31:0]                ), //i
    .io_cmd_payload_normalized (1'b0                                                             ), //i
    .io_cmd_payload_iterations (5'bxxxxx                                                         ), //i
    .io_rsp_valid              (early0_DivPlugin_logic_processing_div_io_rsp_valid               ), //o
    .io_rsp_ready              (1'b0                                                             ), //i
    .io_rsp_payload_result     (early0_DivPlugin_logic_processing_div_io_rsp_payload_result[31:0]), //o
    .io_rsp_payload_remain     (early0_DivPlugin_logic_processing_div_io_rsp_payload_remain[31:0]), //o
    .clk_cpu                   (clk_cpu                                                          ), //i
    .reset_cpu                 (reset_cpu                                                        )  //i
  );
  StreamArbiter LsuPlugin_logic_flusher_arbiter (
    .io_inputs_0_valid (TrapPlugin_logic_lsuL1Invalidate_0_cmd_valid     ), //i
    .io_inputs_0_ready (LsuPlugin_logic_flusher_arbiter_io_inputs_0_ready), //o
    .io_output_valid   (LsuPlugin_logic_flusher_arbiter_io_output_valid  ), //o
    .io_output_ready   (LsuPlugin_logic_flusher_arbiter_io_output_ready  ), //i
    .io_chosenOH       (LsuPlugin_logic_flusher_arbiter_io_chosenOH      ), //o
    .clk_cpu           (clk_cpu                                          ), //i
    .reset_cpu         (reset_cpu                                        )  //i
  );
  StreamArbiter_1 streamArbiter_10 (
    .io_inputs_0_valid                                     (late0_BranchPlugin_logic_jumpLogic_learn_m2sPipe_valid                                         ), //i
    .io_inputs_0_ready                                     (streamArbiter_10_io_inputs_0_ready                                                             ), //o
    .io_inputs_0_payload_pcOnLastSlice                     (late0_BranchPlugin_logic_jumpLogic_learn_m2sPipe_payload_pcOnLastSlice[31:0]                   ), //i
    .io_inputs_0_payload_pcTarget                          (late0_BranchPlugin_logic_jumpLogic_learn_m2sPipe_payload_pcTarget[31:0]                        ), //i
    .io_inputs_0_payload_taken                             (late0_BranchPlugin_logic_jumpLogic_learn_m2sPipe_payload_taken                                 ), //i
    .io_inputs_0_payload_isBranch                          (late0_BranchPlugin_logic_jumpLogic_learn_m2sPipe_payload_isBranch                              ), //i
    .io_inputs_0_payload_isPush                            (late0_BranchPlugin_logic_jumpLogic_learn_m2sPipe_payload_isPush                                ), //i
    .io_inputs_0_payload_isPop                             (late0_BranchPlugin_logic_jumpLogic_learn_m2sPipe_payload_isPop                                 ), //i
    .io_inputs_0_payload_wasWrong                          (late0_BranchPlugin_logic_jumpLogic_learn_m2sPipe_payload_wasWrong                              ), //i
    .io_inputs_0_payload_badPredictedTarget                (late0_BranchPlugin_logic_jumpLogic_learn_m2sPipe_payload_badPredictedTarget                    ), //i
    .io_inputs_0_payload_history                           (late0_BranchPlugin_logic_jumpLogic_learn_m2sPipe_payload_history[11:0]                         ), //i
    .io_inputs_0_payload_uopId                             (late0_BranchPlugin_logic_jumpLogic_learn_m2sPipe_payload_uopId[15:0]                           ), //i
    .io_inputs_0_payload_ctx_GSharePlugin_GSHARE_COUNTER_0 (late0_BranchPlugin_logic_jumpLogic_learn_m2sPipe_payload_ctx_GSharePlugin_GSHARE_COUNTER_0[1:0]), //i
    .io_inputs_0_payload_ctx_GSharePlugin_GSHARE_COUNTER_1 (late0_BranchPlugin_logic_jumpLogic_learn_m2sPipe_payload_ctx_GSharePlugin_GSHARE_COUNTER_1[1:0]), //i
    .io_inputs_0_payload_ctx_GSharePlugin_GSHARE_COUNTER_2 (late0_BranchPlugin_logic_jumpLogic_learn_m2sPipe_payload_ctx_GSharePlugin_GSHARE_COUNTER_2[1:0]), //i
    .io_inputs_0_payload_ctx_GSharePlugin_GSHARE_COUNTER_3 (late0_BranchPlugin_logic_jumpLogic_learn_m2sPipe_payload_ctx_GSharePlugin_GSHARE_COUNTER_3[1:0]), //i
    .io_inputs_1_valid                                     (late1_BranchPlugin_logic_jumpLogic_learn_m2sPipe_valid                                         ), //i
    .io_inputs_1_ready                                     (streamArbiter_10_io_inputs_1_ready                                                             ), //o
    .io_inputs_1_payload_pcOnLastSlice                     (late1_BranchPlugin_logic_jumpLogic_learn_m2sPipe_payload_pcOnLastSlice[31:0]                   ), //i
    .io_inputs_1_payload_pcTarget                          (late1_BranchPlugin_logic_jumpLogic_learn_m2sPipe_payload_pcTarget[31:0]                        ), //i
    .io_inputs_1_payload_taken                             (late1_BranchPlugin_logic_jumpLogic_learn_m2sPipe_payload_taken                                 ), //i
    .io_inputs_1_payload_isBranch                          (late1_BranchPlugin_logic_jumpLogic_learn_m2sPipe_payload_isBranch                              ), //i
    .io_inputs_1_payload_isPush                            (late1_BranchPlugin_logic_jumpLogic_learn_m2sPipe_payload_isPush                                ), //i
    .io_inputs_1_payload_isPop                             (late1_BranchPlugin_logic_jumpLogic_learn_m2sPipe_payload_isPop                                 ), //i
    .io_inputs_1_payload_wasWrong                          (late1_BranchPlugin_logic_jumpLogic_learn_m2sPipe_payload_wasWrong                              ), //i
    .io_inputs_1_payload_badPredictedTarget                (late1_BranchPlugin_logic_jumpLogic_learn_m2sPipe_payload_badPredictedTarget                    ), //i
    .io_inputs_1_payload_history                           (late1_BranchPlugin_logic_jumpLogic_learn_m2sPipe_payload_history[11:0]                         ), //i
    .io_inputs_1_payload_uopId                             (late1_BranchPlugin_logic_jumpLogic_learn_m2sPipe_payload_uopId[15:0]                           ), //i
    .io_inputs_1_payload_ctx_GSharePlugin_GSHARE_COUNTER_0 (late1_BranchPlugin_logic_jumpLogic_learn_m2sPipe_payload_ctx_GSharePlugin_GSHARE_COUNTER_0[1:0]), //i
    .io_inputs_1_payload_ctx_GSharePlugin_GSHARE_COUNTER_1 (late1_BranchPlugin_logic_jumpLogic_learn_m2sPipe_payload_ctx_GSharePlugin_GSHARE_COUNTER_1[1:0]), //i
    .io_inputs_1_payload_ctx_GSharePlugin_GSHARE_COUNTER_2 (late1_BranchPlugin_logic_jumpLogic_learn_m2sPipe_payload_ctx_GSharePlugin_GSHARE_COUNTER_2[1:0]), //i
    .io_inputs_1_payload_ctx_GSharePlugin_GSHARE_COUNTER_3 (late1_BranchPlugin_logic_jumpLogic_learn_m2sPipe_payload_ctx_GSharePlugin_GSHARE_COUNTER_3[1:0]), //i
    .io_output_valid                                       (streamArbiter_10_io_output_valid                                                               ), //o
    .io_output_ready                                       (streamArbiter_10_io_output_combStage_ready                                                     ), //i
    .io_output_payload_pcOnLastSlice                       (streamArbiter_10_io_output_payload_pcOnLastSlice[31:0]                                         ), //o
    .io_output_payload_pcTarget                            (streamArbiter_10_io_output_payload_pcTarget[31:0]                                              ), //o
    .io_output_payload_taken                               (streamArbiter_10_io_output_payload_taken                                                       ), //o
    .io_output_payload_isBranch                            (streamArbiter_10_io_output_payload_isBranch                                                    ), //o
    .io_output_payload_isPush                              (streamArbiter_10_io_output_payload_isPush                                                      ), //o
    .io_output_payload_isPop                               (streamArbiter_10_io_output_payload_isPop                                                       ), //o
    .io_output_payload_wasWrong                            (streamArbiter_10_io_output_payload_wasWrong                                                    ), //o
    .io_output_payload_badPredictedTarget                  (streamArbiter_10_io_output_payload_badPredictedTarget                                          ), //o
    .io_output_payload_history                             (streamArbiter_10_io_output_payload_history[11:0]                                               ), //o
    .io_output_payload_uopId                               (streamArbiter_10_io_output_payload_uopId[15:0]                                                 ), //o
    .io_output_payload_ctx_GSharePlugin_GSHARE_COUNTER_0   (streamArbiter_10_io_output_payload_ctx_GSharePlugin_GSHARE_COUNTER_0[1:0]                      ), //o
    .io_output_payload_ctx_GSharePlugin_GSHARE_COUNTER_1   (streamArbiter_10_io_output_payload_ctx_GSharePlugin_GSHARE_COUNTER_1[1:0]                      ), //o
    .io_output_payload_ctx_GSharePlugin_GSHARE_COUNTER_2   (streamArbiter_10_io_output_payload_ctx_GSharePlugin_GSHARE_COUNTER_2[1:0]                      ), //o
    .io_output_payload_ctx_GSharePlugin_GSHARE_COUNTER_3   (streamArbiter_10_io_output_payload_ctx_GSharePlugin_GSHARE_COUNTER_3[1:0]                      ), //o
    .io_chosen                                             (streamArbiter_10_io_chosen                                                                     ), //o
    .io_chosenOH                                           (streamArbiter_10_io_chosenOH[1:0]                                                              ), //o
    .clk_cpu                                               (clk_cpu                                                                                        ), //i
    .reset_cpu                                             (reset_cpu                                                                                      )  //i
  );
  StreamArbiter_2 LsuPlugin_logic_onAddress0_arbiter (
    .io_inputs_0_valid           (LsuPlugin_logic_onAddress0_ls_port_valid                          ), //i
    .io_inputs_0_ready           (LsuPlugin_logic_onAddress0_arbiter_io_inputs_0_ready              ), //o
    .io_inputs_0_payload_op      (LsuPlugin_logic_onAddress0_ls_port_payload_op[2:0]                ), //i
    .io_inputs_0_payload_address (LsuPlugin_logic_onAddress0_ls_port_payload_address[31:0]          ), //i
    .io_inputs_0_payload_size    (LsuPlugin_logic_onAddress0_ls_port_payload_size[1:0]              ), //i
    .io_inputs_0_payload_load    (LsuPlugin_logic_onAddress0_ls_port_payload_load                   ), //i
    .io_inputs_0_payload_store   (LsuPlugin_logic_onAddress0_ls_port_payload_store                  ), //i
    .io_inputs_0_payload_atomic  (LsuPlugin_logic_onAddress0_ls_port_payload_atomic                 ), //i
    .io_inputs_0_payload_storeId (LsuPlugin_logic_onAddress0_ls_port_payload_storeId[11:0]          ), //i
    .io_inputs_1_valid           (LsuPlugin_logic_onAddress0_access_port_valid                      ), //i
    .io_inputs_1_ready           (LsuPlugin_logic_onAddress0_arbiter_io_inputs_1_ready              ), //o
    .io_inputs_1_payload_op      (LsuPlugin_logic_onAddress0_access_port_payload_op[2:0]            ), //i
    .io_inputs_1_payload_address (LsuPlugin_logic_onAddress0_access_port_payload_address[31:0]      ), //i
    .io_inputs_1_payload_size    (LsuPlugin_logic_onAddress0_access_port_payload_size[1:0]          ), //i
    .io_inputs_1_payload_load    (LsuPlugin_logic_onAddress0_access_port_payload_load               ), //i
    .io_inputs_1_payload_store   (LsuPlugin_logic_onAddress0_access_port_payload_store              ), //i
    .io_inputs_1_payload_atomic  (LsuPlugin_logic_onAddress0_access_port_payload_atomic             ), //i
    .io_inputs_1_payload_storeId (LsuPlugin_logic_onAddress0_access_port_payload_storeId[11:0]      ), //i
    .io_inputs_2_valid           (LsuPlugin_logic_onAddress0_flush_port_valid                       ), //i
    .io_inputs_2_ready           (LsuPlugin_logic_onAddress0_arbiter_io_inputs_2_ready              ), //o
    .io_inputs_2_payload_op      (LsuPlugin_logic_onAddress0_flush_port_payload_op[2:0]             ), //i
    .io_inputs_2_payload_address (LsuPlugin_logic_onAddress0_flush_port_payload_address[31:0]       ), //i
    .io_inputs_2_payload_size    (LsuPlugin_logic_onAddress0_flush_port_payload_size[1:0]           ), //i
    .io_inputs_2_payload_load    (LsuPlugin_logic_onAddress0_flush_port_payload_load                ), //i
    .io_inputs_2_payload_store   (LsuPlugin_logic_onAddress0_flush_port_payload_store               ), //i
    .io_inputs_2_payload_atomic  (LsuPlugin_logic_onAddress0_flush_port_payload_atomic              ), //i
    .io_inputs_2_payload_storeId (LsuPlugin_logic_onAddress0_flush_port_payload_storeId[11:0]       ), //i
    .io_output_valid             (LsuPlugin_logic_onAddress0_arbiter_io_output_valid                ), //o
    .io_output_ready             (LsuPlugin_logic_onAddress0_arbiter_io_output_ready                ), //i
    .io_output_payload_op        (LsuPlugin_logic_onAddress0_arbiter_io_output_payload_op[2:0]      ), //o
    .io_output_payload_address   (LsuPlugin_logic_onAddress0_arbiter_io_output_payload_address[31:0]), //o
    .io_output_payload_size      (LsuPlugin_logic_onAddress0_arbiter_io_output_payload_size[1:0]    ), //o
    .io_output_payload_load      (LsuPlugin_logic_onAddress0_arbiter_io_output_payload_load         ), //o
    .io_output_payload_store     (LsuPlugin_logic_onAddress0_arbiter_io_output_payload_store        ), //o
    .io_output_payload_atomic    (LsuPlugin_logic_onAddress0_arbiter_io_output_payload_atomic       ), //o
    .io_output_payload_storeId   (LsuPlugin_logic_onAddress0_arbiter_io_output_payload_storeId[11:0]), //o
    .io_chosen                   (LsuPlugin_logic_onAddress0_arbiter_io_chosen[1:0]                 ), //o
    .io_chosenOH                 (LsuPlugin_logic_onAddress0_arbiter_io_chosenOH[2:0]               ), //o
    .clk_cpu                     (clk_cpu                                                           ), //i
    .reset_cpu                   (reset_cpu                                                         )  //i
  );
  StreamArbiter_3 MmuPlugin_logic_refill_arbiter (
    .io_inputs_0_valid             (TrapPlugin_logic_harts_0_trap_fsm_atsPorts_refill_cmd_valid                ), //i
    .io_inputs_0_ready             (MmuPlugin_logic_refill_arbiter_io_inputs_0_ready                           ), //o
    .io_inputs_0_payload_address   (TrapPlugin_logic_harts_0_trap_fsm_atsPorts_refill_cmd_payload_address[31:0]), //i
    .io_inputs_0_payload_storageId (TrapPlugin_logic_harts_0_trap_fsm_atsPorts_refill_cmd_payload_storageId    ), //i
    .io_output_valid               (MmuPlugin_logic_refill_arbiter_io_output_valid                             ), //o
    .io_output_ready               (MmuPlugin_logic_refill_arbiter_io_output_ready                             ), //i
    .io_output_payload_address     (MmuPlugin_logic_refill_arbiter_io_output_payload_address[31:0]             ), //o
    .io_output_payload_storageId   (MmuPlugin_logic_refill_arbiter_io_output_payload_storageId                 ), //o
    .io_chosenOH                   (MmuPlugin_logic_refill_arbiter_io_chosenOH                                 ), //o
    .clk_cpu                       (clk_cpu                                                                    ), //i
    .reset_cpu                     (reset_cpu                                                                  )  //i
  );
  StreamArbiter_4 MmuPlugin_logic_invalidate_arbiter (
    .io_inputs_0_valid (TrapPlugin_logic_harts_0_trap_fsm_atsPorts_invalidate_cmd_valid), //i
    .io_inputs_0_ready (MmuPlugin_logic_invalidate_arbiter_io_inputs_0_ready           ), //o
    .io_output_valid   (MmuPlugin_logic_invalidate_arbiter_io_output_valid             ), //o
    .io_output_ready   (MmuPlugin_logic_invalidate_arbiter_io_output_ready             ), //i
    .io_chosenOH       (MmuPlugin_logic_invalidate_arbiter_io_chosenOH                 ), //o
    .clk_cpu           (clk_cpu                                                        ), //i
    .reset_cpu         (reset_cpu                                                      )  //i
  );
  RegFileMem integer_RegFilePlugin_logic_regfile_fpga (
    .io_writes_0_valid   (integer_RegFilePlugin_logic_regfile_fpga_io_writes_0_valid       ), //i
    .io_writes_0_address (integer_RegFilePlugin_logic_regfile_fpga_io_writes_0_address[4:0]), //i
    .io_writes_0_data    (integer_RegFilePlugin_logic_regfile_fpga_io_writes_0_data[31:0]  ), //i
    .io_writes_0_uopId   (integer_RegFilePlugin_logic_writeMerges_0_bus_uopId[15:0]        ), //i
    .io_writes_1_valid   (integer_RegFilePlugin_logic_writeMerges_1_bus_valid              ), //i
    .io_writes_1_address (integer_RegFilePlugin_logic_writeMerges_1_bus_address[4:0]       ), //i
    .io_writes_1_data    (integer_RegFilePlugin_logic_writeMerges_1_bus_data[31:0]         ), //i
    .io_writes_1_uopId   (integer_RegFilePlugin_logic_writeMerges_1_bus_uopId[15:0]        ), //i
    .io_reads_0_valid    (toplevel_execute_lane1_bypasser_integer_RS1_port_valid           ), //i
    .io_reads_0_address  (toplevel_execute_lane1_bypasser_integer_RS1_port_address[4:0]    ), //i
    .io_reads_0_data     (integer_RegFilePlugin_logic_regfile_fpga_io_reads_0_data[31:0]   ), //o
    .io_reads_1_valid    (toplevel_execute_lane0_bypasser_integer_RS1_port_valid           ), //i
    .io_reads_1_address  (toplevel_execute_lane0_bypasser_integer_RS1_port_address[4:0]    ), //i
    .io_reads_1_data     (integer_RegFilePlugin_logic_regfile_fpga_io_reads_1_data[31:0]   ), //o
    .io_reads_2_valid    (toplevel_execute_lane0_bypasser_integer_RS2_port_valid           ), //i
    .io_reads_2_address  (toplevel_execute_lane0_bypasser_integer_RS2_port_address[4:0]    ), //i
    .io_reads_2_data     (integer_RegFilePlugin_logic_regfile_fpga_io_reads_2_data[31:0]   ), //o
    .io_reads_3_valid    (toplevel_execute_lane1_bypasser_integer_RS2_port_valid           ), //i
    .io_reads_3_address  (toplevel_execute_lane1_bypasser_integer_RS2_port_address[4:0]    ), //i
    .io_reads_3_data     (integer_RegFilePlugin_logic_regfile_fpga_io_reads_3_data[31:0]   ), //o
    .clk_cpu             (clk_cpu                                                          ), //i
    .reset_cpu           (reset_cpu                                                        )  //i
  );
  always @(*) begin
    case(_zz_fetch_logic_ctrls_2_down_AlignerPlugin_logic_FETCH_MASK_1)
      2'b00 : _zz_fetch_logic_ctrls_2_down_AlignerPlugin_logic_FETCH_MASK = AlignerPlugin_logic_maskGen_frontMasks_0;
      2'b01 : _zz_fetch_logic_ctrls_2_down_AlignerPlugin_logic_FETCH_MASK = AlignerPlugin_logic_maskGen_frontMasks_1;
      2'b10 : _zz_fetch_logic_ctrls_2_down_AlignerPlugin_logic_FETCH_MASK = AlignerPlugin_logic_maskGen_frontMasks_2;
      default : _zz_fetch_logic_ctrls_2_down_AlignerPlugin_logic_FETCH_MASK = AlignerPlugin_logic_maskGen_frontMasks_3;
    endcase
  end

  always @(*) begin
    case(fetch_logic_ctrls_2_down_Prediction_WORD_JUMP_SLICE)
      2'b00 : _zz_fetch_logic_ctrls_2_down_AlignerPlugin_logic_FETCH_MASK_2 = AlignerPlugin_logic_maskGen_backMasks_0;
      2'b01 : _zz_fetch_logic_ctrls_2_down_AlignerPlugin_logic_FETCH_MASK_2 = AlignerPlugin_logic_maskGen_backMasks_1;
      2'b10 : _zz_fetch_logic_ctrls_2_down_AlignerPlugin_logic_FETCH_MASK_2 = AlignerPlugin_logic_maskGen_backMasks_2;
      default : _zz_fetch_logic_ctrls_2_down_AlignerPlugin_logic_FETCH_MASK_2 = AlignerPlugin_logic_maskGen_backMasks_3;
    endcase
  end

  always @(*) begin
    case(_zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_28)
      2'b00 : _zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_27 = _zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_22;
      2'b01 : _zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_27 = (_zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_22 | 32'h40000000);
      2'b10 : _zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_27 = {{{{_zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_5,_zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst},3'b111},_zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst},7'h13};
      default : _zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_27 = ({{{{{7'h0,_zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_1},_zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst},_zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_29},_zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst},(AlignerPlugin_logic_extractors_0_ctx_instruction[12] ? 7'h3b : 7'h33)} | ((AlignerPlugin_logic_extractors_0_ctx_instruction[6 : 5] == 2'b00) ? 32'h40000000 : 32'h0));
    endcase
  end

  always @(*) begin
    case(_zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_30)
      3'b000 : _zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_29 = 3'b000;
      3'b001 : _zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_29 = 3'b100;
      3'b010 : _zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_29 = 3'b110;
      3'b011 : _zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_29 = 3'b111;
      3'b100 : _zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_29 = 3'b000;
      3'b101 : _zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_29 = 3'b000;
      3'b110 : _zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_29 = 3'b010;
      default : _zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_29 = 3'b011;
    endcase
  end

  always @(*) begin
    case(_zz_AlignerPlugin_logic_feeder_lanes_1_withRvc_dec_inst_28)
      2'b00 : _zz_AlignerPlugin_logic_feeder_lanes_1_withRvc_dec_inst_27 = _zz_AlignerPlugin_logic_feeder_lanes_1_withRvc_dec_inst_22;
      2'b01 : _zz_AlignerPlugin_logic_feeder_lanes_1_withRvc_dec_inst_27 = (_zz_AlignerPlugin_logic_feeder_lanes_1_withRvc_dec_inst_22 | 32'h40000000);
      2'b10 : _zz_AlignerPlugin_logic_feeder_lanes_1_withRvc_dec_inst_27 = {{{{_zz_AlignerPlugin_logic_feeder_lanes_1_withRvc_dec_inst_5,_zz_AlignerPlugin_logic_feeder_lanes_1_withRvc_dec_inst},3'b111},_zz_AlignerPlugin_logic_feeder_lanes_1_withRvc_dec_inst},7'h13};
      default : _zz_AlignerPlugin_logic_feeder_lanes_1_withRvc_dec_inst_27 = ({{{{{7'h0,_zz_AlignerPlugin_logic_feeder_lanes_1_withRvc_dec_inst_1},_zz_AlignerPlugin_logic_feeder_lanes_1_withRvc_dec_inst},_zz_AlignerPlugin_logic_feeder_lanes_1_withRvc_dec_inst_29},_zz_AlignerPlugin_logic_feeder_lanes_1_withRvc_dec_inst},(AlignerPlugin_logic_extractors_1_ctx_instruction[12] ? 7'h3b : 7'h33)} | ((AlignerPlugin_logic_extractors_1_ctx_instruction[6 : 5] == 2'b00) ? 32'h40000000 : 32'h0));
    endcase
  end

  always @(*) begin
    case(_zz_AlignerPlugin_logic_feeder_lanes_1_withRvc_dec_inst_30)
      3'b000 : _zz_AlignerPlugin_logic_feeder_lanes_1_withRvc_dec_inst_29 = 3'b000;
      3'b001 : _zz_AlignerPlugin_logic_feeder_lanes_1_withRvc_dec_inst_29 = 3'b100;
      3'b010 : _zz_AlignerPlugin_logic_feeder_lanes_1_withRvc_dec_inst_29 = 3'b110;
      3'b011 : _zz_AlignerPlugin_logic_feeder_lanes_1_withRvc_dec_inst_29 = 3'b111;
      3'b100 : _zz_AlignerPlugin_logic_feeder_lanes_1_withRvc_dec_inst_29 = 3'b000;
      3'b101 : _zz_AlignerPlugin_logic_feeder_lanes_1_withRvc_dec_inst_29 = 3'b000;
      3'b110 : _zz_AlignerPlugin_logic_feeder_lanes_1_withRvc_dec_inst_29 = 3'b010;
      default : _zz_AlignerPlugin_logic_feeder_lanes_1_withRvc_dec_inst_29 = 3'b011;
    endcase
  end

  always @(*) begin
    case(_zz_DispatchPlugin_logic_candidates_1_age_1)
      1'b0 : _zz_DispatchPlugin_logic_candidates_1_age = 1'b0;
      default : _zz_DispatchPlugin_logic_candidates_1_age = 1'b1;
    endcase
  end

  always @(*) begin
    case(_zz_DispatchPlugin_logic_candidates_2_age_1)
      2'b00 : _zz_DispatchPlugin_logic_candidates_2_age = 2'b00;
      2'b01 : _zz_DispatchPlugin_logic_candidates_2_age = 2'b01;
      2'b10 : _zz_DispatchPlugin_logic_candidates_2_age = 2'b01;
      default : _zz_DispatchPlugin_logic_candidates_2_age = 2'b10;
    endcase
  end

  always @(*) begin
    case(_zz_DispatchPlugin_logic_slotsFeeds_fit_1)
      2'b00 : _zz_DispatchPlugin_logic_slotsFeeds_fit = 2'b00;
      2'b01 : _zz_DispatchPlugin_logic_slotsFeeds_fit = 2'b01;
      2'b10 : _zz_DispatchPlugin_logic_slotsFeeds_fit = 2'b01;
      default : _zz_DispatchPlugin_logic_slotsFeeds_fit = 2'b10;
    endcase
  end

  always @(*) begin
    case(LsuL1Plugin_logic_writeback_read_slotReadLast_payload_way)
      1'b0 : _zz_LsuL1Plugin_logic_writeback_read_readedData = LsuL1Plugin_logic_banks_0_read_rsp;
      default : _zz_LsuL1Plugin_logic_writeback_read_readedData = LsuL1Plugin_logic_banks_1_read_rsp;
    endcase
  end

  always @(*) begin
    case(_zz_toplevel_execute_ctrl3_down_LsuL1Plugin_logic_BANKS_MUXES_lane0_0_1)
      1'b0 : _zz_toplevel_execute_ctrl3_down_LsuL1Plugin_logic_BANKS_MUXES_lane0_0 = toplevel_execute_ctrl3_down_LsuL1Plugin_logic_BANKS_WORDS_lane0_0[31 : 0];
      default : _zz_toplevel_execute_ctrl3_down_LsuL1Plugin_logic_BANKS_MUXES_lane0_0 = toplevel_execute_ctrl3_down_LsuL1Plugin_logic_BANKS_WORDS_lane0_0[63 : 32];
    endcase
  end

  always @(*) begin
    case(_zz_toplevel_execute_ctrl3_down_LsuL1Plugin_logic_BANKS_MUXES_lane0_1_1)
      1'b0 : _zz_toplevel_execute_ctrl3_down_LsuL1Plugin_logic_BANKS_MUXES_lane0_1 = toplevel_execute_ctrl3_down_LsuL1Plugin_logic_BANKS_WORDS_lane0_1[31 : 0];
      default : _zz_toplevel_execute_ctrl3_down_LsuL1Plugin_logic_BANKS_MUXES_lane0_1 = toplevel_execute_ctrl3_down_LsuL1Plugin_logic_BANKS_WORDS_lane0_1[63 : 32];
    endcase
  end

  always @(*) begin
    case(_zz_56)
      2'b00 : _zz_55 = 2'b00;
      2'b01 : _zz_55 = 2'b01;
      2'b10 : _zz_55 = 2'b01;
      default : _zz_55 = 2'b10;
    endcase
  end

  always @(*) begin
    case(_zz_58)
      3'b000 : _zz_57 = 2'b00;
      3'b001 : _zz_57 = 2'b01;
      3'b010 : _zz_57 = 2'b01;
      3'b011 : _zz_57 = 2'b10;
      3'b100 : _zz_57 = 2'b01;
      3'b101 : _zz_57 = 2'b10;
      3'b110 : _zz_57 = 2'b10;
      default : _zz_57 = 2'b11;
    endcase
  end

  always @(*) begin
    case(LsuL1Plugin_logic_ls_ctrl_needFlushSel)
      1'b0 : begin
        _zz__zz_LsuL1Plugin_logic_waysWrite_tag_address = toplevel_execute_ctrl4_down_LsuL1Plugin_logic_WAYS_TAGS_lane0_0_address;
        _zz_LsuL1Plugin_logic_waysWrite_tag_fault = toplevel_execute_ctrl4_down_LsuL1Plugin_logic_WAYS_TAGS_lane0_0_fault;
      end
      default : begin
        _zz__zz_LsuL1Plugin_logic_waysWrite_tag_address = toplevel_execute_ctrl4_down_LsuL1Plugin_logic_WAYS_TAGS_lane0_1_address;
        _zz_LsuL1Plugin_logic_waysWrite_tag_fault = toplevel_execute_ctrl4_down_LsuL1Plugin_logic_WAYS_TAGS_lane0_1_fault;
      end
    endcase
  end

  always @(*) begin
    case(LsuL1Plugin_logic_ls_ctrl_targetWay)
      1'b0 : _zz_LsuL1Plugin_logic_writeback_push_payload_address = toplevel_execute_ctrl4_down_LsuL1Plugin_logic_WAYS_TAGS_lane0_0_address;
      default : _zz_LsuL1Plugin_logic_writeback_push_payload_address = toplevel_execute_ctrl4_down_LsuL1Plugin_logic_WAYS_TAGS_lane0_1_address;
    endcase
  end

  always @(*) begin
    case(_zz_LsuPlugin_logic_onCtrl_loadData_shited_1)
      2'b00 : _zz_LsuPlugin_logic_onCtrl_loadData_shited = LsuPlugin_logic_onCtrl_loadData_splited_0;
      2'b01 : _zz_LsuPlugin_logic_onCtrl_loadData_shited = LsuPlugin_logic_onCtrl_loadData_splited_1;
      2'b10 : _zz_LsuPlugin_logic_onCtrl_loadData_shited = LsuPlugin_logic_onCtrl_loadData_splited_2;
      default : _zz_LsuPlugin_logic_onCtrl_loadData_shited = LsuPlugin_logic_onCtrl_loadData_splited_3;
    endcase
  end

  always @(*) begin
    case(_zz_LsuPlugin_logic_onCtrl_loadData_shited_3)
      1'b0 : _zz_LsuPlugin_logic_onCtrl_loadData_shited_2 = LsuPlugin_logic_onCtrl_loadData_splited_1;
      default : _zz_LsuPlugin_logic_onCtrl_loadData_shited_2 = LsuPlugin_logic_onCtrl_loadData_splited_3;
    endcase
  end

  always @(*) begin
    case(LsuL1TileLinkPlugin_logic_down_a_payload_size)
      3'b000 : _zz_LsuL1TileLinkPlugin_logic_down_a_tracker_last = 3'b000;
      3'b001 : _zz_LsuL1TileLinkPlugin_logic_down_a_tracker_last = 3'b000;
      3'b010 : _zz_LsuL1TileLinkPlugin_logic_down_a_tracker_last = 3'b000;
      3'b011 : _zz_LsuL1TileLinkPlugin_logic_down_a_tracker_last = 3'b000;
      3'b100 : _zz_LsuL1TileLinkPlugin_logic_down_a_tracker_last = 3'b001;
      3'b101 : _zz_LsuL1TileLinkPlugin_logic_down_a_tracker_last = 3'b011;
      default : _zz_LsuL1TileLinkPlugin_logic_down_a_tracker_last = 3'b111;
    endcase
  end

  always @(*) begin
    case(CsrRamPlugin_logic_readLogic_sel)
      1'b0 : _zz_CsrRamPlugin_logic_readLogic_port_cmd_payload = TrapPlugin_logic_harts_0_crsPorts_read_address;
      default : _zz_CsrRamPlugin_logic_readLogic_port_cmd_payload = CsrRamPlugin_csrMapper_read_address;
    endcase
  end

  always @(*) begin
    case(_zz_WhiteboxerPlugin_logic_perf_candidatesCount_1)
      3'b000 : _zz_WhiteboxerPlugin_logic_perf_candidatesCount = 2'b00;
      3'b001 : _zz_WhiteboxerPlugin_logic_perf_candidatesCount = 2'b01;
      3'b010 : _zz_WhiteboxerPlugin_logic_perf_candidatesCount = 2'b01;
      3'b011 : _zz_WhiteboxerPlugin_logic_perf_candidatesCount = 2'b10;
      3'b100 : _zz_WhiteboxerPlugin_logic_perf_candidatesCount = 2'b01;
      3'b101 : _zz_WhiteboxerPlugin_logic_perf_candidatesCount = 2'b10;
      3'b110 : _zz_WhiteboxerPlugin_logic_perf_candidatesCount = 2'b10;
      default : _zz_WhiteboxerPlugin_logic_perf_candidatesCount = 2'b11;
    endcase
  end

  always @(*) begin
    case(_zz_WhiteboxerPlugin_logic_perf_dispatchFeedCount_1)
      2'b00 : _zz_WhiteboxerPlugin_logic_perf_dispatchFeedCount = 2'b00;
      2'b01 : _zz_WhiteboxerPlugin_logic_perf_dispatchFeedCount = 2'b01;
      2'b10 : _zz_WhiteboxerPlugin_logic_perf_dispatchFeedCount = 2'b01;
      default : _zz_WhiteboxerPlugin_logic_perf_dispatchFeedCount = 2'b10;
    endcase
  end

  `ifndef SYNTHESIS
  always @(*) begin
    case(toplevel_execute_ctrl3_down_late1_IntAluPlugin_ALU_BITWISE_CTRL_lane1)
      IntAluPlugin_AluBitwiseCtrlEnum_XOR_1 : toplevel_execute_ctrl3_down_late1_IntAluPlugin_ALU_BITWISE_CTRL_lane1_string = "XOR_1";
      IntAluPlugin_AluBitwiseCtrlEnum_OR_1 : toplevel_execute_ctrl3_down_late1_IntAluPlugin_ALU_BITWISE_CTRL_lane1_string = "OR_1 ";
      IntAluPlugin_AluBitwiseCtrlEnum_AND_1 : toplevel_execute_ctrl3_down_late1_IntAluPlugin_ALU_BITWISE_CTRL_lane1_string = "AND_1";
      IntAluPlugin_AluBitwiseCtrlEnum_ZERO : toplevel_execute_ctrl3_down_late1_IntAluPlugin_ALU_BITWISE_CTRL_lane1_string = "ZERO ";
      default : toplevel_execute_ctrl3_down_late1_IntAluPlugin_ALU_BITWISE_CTRL_lane1_string = "?????";
    endcase
  end
  always @(*) begin
    case(toplevel_execute_ctrl3_down_late0_IntAluPlugin_ALU_BITWISE_CTRL_lane0)
      IntAluPlugin_AluBitwiseCtrlEnum_XOR_1 : toplevel_execute_ctrl3_down_late0_IntAluPlugin_ALU_BITWISE_CTRL_lane0_string = "XOR_1";
      IntAluPlugin_AluBitwiseCtrlEnum_OR_1 : toplevel_execute_ctrl3_down_late0_IntAluPlugin_ALU_BITWISE_CTRL_lane0_string = "OR_1 ";
      IntAluPlugin_AluBitwiseCtrlEnum_AND_1 : toplevel_execute_ctrl3_down_late0_IntAluPlugin_ALU_BITWISE_CTRL_lane0_string = "AND_1";
      IntAluPlugin_AluBitwiseCtrlEnum_ZERO : toplevel_execute_ctrl3_down_late0_IntAluPlugin_ALU_BITWISE_CTRL_lane0_string = "ZERO ";
      default : toplevel_execute_ctrl3_down_late0_IntAluPlugin_ALU_BITWISE_CTRL_lane0_string = "?????";
    endcase
  end
  always @(*) begin
    case(toplevel_execute_ctrl4_up_late1_IntAluPlugin_ALU_BITWISE_CTRL_lane1)
      IntAluPlugin_AluBitwiseCtrlEnum_XOR_1 : toplevel_execute_ctrl4_up_late1_IntAluPlugin_ALU_BITWISE_CTRL_lane1_string = "XOR_1";
      IntAluPlugin_AluBitwiseCtrlEnum_OR_1 : toplevel_execute_ctrl4_up_late1_IntAluPlugin_ALU_BITWISE_CTRL_lane1_string = "OR_1 ";
      IntAluPlugin_AluBitwiseCtrlEnum_AND_1 : toplevel_execute_ctrl4_up_late1_IntAluPlugin_ALU_BITWISE_CTRL_lane1_string = "AND_1";
      IntAluPlugin_AluBitwiseCtrlEnum_ZERO : toplevel_execute_ctrl4_up_late1_IntAluPlugin_ALU_BITWISE_CTRL_lane1_string = "ZERO ";
      default : toplevel_execute_ctrl4_up_late1_IntAluPlugin_ALU_BITWISE_CTRL_lane1_string = "?????";
    endcase
  end
  always @(*) begin
    case(toplevel_execute_ctrl4_up_BranchPlugin_BRANCH_CTRL_lane1)
      BranchPlugin_BranchCtrlEnum_B : toplevel_execute_ctrl4_up_BranchPlugin_BRANCH_CTRL_lane1_string = "B   ";
      BranchPlugin_BranchCtrlEnum_JAL : toplevel_execute_ctrl4_up_BranchPlugin_BRANCH_CTRL_lane1_string = "JAL ";
      BranchPlugin_BranchCtrlEnum_JALR : toplevel_execute_ctrl4_up_BranchPlugin_BRANCH_CTRL_lane1_string = "JALR";
      default : toplevel_execute_ctrl4_up_BranchPlugin_BRANCH_CTRL_lane1_string = "????";
    endcase
  end
  always @(*) begin
    case(toplevel_execute_ctrl4_up_late0_IntAluPlugin_ALU_BITWISE_CTRL_lane0)
      IntAluPlugin_AluBitwiseCtrlEnum_XOR_1 : toplevel_execute_ctrl4_up_late0_IntAluPlugin_ALU_BITWISE_CTRL_lane0_string = "XOR_1";
      IntAluPlugin_AluBitwiseCtrlEnum_OR_1 : toplevel_execute_ctrl4_up_late0_IntAluPlugin_ALU_BITWISE_CTRL_lane0_string = "OR_1 ";
      IntAluPlugin_AluBitwiseCtrlEnum_AND_1 : toplevel_execute_ctrl4_up_late0_IntAluPlugin_ALU_BITWISE_CTRL_lane0_string = "AND_1";
      IntAluPlugin_AluBitwiseCtrlEnum_ZERO : toplevel_execute_ctrl4_up_late0_IntAluPlugin_ALU_BITWISE_CTRL_lane0_string = "ZERO ";
      default : toplevel_execute_ctrl4_up_late0_IntAluPlugin_ALU_BITWISE_CTRL_lane0_string = "?????";
    endcase
  end
  always @(*) begin
    case(toplevel_execute_ctrl4_up_BranchPlugin_BRANCH_CTRL_lane0)
      BranchPlugin_BranchCtrlEnum_B : toplevel_execute_ctrl4_up_BranchPlugin_BRANCH_CTRL_lane0_string = "B   ";
      BranchPlugin_BranchCtrlEnum_JAL : toplevel_execute_ctrl4_up_BranchPlugin_BRANCH_CTRL_lane0_string = "JAL ";
      BranchPlugin_BranchCtrlEnum_JALR : toplevel_execute_ctrl4_up_BranchPlugin_BRANCH_CTRL_lane0_string = "JALR";
      default : toplevel_execute_ctrl4_up_BranchPlugin_BRANCH_CTRL_lane0_string = "????";
    endcase
  end
  always @(*) begin
    case(toplevel_execute_ctrl2_down_late1_IntAluPlugin_ALU_BITWISE_CTRL_lane1)
      IntAluPlugin_AluBitwiseCtrlEnum_XOR_1 : toplevel_execute_ctrl2_down_late1_IntAluPlugin_ALU_BITWISE_CTRL_lane1_string = "XOR_1";
      IntAluPlugin_AluBitwiseCtrlEnum_OR_1 : toplevel_execute_ctrl2_down_late1_IntAluPlugin_ALU_BITWISE_CTRL_lane1_string = "OR_1 ";
      IntAluPlugin_AluBitwiseCtrlEnum_AND_1 : toplevel_execute_ctrl2_down_late1_IntAluPlugin_ALU_BITWISE_CTRL_lane1_string = "AND_1";
      IntAluPlugin_AluBitwiseCtrlEnum_ZERO : toplevel_execute_ctrl2_down_late1_IntAluPlugin_ALU_BITWISE_CTRL_lane1_string = "ZERO ";
      default : toplevel_execute_ctrl2_down_late1_IntAluPlugin_ALU_BITWISE_CTRL_lane1_string = "?????";
    endcase
  end
  always @(*) begin
    case(toplevel_execute_ctrl2_down_late0_IntAluPlugin_ALU_BITWISE_CTRL_lane0)
      IntAluPlugin_AluBitwiseCtrlEnum_XOR_1 : toplevel_execute_ctrl2_down_late0_IntAluPlugin_ALU_BITWISE_CTRL_lane0_string = "XOR_1";
      IntAluPlugin_AluBitwiseCtrlEnum_OR_1 : toplevel_execute_ctrl2_down_late0_IntAluPlugin_ALU_BITWISE_CTRL_lane0_string = "OR_1 ";
      IntAluPlugin_AluBitwiseCtrlEnum_AND_1 : toplevel_execute_ctrl2_down_late0_IntAluPlugin_ALU_BITWISE_CTRL_lane0_string = "AND_1";
      IntAluPlugin_AluBitwiseCtrlEnum_ZERO : toplevel_execute_ctrl2_down_late0_IntAluPlugin_ALU_BITWISE_CTRL_lane0_string = "ZERO ";
      default : toplevel_execute_ctrl2_down_late0_IntAluPlugin_ALU_BITWISE_CTRL_lane0_string = "?????";
    endcase
  end
  always @(*) begin
    case(toplevel_execute_ctrl3_up_late1_IntAluPlugin_ALU_BITWISE_CTRL_lane1)
      IntAluPlugin_AluBitwiseCtrlEnum_XOR_1 : toplevel_execute_ctrl3_up_late1_IntAluPlugin_ALU_BITWISE_CTRL_lane1_string = "XOR_1";
      IntAluPlugin_AluBitwiseCtrlEnum_OR_1 : toplevel_execute_ctrl3_up_late1_IntAluPlugin_ALU_BITWISE_CTRL_lane1_string = "OR_1 ";
      IntAluPlugin_AluBitwiseCtrlEnum_AND_1 : toplevel_execute_ctrl3_up_late1_IntAluPlugin_ALU_BITWISE_CTRL_lane1_string = "AND_1";
      IntAluPlugin_AluBitwiseCtrlEnum_ZERO : toplevel_execute_ctrl3_up_late1_IntAluPlugin_ALU_BITWISE_CTRL_lane1_string = "ZERO ";
      default : toplevel_execute_ctrl3_up_late1_IntAluPlugin_ALU_BITWISE_CTRL_lane1_string = "?????";
    endcase
  end
  always @(*) begin
    case(toplevel_execute_ctrl3_up_BranchPlugin_BRANCH_CTRL_lane1)
      BranchPlugin_BranchCtrlEnum_B : toplevel_execute_ctrl3_up_BranchPlugin_BRANCH_CTRL_lane1_string = "B   ";
      BranchPlugin_BranchCtrlEnum_JAL : toplevel_execute_ctrl3_up_BranchPlugin_BRANCH_CTRL_lane1_string = "JAL ";
      BranchPlugin_BranchCtrlEnum_JALR : toplevel_execute_ctrl3_up_BranchPlugin_BRANCH_CTRL_lane1_string = "JALR";
      default : toplevel_execute_ctrl3_up_BranchPlugin_BRANCH_CTRL_lane1_string = "????";
    endcase
  end
  always @(*) begin
    case(toplevel_execute_ctrl3_up_late0_IntAluPlugin_ALU_BITWISE_CTRL_lane0)
      IntAluPlugin_AluBitwiseCtrlEnum_XOR_1 : toplevel_execute_ctrl3_up_late0_IntAluPlugin_ALU_BITWISE_CTRL_lane0_string = "XOR_1";
      IntAluPlugin_AluBitwiseCtrlEnum_OR_1 : toplevel_execute_ctrl3_up_late0_IntAluPlugin_ALU_BITWISE_CTRL_lane0_string = "OR_1 ";
      IntAluPlugin_AluBitwiseCtrlEnum_AND_1 : toplevel_execute_ctrl3_up_late0_IntAluPlugin_ALU_BITWISE_CTRL_lane0_string = "AND_1";
      IntAluPlugin_AluBitwiseCtrlEnum_ZERO : toplevel_execute_ctrl3_up_late0_IntAluPlugin_ALU_BITWISE_CTRL_lane0_string = "ZERO ";
      default : toplevel_execute_ctrl3_up_late0_IntAluPlugin_ALU_BITWISE_CTRL_lane0_string = "?????";
    endcase
  end
  always @(*) begin
    case(toplevel_execute_ctrl3_up_BranchPlugin_BRANCH_CTRL_lane0)
      BranchPlugin_BranchCtrlEnum_B : toplevel_execute_ctrl3_up_BranchPlugin_BRANCH_CTRL_lane0_string = "B   ";
      BranchPlugin_BranchCtrlEnum_JAL : toplevel_execute_ctrl3_up_BranchPlugin_BRANCH_CTRL_lane0_string = "JAL ";
      BranchPlugin_BranchCtrlEnum_JALR : toplevel_execute_ctrl3_up_BranchPlugin_BRANCH_CTRL_lane0_string = "JALR";
      default : toplevel_execute_ctrl3_up_BranchPlugin_BRANCH_CTRL_lane0_string = "????";
    endcase
  end
  always @(*) begin
    case(toplevel_execute_ctrl2_up_late1_IntAluPlugin_ALU_BITWISE_CTRL_lane1)
      IntAluPlugin_AluBitwiseCtrlEnum_XOR_1 : toplevel_execute_ctrl2_up_late1_IntAluPlugin_ALU_BITWISE_CTRL_lane1_string = "XOR_1";
      IntAluPlugin_AluBitwiseCtrlEnum_OR_1 : toplevel_execute_ctrl2_up_late1_IntAluPlugin_ALU_BITWISE_CTRL_lane1_string = "OR_1 ";
      IntAluPlugin_AluBitwiseCtrlEnum_AND_1 : toplevel_execute_ctrl2_up_late1_IntAluPlugin_ALU_BITWISE_CTRL_lane1_string = "AND_1";
      IntAluPlugin_AluBitwiseCtrlEnum_ZERO : toplevel_execute_ctrl2_up_late1_IntAluPlugin_ALU_BITWISE_CTRL_lane1_string = "ZERO ";
      default : toplevel_execute_ctrl2_up_late1_IntAluPlugin_ALU_BITWISE_CTRL_lane1_string = "?????";
    endcase
  end
  always @(*) begin
    case(toplevel_execute_ctrl2_up_BranchPlugin_BRANCH_CTRL_lane1)
      BranchPlugin_BranchCtrlEnum_B : toplevel_execute_ctrl2_up_BranchPlugin_BRANCH_CTRL_lane1_string = "B   ";
      BranchPlugin_BranchCtrlEnum_JAL : toplevel_execute_ctrl2_up_BranchPlugin_BRANCH_CTRL_lane1_string = "JAL ";
      BranchPlugin_BranchCtrlEnum_JALR : toplevel_execute_ctrl2_up_BranchPlugin_BRANCH_CTRL_lane1_string = "JALR";
      default : toplevel_execute_ctrl2_up_BranchPlugin_BRANCH_CTRL_lane1_string = "????";
    endcase
  end
  always @(*) begin
    case(toplevel_execute_ctrl2_up_early1_IntAluPlugin_ALU_BITWISE_CTRL_lane1)
      IntAluPlugin_AluBitwiseCtrlEnum_XOR_1 : toplevel_execute_ctrl2_up_early1_IntAluPlugin_ALU_BITWISE_CTRL_lane1_string = "XOR_1";
      IntAluPlugin_AluBitwiseCtrlEnum_OR_1 : toplevel_execute_ctrl2_up_early1_IntAluPlugin_ALU_BITWISE_CTRL_lane1_string = "OR_1 ";
      IntAluPlugin_AluBitwiseCtrlEnum_AND_1 : toplevel_execute_ctrl2_up_early1_IntAluPlugin_ALU_BITWISE_CTRL_lane1_string = "AND_1";
      IntAluPlugin_AluBitwiseCtrlEnum_ZERO : toplevel_execute_ctrl2_up_early1_IntAluPlugin_ALU_BITWISE_CTRL_lane1_string = "ZERO ";
      default : toplevel_execute_ctrl2_up_early1_IntAluPlugin_ALU_BITWISE_CTRL_lane1_string = "?????";
    endcase
  end
  always @(*) begin
    case(toplevel_execute_ctrl2_up_late0_IntAluPlugin_ALU_BITWISE_CTRL_lane0)
      IntAluPlugin_AluBitwiseCtrlEnum_XOR_1 : toplevel_execute_ctrl2_up_late0_IntAluPlugin_ALU_BITWISE_CTRL_lane0_string = "XOR_1";
      IntAluPlugin_AluBitwiseCtrlEnum_OR_1 : toplevel_execute_ctrl2_up_late0_IntAluPlugin_ALU_BITWISE_CTRL_lane0_string = "OR_1 ";
      IntAluPlugin_AluBitwiseCtrlEnum_AND_1 : toplevel_execute_ctrl2_up_late0_IntAluPlugin_ALU_BITWISE_CTRL_lane0_string = "AND_1";
      IntAluPlugin_AluBitwiseCtrlEnum_ZERO : toplevel_execute_ctrl2_up_late0_IntAluPlugin_ALU_BITWISE_CTRL_lane0_string = "ZERO ";
      default : toplevel_execute_ctrl2_up_late0_IntAluPlugin_ALU_BITWISE_CTRL_lane0_string = "?????";
    endcase
  end
  always @(*) begin
    case(toplevel_execute_ctrl2_up_early0_EnvPlugin_OP_lane0)
      EnvPluginOp_ECALL : toplevel_execute_ctrl2_up_early0_EnvPlugin_OP_lane0_string = "ECALL     ";
      EnvPluginOp_EBREAK : toplevel_execute_ctrl2_up_early0_EnvPlugin_OP_lane0_string = "EBREAK    ";
      EnvPluginOp_PRIV_RET : toplevel_execute_ctrl2_up_early0_EnvPlugin_OP_lane0_string = "PRIV_RET  ";
      EnvPluginOp_FENCE_I : toplevel_execute_ctrl2_up_early0_EnvPlugin_OP_lane0_string = "FENCE_I   ";
      EnvPluginOp_SFENCE_VMA : toplevel_execute_ctrl2_up_early0_EnvPlugin_OP_lane0_string = "SFENCE_VMA";
      EnvPluginOp_WFI : toplevel_execute_ctrl2_up_early0_EnvPlugin_OP_lane0_string = "WFI       ";
      default : toplevel_execute_ctrl2_up_early0_EnvPlugin_OP_lane0_string = "??????????";
    endcase
  end
  always @(*) begin
    case(toplevel_execute_ctrl2_up_BranchPlugin_BRANCH_CTRL_lane0)
      BranchPlugin_BranchCtrlEnum_B : toplevel_execute_ctrl2_up_BranchPlugin_BRANCH_CTRL_lane0_string = "B   ";
      BranchPlugin_BranchCtrlEnum_JAL : toplevel_execute_ctrl2_up_BranchPlugin_BRANCH_CTRL_lane0_string = "JAL ";
      BranchPlugin_BranchCtrlEnum_JALR : toplevel_execute_ctrl2_up_BranchPlugin_BRANCH_CTRL_lane0_string = "JALR";
      default : toplevel_execute_ctrl2_up_BranchPlugin_BRANCH_CTRL_lane0_string = "????";
    endcase
  end
  always @(*) begin
    case(toplevel_execute_ctrl2_up_early0_IntAluPlugin_ALU_BITWISE_CTRL_lane0)
      IntAluPlugin_AluBitwiseCtrlEnum_XOR_1 : toplevel_execute_ctrl2_up_early0_IntAluPlugin_ALU_BITWISE_CTRL_lane0_string = "XOR_1";
      IntAluPlugin_AluBitwiseCtrlEnum_OR_1 : toplevel_execute_ctrl2_up_early0_IntAluPlugin_ALU_BITWISE_CTRL_lane0_string = "OR_1 ";
      IntAluPlugin_AluBitwiseCtrlEnum_AND_1 : toplevel_execute_ctrl2_up_early0_IntAluPlugin_ALU_BITWISE_CTRL_lane0_string = "AND_1";
      IntAluPlugin_AluBitwiseCtrlEnum_ZERO : toplevel_execute_ctrl2_up_early0_IntAluPlugin_ALU_BITWISE_CTRL_lane0_string = "ZERO ";
      default : toplevel_execute_ctrl2_up_early0_IntAluPlugin_ALU_BITWISE_CTRL_lane0_string = "?????";
    endcase
  end
  always @(*) begin
    case(toplevel_execute_ctrl1_down_late1_IntAluPlugin_ALU_BITWISE_CTRL_lane1)
      IntAluPlugin_AluBitwiseCtrlEnum_XOR_1 : toplevel_execute_ctrl1_down_late1_IntAluPlugin_ALU_BITWISE_CTRL_lane1_string = "XOR_1";
      IntAluPlugin_AluBitwiseCtrlEnum_OR_1 : toplevel_execute_ctrl1_down_late1_IntAluPlugin_ALU_BITWISE_CTRL_lane1_string = "OR_1 ";
      IntAluPlugin_AluBitwiseCtrlEnum_AND_1 : toplevel_execute_ctrl1_down_late1_IntAluPlugin_ALU_BITWISE_CTRL_lane1_string = "AND_1";
      IntAluPlugin_AluBitwiseCtrlEnum_ZERO : toplevel_execute_ctrl1_down_late1_IntAluPlugin_ALU_BITWISE_CTRL_lane1_string = "ZERO ";
      default : toplevel_execute_ctrl1_down_late1_IntAluPlugin_ALU_BITWISE_CTRL_lane1_string = "?????";
    endcase
  end
  always @(*) begin
    case(toplevel_execute_ctrl1_down_BranchPlugin_BRANCH_CTRL_lane1)
      BranchPlugin_BranchCtrlEnum_B : toplevel_execute_ctrl1_down_BranchPlugin_BRANCH_CTRL_lane1_string = "B   ";
      BranchPlugin_BranchCtrlEnum_JAL : toplevel_execute_ctrl1_down_BranchPlugin_BRANCH_CTRL_lane1_string = "JAL ";
      BranchPlugin_BranchCtrlEnum_JALR : toplevel_execute_ctrl1_down_BranchPlugin_BRANCH_CTRL_lane1_string = "JALR";
      default : toplevel_execute_ctrl1_down_BranchPlugin_BRANCH_CTRL_lane1_string = "????";
    endcase
  end
  always @(*) begin
    case(toplevel_execute_ctrl1_down_early1_IntAluPlugin_ALU_BITWISE_CTRL_lane1)
      IntAluPlugin_AluBitwiseCtrlEnum_XOR_1 : toplevel_execute_ctrl1_down_early1_IntAluPlugin_ALU_BITWISE_CTRL_lane1_string = "XOR_1";
      IntAluPlugin_AluBitwiseCtrlEnum_OR_1 : toplevel_execute_ctrl1_down_early1_IntAluPlugin_ALU_BITWISE_CTRL_lane1_string = "OR_1 ";
      IntAluPlugin_AluBitwiseCtrlEnum_AND_1 : toplevel_execute_ctrl1_down_early1_IntAluPlugin_ALU_BITWISE_CTRL_lane1_string = "AND_1";
      IntAluPlugin_AluBitwiseCtrlEnum_ZERO : toplevel_execute_ctrl1_down_early1_IntAluPlugin_ALU_BITWISE_CTRL_lane1_string = "ZERO ";
      default : toplevel_execute_ctrl1_down_early1_IntAluPlugin_ALU_BITWISE_CTRL_lane1_string = "?????";
    endcase
  end
  always @(*) begin
    case(toplevel_execute_ctrl1_down_late0_IntAluPlugin_ALU_BITWISE_CTRL_lane0)
      IntAluPlugin_AluBitwiseCtrlEnum_XOR_1 : toplevel_execute_ctrl1_down_late0_IntAluPlugin_ALU_BITWISE_CTRL_lane0_string = "XOR_1";
      IntAluPlugin_AluBitwiseCtrlEnum_OR_1 : toplevel_execute_ctrl1_down_late0_IntAluPlugin_ALU_BITWISE_CTRL_lane0_string = "OR_1 ";
      IntAluPlugin_AluBitwiseCtrlEnum_AND_1 : toplevel_execute_ctrl1_down_late0_IntAluPlugin_ALU_BITWISE_CTRL_lane0_string = "AND_1";
      IntAluPlugin_AluBitwiseCtrlEnum_ZERO : toplevel_execute_ctrl1_down_late0_IntAluPlugin_ALU_BITWISE_CTRL_lane0_string = "ZERO ";
      default : toplevel_execute_ctrl1_down_late0_IntAluPlugin_ALU_BITWISE_CTRL_lane0_string = "?????";
    endcase
  end
  always @(*) begin
    case(toplevel_execute_ctrl1_down_early0_EnvPlugin_OP_lane0)
      EnvPluginOp_ECALL : toplevel_execute_ctrl1_down_early0_EnvPlugin_OP_lane0_string = "ECALL     ";
      EnvPluginOp_EBREAK : toplevel_execute_ctrl1_down_early0_EnvPlugin_OP_lane0_string = "EBREAK    ";
      EnvPluginOp_PRIV_RET : toplevel_execute_ctrl1_down_early0_EnvPlugin_OP_lane0_string = "PRIV_RET  ";
      EnvPluginOp_FENCE_I : toplevel_execute_ctrl1_down_early0_EnvPlugin_OP_lane0_string = "FENCE_I   ";
      EnvPluginOp_SFENCE_VMA : toplevel_execute_ctrl1_down_early0_EnvPlugin_OP_lane0_string = "SFENCE_VMA";
      EnvPluginOp_WFI : toplevel_execute_ctrl1_down_early0_EnvPlugin_OP_lane0_string = "WFI       ";
      default : toplevel_execute_ctrl1_down_early0_EnvPlugin_OP_lane0_string = "??????????";
    endcase
  end
  always @(*) begin
    case(toplevel_execute_ctrl1_down_BranchPlugin_BRANCH_CTRL_lane0)
      BranchPlugin_BranchCtrlEnum_B : toplevel_execute_ctrl1_down_BranchPlugin_BRANCH_CTRL_lane0_string = "B   ";
      BranchPlugin_BranchCtrlEnum_JAL : toplevel_execute_ctrl1_down_BranchPlugin_BRANCH_CTRL_lane0_string = "JAL ";
      BranchPlugin_BranchCtrlEnum_JALR : toplevel_execute_ctrl1_down_BranchPlugin_BRANCH_CTRL_lane0_string = "JALR";
      default : toplevel_execute_ctrl1_down_BranchPlugin_BRANCH_CTRL_lane0_string = "????";
    endcase
  end
  always @(*) begin
    case(toplevel_execute_ctrl1_down_early0_IntAluPlugin_ALU_BITWISE_CTRL_lane0)
      IntAluPlugin_AluBitwiseCtrlEnum_XOR_1 : toplevel_execute_ctrl1_down_early0_IntAluPlugin_ALU_BITWISE_CTRL_lane0_string = "XOR_1";
      IntAluPlugin_AluBitwiseCtrlEnum_OR_1 : toplevel_execute_ctrl1_down_early0_IntAluPlugin_ALU_BITWISE_CTRL_lane0_string = "OR_1 ";
      IntAluPlugin_AluBitwiseCtrlEnum_AND_1 : toplevel_execute_ctrl1_down_early0_IntAluPlugin_ALU_BITWISE_CTRL_lane0_string = "AND_1";
      IntAluPlugin_AluBitwiseCtrlEnum_ZERO : toplevel_execute_ctrl1_down_early0_IntAluPlugin_ALU_BITWISE_CTRL_lane0_string = "ZERO ";
      default : toplevel_execute_ctrl1_down_early0_IntAluPlugin_ALU_BITWISE_CTRL_lane0_string = "?????";
    endcase
  end
  always @(*) begin
    case(toplevel_execute_ctrl4_down_BranchPlugin_BRANCH_CTRL_lane1)
      BranchPlugin_BranchCtrlEnum_B : toplevel_execute_ctrl4_down_BranchPlugin_BRANCH_CTRL_lane1_string = "B   ";
      BranchPlugin_BranchCtrlEnum_JAL : toplevel_execute_ctrl4_down_BranchPlugin_BRANCH_CTRL_lane1_string = "JAL ";
      BranchPlugin_BranchCtrlEnum_JALR : toplevel_execute_ctrl4_down_BranchPlugin_BRANCH_CTRL_lane1_string = "JALR";
      default : toplevel_execute_ctrl4_down_BranchPlugin_BRANCH_CTRL_lane1_string = "????";
    endcase
  end
  always @(*) begin
    case(toplevel_execute_ctrl4_down_BranchPlugin_BRANCH_CTRL_lane0)
      BranchPlugin_BranchCtrlEnum_B : toplevel_execute_ctrl4_down_BranchPlugin_BRANCH_CTRL_lane0_string = "B   ";
      BranchPlugin_BranchCtrlEnum_JAL : toplevel_execute_ctrl4_down_BranchPlugin_BRANCH_CTRL_lane0_string = "JAL ";
      BranchPlugin_BranchCtrlEnum_JALR : toplevel_execute_ctrl4_down_BranchPlugin_BRANCH_CTRL_lane0_string = "JALR";
      default : toplevel_execute_ctrl4_down_BranchPlugin_BRANCH_CTRL_lane0_string = "????";
    endcase
  end
  always @(*) begin
    case(toplevel_execute_ctrl3_down_BranchPlugin_BRANCH_CTRL_lane1)
      BranchPlugin_BranchCtrlEnum_B : toplevel_execute_ctrl3_down_BranchPlugin_BRANCH_CTRL_lane1_string = "B   ";
      BranchPlugin_BranchCtrlEnum_JAL : toplevel_execute_ctrl3_down_BranchPlugin_BRANCH_CTRL_lane1_string = "JAL ";
      BranchPlugin_BranchCtrlEnum_JALR : toplevel_execute_ctrl3_down_BranchPlugin_BRANCH_CTRL_lane1_string = "JALR";
      default : toplevel_execute_ctrl3_down_BranchPlugin_BRANCH_CTRL_lane1_string = "????";
    endcase
  end
  always @(*) begin
    case(toplevel_execute_ctrl2_down_early0_EnvPlugin_OP_lane0)
      EnvPluginOp_ECALL : toplevel_execute_ctrl2_down_early0_EnvPlugin_OP_lane0_string = "ECALL     ";
      EnvPluginOp_EBREAK : toplevel_execute_ctrl2_down_early0_EnvPlugin_OP_lane0_string = "EBREAK    ";
      EnvPluginOp_PRIV_RET : toplevel_execute_ctrl2_down_early0_EnvPlugin_OP_lane0_string = "PRIV_RET  ";
      EnvPluginOp_FENCE_I : toplevel_execute_ctrl2_down_early0_EnvPlugin_OP_lane0_string = "FENCE_I   ";
      EnvPluginOp_SFENCE_VMA : toplevel_execute_ctrl2_down_early0_EnvPlugin_OP_lane0_string = "SFENCE_VMA";
      EnvPluginOp_WFI : toplevel_execute_ctrl2_down_early0_EnvPlugin_OP_lane0_string = "WFI       ";
      default : toplevel_execute_ctrl2_down_early0_EnvPlugin_OP_lane0_string = "??????????";
    endcase
  end
  always @(*) begin
    case(toplevel_execute_ctrl3_down_BranchPlugin_BRANCH_CTRL_lane0)
      BranchPlugin_BranchCtrlEnum_B : toplevel_execute_ctrl3_down_BranchPlugin_BRANCH_CTRL_lane0_string = "B   ";
      BranchPlugin_BranchCtrlEnum_JAL : toplevel_execute_ctrl3_down_BranchPlugin_BRANCH_CTRL_lane0_string = "JAL ";
      BranchPlugin_BranchCtrlEnum_JALR : toplevel_execute_ctrl3_down_BranchPlugin_BRANCH_CTRL_lane0_string = "JALR";
      default : toplevel_execute_ctrl3_down_BranchPlugin_BRANCH_CTRL_lane0_string = "????";
    endcase
  end
  always @(*) begin
    case(toplevel_execute_ctrl2_down_BranchPlugin_BRANCH_CTRL_lane1)
      BranchPlugin_BranchCtrlEnum_B : toplevel_execute_ctrl2_down_BranchPlugin_BRANCH_CTRL_lane1_string = "B   ";
      BranchPlugin_BranchCtrlEnum_JAL : toplevel_execute_ctrl2_down_BranchPlugin_BRANCH_CTRL_lane1_string = "JAL ";
      BranchPlugin_BranchCtrlEnum_JALR : toplevel_execute_ctrl2_down_BranchPlugin_BRANCH_CTRL_lane1_string = "JALR";
      default : toplevel_execute_ctrl2_down_BranchPlugin_BRANCH_CTRL_lane1_string = "????";
    endcase
  end
  always @(*) begin
    case(toplevel_execute_ctrl2_down_BranchPlugin_BRANCH_CTRL_lane0)
      BranchPlugin_BranchCtrlEnum_B : toplevel_execute_ctrl2_down_BranchPlugin_BRANCH_CTRL_lane0_string = "B   ";
      BranchPlugin_BranchCtrlEnum_JAL : toplevel_execute_ctrl2_down_BranchPlugin_BRANCH_CTRL_lane0_string = "JAL ";
      BranchPlugin_BranchCtrlEnum_JALR : toplevel_execute_ctrl2_down_BranchPlugin_BRANCH_CTRL_lane0_string = "JALR";
      default : toplevel_execute_ctrl2_down_BranchPlugin_BRANCH_CTRL_lane0_string = "????";
    endcase
  end
  always @(*) begin
    case(toplevel_execute_ctrl4_down_late1_IntAluPlugin_ALU_BITWISE_CTRL_lane1)
      IntAluPlugin_AluBitwiseCtrlEnum_XOR_1 : toplevel_execute_ctrl4_down_late1_IntAluPlugin_ALU_BITWISE_CTRL_lane1_string = "XOR_1";
      IntAluPlugin_AluBitwiseCtrlEnum_OR_1 : toplevel_execute_ctrl4_down_late1_IntAluPlugin_ALU_BITWISE_CTRL_lane1_string = "OR_1 ";
      IntAluPlugin_AluBitwiseCtrlEnum_AND_1 : toplevel_execute_ctrl4_down_late1_IntAluPlugin_ALU_BITWISE_CTRL_lane1_string = "AND_1";
      IntAluPlugin_AluBitwiseCtrlEnum_ZERO : toplevel_execute_ctrl4_down_late1_IntAluPlugin_ALU_BITWISE_CTRL_lane1_string = "ZERO ";
      default : toplevel_execute_ctrl4_down_late1_IntAluPlugin_ALU_BITWISE_CTRL_lane1_string = "?????";
    endcase
  end
  always @(*) begin
    case(toplevel_execute_ctrl2_down_early1_IntAluPlugin_ALU_BITWISE_CTRL_lane1)
      IntAluPlugin_AluBitwiseCtrlEnum_XOR_1 : toplevel_execute_ctrl2_down_early1_IntAluPlugin_ALU_BITWISE_CTRL_lane1_string = "XOR_1";
      IntAluPlugin_AluBitwiseCtrlEnum_OR_1 : toplevel_execute_ctrl2_down_early1_IntAluPlugin_ALU_BITWISE_CTRL_lane1_string = "OR_1 ";
      IntAluPlugin_AluBitwiseCtrlEnum_AND_1 : toplevel_execute_ctrl2_down_early1_IntAluPlugin_ALU_BITWISE_CTRL_lane1_string = "AND_1";
      IntAluPlugin_AluBitwiseCtrlEnum_ZERO : toplevel_execute_ctrl2_down_early1_IntAluPlugin_ALU_BITWISE_CTRL_lane1_string = "ZERO ";
      default : toplevel_execute_ctrl2_down_early1_IntAluPlugin_ALU_BITWISE_CTRL_lane1_string = "?????";
    endcase
  end
  always @(*) begin
    case(toplevel_execute_ctrl4_down_late0_IntAluPlugin_ALU_BITWISE_CTRL_lane0)
      IntAluPlugin_AluBitwiseCtrlEnum_XOR_1 : toplevel_execute_ctrl4_down_late0_IntAluPlugin_ALU_BITWISE_CTRL_lane0_string = "XOR_1";
      IntAluPlugin_AluBitwiseCtrlEnum_OR_1 : toplevel_execute_ctrl4_down_late0_IntAluPlugin_ALU_BITWISE_CTRL_lane0_string = "OR_1 ";
      IntAluPlugin_AluBitwiseCtrlEnum_AND_1 : toplevel_execute_ctrl4_down_late0_IntAluPlugin_ALU_BITWISE_CTRL_lane0_string = "AND_1";
      IntAluPlugin_AluBitwiseCtrlEnum_ZERO : toplevel_execute_ctrl4_down_late0_IntAluPlugin_ALU_BITWISE_CTRL_lane0_string = "ZERO ";
      default : toplevel_execute_ctrl4_down_late0_IntAluPlugin_ALU_BITWISE_CTRL_lane0_string = "?????";
    endcase
  end
  always @(*) begin
    case(toplevel_execute_ctrl2_down_early0_IntAluPlugin_ALU_BITWISE_CTRL_lane0)
      IntAluPlugin_AluBitwiseCtrlEnum_XOR_1 : toplevel_execute_ctrl2_down_early0_IntAluPlugin_ALU_BITWISE_CTRL_lane0_string = "XOR_1";
      IntAluPlugin_AluBitwiseCtrlEnum_OR_1 : toplevel_execute_ctrl2_down_early0_IntAluPlugin_ALU_BITWISE_CTRL_lane0_string = "OR_1 ";
      IntAluPlugin_AluBitwiseCtrlEnum_AND_1 : toplevel_execute_ctrl2_down_early0_IntAluPlugin_ALU_BITWISE_CTRL_lane0_string = "AND_1";
      IntAluPlugin_AluBitwiseCtrlEnum_ZERO : toplevel_execute_ctrl2_down_early0_IntAluPlugin_ALU_BITWISE_CTRL_lane0_string = "ZERO ";
      default : toplevel_execute_ctrl2_down_early0_IntAluPlugin_ALU_BITWISE_CTRL_lane0_string = "?????";
    endcase
  end
  always @(*) begin
    case(FetchL1TileLinkPlugin_logic_down_a_payload_opcode)
      A_PUT_FULL_DATA : FetchL1TileLinkPlugin_logic_down_a_payload_opcode_string = "PUT_FULL_DATA   ";
      A_PUT_PARTIAL_DATA : FetchL1TileLinkPlugin_logic_down_a_payload_opcode_string = "PUT_PARTIAL_DATA";
      A_GET : FetchL1TileLinkPlugin_logic_down_a_payload_opcode_string = "GET             ";
      A_ACQUIRE_BLOCK : FetchL1TileLinkPlugin_logic_down_a_payload_opcode_string = "ACQUIRE_BLOCK   ";
      A_ACQUIRE_PERM : FetchL1TileLinkPlugin_logic_down_a_payload_opcode_string = "ACQUIRE_PERM    ";
      default : FetchL1TileLinkPlugin_logic_down_a_payload_opcode_string = "????????????????";
    endcase
  end
  always @(*) begin
    case(FetchL1TileLinkPlugin_logic_down_d_payload_opcode)
      D_ACCESS_ACK : FetchL1TileLinkPlugin_logic_down_d_payload_opcode_string = "ACCESS_ACK     ";
      D_ACCESS_ACK_DATA : FetchL1TileLinkPlugin_logic_down_d_payload_opcode_string = "ACCESS_ACK_DATA";
      D_GRANT : FetchL1TileLinkPlugin_logic_down_d_payload_opcode_string = "GRANT          ";
      D_GRANT_DATA : FetchL1TileLinkPlugin_logic_down_d_payload_opcode_string = "GRANT_DATA     ";
      D_RELEASE_ACK : FetchL1TileLinkPlugin_logic_down_d_payload_opcode_string = "RELEASE_ACK    ";
      default : FetchL1TileLinkPlugin_logic_down_d_payload_opcode_string = "???????????????";
    endcase
  end
  always @(*) begin
    case(LsuPlugin_logic_onAddress0_ls_port_payload_op)
      LsuL1CmdOpcode_LSU : LsuPlugin_logic_onAddress0_ls_port_payload_op_string = "LSU         ";
      LsuL1CmdOpcode_ACCESS_1 : LsuPlugin_logic_onAddress0_ls_port_payload_op_string = "ACCESS_1    ";
      LsuL1CmdOpcode_STORE_BUFFER : LsuPlugin_logic_onAddress0_ls_port_payload_op_string = "STORE_BUFFER";
      LsuL1CmdOpcode_FLUSH : LsuPlugin_logic_onAddress0_ls_port_payload_op_string = "FLUSH       ";
      LsuL1CmdOpcode_PREFETCH : LsuPlugin_logic_onAddress0_ls_port_payload_op_string = "PREFETCH    ";
      default : LsuPlugin_logic_onAddress0_ls_port_payload_op_string = "????????????";
    endcase
  end
  always @(*) begin
    case(LsuPlugin_logic_onAddress0_access_port_payload_op)
      LsuL1CmdOpcode_LSU : LsuPlugin_logic_onAddress0_access_port_payload_op_string = "LSU         ";
      LsuL1CmdOpcode_ACCESS_1 : LsuPlugin_logic_onAddress0_access_port_payload_op_string = "ACCESS_1    ";
      LsuL1CmdOpcode_STORE_BUFFER : LsuPlugin_logic_onAddress0_access_port_payload_op_string = "STORE_BUFFER";
      LsuL1CmdOpcode_FLUSH : LsuPlugin_logic_onAddress0_access_port_payload_op_string = "FLUSH       ";
      LsuL1CmdOpcode_PREFETCH : LsuPlugin_logic_onAddress0_access_port_payload_op_string = "PREFETCH    ";
      default : LsuPlugin_logic_onAddress0_access_port_payload_op_string = "????????????";
    endcase
  end
  always @(*) begin
    case(LsuPlugin_logic_onAddress0_flush_port_payload_op)
      LsuL1CmdOpcode_LSU : LsuPlugin_logic_onAddress0_flush_port_payload_op_string = "LSU         ";
      LsuL1CmdOpcode_ACCESS_1 : LsuPlugin_logic_onAddress0_flush_port_payload_op_string = "ACCESS_1    ";
      LsuL1CmdOpcode_STORE_BUFFER : LsuPlugin_logic_onAddress0_flush_port_payload_op_string = "STORE_BUFFER";
      LsuL1CmdOpcode_FLUSH : LsuPlugin_logic_onAddress0_flush_port_payload_op_string = "FLUSH       ";
      LsuL1CmdOpcode_PREFETCH : LsuPlugin_logic_onAddress0_flush_port_payload_op_string = "PREFETCH    ";
      default : LsuPlugin_logic_onAddress0_flush_port_payload_op_string = "????????????";
    endcase
  end
  always @(*) begin
    case(LsuL1TileLinkPlugin_logic_down_a_payload_opcode)
      A_PUT_FULL_DATA : LsuL1TileLinkPlugin_logic_down_a_payload_opcode_string = "PUT_FULL_DATA   ";
      A_PUT_PARTIAL_DATA : LsuL1TileLinkPlugin_logic_down_a_payload_opcode_string = "PUT_PARTIAL_DATA";
      A_GET : LsuL1TileLinkPlugin_logic_down_a_payload_opcode_string = "GET             ";
      A_ACQUIRE_BLOCK : LsuL1TileLinkPlugin_logic_down_a_payload_opcode_string = "ACQUIRE_BLOCK   ";
      A_ACQUIRE_PERM : LsuL1TileLinkPlugin_logic_down_a_payload_opcode_string = "ACQUIRE_PERM    ";
      default : LsuL1TileLinkPlugin_logic_down_a_payload_opcode_string = "????????????????";
    endcase
  end
  always @(*) begin
    case(LsuL1TileLinkPlugin_logic_down_d_payload_opcode)
      D_ACCESS_ACK : LsuL1TileLinkPlugin_logic_down_d_payload_opcode_string = "ACCESS_ACK     ";
      D_ACCESS_ACK_DATA : LsuL1TileLinkPlugin_logic_down_d_payload_opcode_string = "ACCESS_ACK_DATA";
      D_GRANT : LsuL1TileLinkPlugin_logic_down_d_payload_opcode_string = "GRANT          ";
      D_GRANT_DATA : LsuL1TileLinkPlugin_logic_down_d_payload_opcode_string = "GRANT_DATA     ";
      D_RELEASE_ACK : LsuL1TileLinkPlugin_logic_down_d_payload_opcode_string = "RELEASE_ACK    ";
      default : LsuL1TileLinkPlugin_logic_down_d_payload_opcode_string = "???????????????";
    endcase
  end
  always @(*) begin
    case(LsuTileLinkPlugin_logic_bridge_down_a_payload_opcode)
      A_PUT_FULL_DATA : LsuTileLinkPlugin_logic_bridge_down_a_payload_opcode_string = "PUT_FULL_DATA   ";
      A_PUT_PARTIAL_DATA : LsuTileLinkPlugin_logic_bridge_down_a_payload_opcode_string = "PUT_PARTIAL_DATA";
      A_GET : LsuTileLinkPlugin_logic_bridge_down_a_payload_opcode_string = "GET             ";
      A_ACQUIRE_BLOCK : LsuTileLinkPlugin_logic_bridge_down_a_payload_opcode_string = "ACQUIRE_BLOCK   ";
      A_ACQUIRE_PERM : LsuTileLinkPlugin_logic_bridge_down_a_payload_opcode_string = "ACQUIRE_PERM    ";
      default : LsuTileLinkPlugin_logic_bridge_down_a_payload_opcode_string = "????????????????";
    endcase
  end
  always @(*) begin
    case(LsuTileLinkPlugin_logic_bridge_down_d_payload_opcode)
      D_ACCESS_ACK : LsuTileLinkPlugin_logic_bridge_down_d_payload_opcode_string = "ACCESS_ACK     ";
      D_ACCESS_ACK_DATA : LsuTileLinkPlugin_logic_bridge_down_d_payload_opcode_string = "ACCESS_ACK_DATA";
      D_GRANT : LsuTileLinkPlugin_logic_bridge_down_d_payload_opcode_string = "GRANT          ";
      D_GRANT_DATA : LsuTileLinkPlugin_logic_bridge_down_d_payload_opcode_string = "GRANT_DATA     ";
      D_RELEASE_ACK : LsuTileLinkPlugin_logic_bridge_down_d_payload_opcode_string = "RELEASE_ACK    ";
      default : LsuTileLinkPlugin_logic_bridge_down_d_payload_opcode_string = "???????????????";
    endcase
  end
  always @(*) begin
    case(_zz_LsuTileLinkPlugin_logic_bridge_down_a_payload_opcode)
      A_PUT_FULL_DATA : _zz_LsuTileLinkPlugin_logic_bridge_down_a_payload_opcode_string = "PUT_FULL_DATA   ";
      A_PUT_PARTIAL_DATA : _zz_LsuTileLinkPlugin_logic_bridge_down_a_payload_opcode_string = "PUT_PARTIAL_DATA";
      A_GET : _zz_LsuTileLinkPlugin_logic_bridge_down_a_payload_opcode_string = "GET             ";
      A_ACQUIRE_BLOCK : _zz_LsuTileLinkPlugin_logic_bridge_down_a_payload_opcode_string = "ACQUIRE_BLOCK   ";
      A_ACQUIRE_PERM : _zz_LsuTileLinkPlugin_logic_bridge_down_a_payload_opcode_string = "ACQUIRE_PERM    ";
      default : _zz_LsuTileLinkPlugin_logic_bridge_down_a_payload_opcode_string = "????????????????";
    endcase
  end
  always @(*) begin
    case(_zz_toplevel_execute_ctrl1_down_early0_IntAluPlugin_ALU_BITWISE_CTRL_lane0)
      IntAluPlugin_AluBitwiseCtrlEnum_XOR_1 : _zz_toplevel_execute_ctrl1_down_early0_IntAluPlugin_ALU_BITWISE_CTRL_lane0_string = "XOR_1";
      IntAluPlugin_AluBitwiseCtrlEnum_OR_1 : _zz_toplevel_execute_ctrl1_down_early0_IntAluPlugin_ALU_BITWISE_CTRL_lane0_string = "OR_1 ";
      IntAluPlugin_AluBitwiseCtrlEnum_AND_1 : _zz_toplevel_execute_ctrl1_down_early0_IntAluPlugin_ALU_BITWISE_CTRL_lane0_string = "AND_1";
      IntAluPlugin_AluBitwiseCtrlEnum_ZERO : _zz_toplevel_execute_ctrl1_down_early0_IntAluPlugin_ALU_BITWISE_CTRL_lane0_string = "ZERO ";
      default : _zz_toplevel_execute_ctrl1_down_early0_IntAluPlugin_ALU_BITWISE_CTRL_lane0_string = "?????";
    endcase
  end
  always @(*) begin
    case(_zz_toplevel_execute_ctrl1_down_early0_IntAluPlugin_ALU_BITWISE_CTRL_lane0_1)
      IntAluPlugin_AluBitwiseCtrlEnum_XOR_1 : _zz_toplevel_execute_ctrl1_down_early0_IntAluPlugin_ALU_BITWISE_CTRL_lane0_1_string = "XOR_1";
      IntAluPlugin_AluBitwiseCtrlEnum_OR_1 : _zz_toplevel_execute_ctrl1_down_early0_IntAluPlugin_ALU_BITWISE_CTRL_lane0_1_string = "OR_1 ";
      IntAluPlugin_AluBitwiseCtrlEnum_AND_1 : _zz_toplevel_execute_ctrl1_down_early0_IntAluPlugin_ALU_BITWISE_CTRL_lane0_1_string = "AND_1";
      IntAluPlugin_AluBitwiseCtrlEnum_ZERO : _zz_toplevel_execute_ctrl1_down_early0_IntAluPlugin_ALU_BITWISE_CTRL_lane0_1_string = "ZERO ";
      default : _zz_toplevel_execute_ctrl1_down_early0_IntAluPlugin_ALU_BITWISE_CTRL_lane0_1_string = "?????";
    endcase
  end
  always @(*) begin
    case(_zz_toplevel_execute_ctrl1_down_early0_IntAluPlugin_ALU_BITWISE_CTRL_lane0_2)
      IntAluPlugin_AluBitwiseCtrlEnum_XOR_1 : _zz_toplevel_execute_ctrl1_down_early0_IntAluPlugin_ALU_BITWISE_CTRL_lane0_2_string = "XOR_1";
      IntAluPlugin_AluBitwiseCtrlEnum_OR_1 : _zz_toplevel_execute_ctrl1_down_early0_IntAluPlugin_ALU_BITWISE_CTRL_lane0_2_string = "OR_1 ";
      IntAluPlugin_AluBitwiseCtrlEnum_AND_1 : _zz_toplevel_execute_ctrl1_down_early0_IntAluPlugin_ALU_BITWISE_CTRL_lane0_2_string = "AND_1";
      IntAluPlugin_AluBitwiseCtrlEnum_ZERO : _zz_toplevel_execute_ctrl1_down_early0_IntAluPlugin_ALU_BITWISE_CTRL_lane0_2_string = "ZERO ";
      default : _zz_toplevel_execute_ctrl1_down_early0_IntAluPlugin_ALU_BITWISE_CTRL_lane0_2_string = "?????";
    endcase
  end
  always @(*) begin
    case(_zz_toplevel_execute_ctrl1_down_BranchPlugin_BRANCH_CTRL_lane0)
      BranchPlugin_BranchCtrlEnum_B : _zz_toplevel_execute_ctrl1_down_BranchPlugin_BRANCH_CTRL_lane0_string = "B   ";
      BranchPlugin_BranchCtrlEnum_JAL : _zz_toplevel_execute_ctrl1_down_BranchPlugin_BRANCH_CTRL_lane0_string = "JAL ";
      BranchPlugin_BranchCtrlEnum_JALR : _zz_toplevel_execute_ctrl1_down_BranchPlugin_BRANCH_CTRL_lane0_string = "JALR";
      default : _zz_toplevel_execute_ctrl1_down_BranchPlugin_BRANCH_CTRL_lane0_string = "????";
    endcase
  end
  always @(*) begin
    case(_zz_toplevel_execute_ctrl1_down_BranchPlugin_BRANCH_CTRL_lane0_1)
      BranchPlugin_BranchCtrlEnum_B : _zz_toplevel_execute_ctrl1_down_BranchPlugin_BRANCH_CTRL_lane0_1_string = "B   ";
      BranchPlugin_BranchCtrlEnum_JAL : _zz_toplevel_execute_ctrl1_down_BranchPlugin_BRANCH_CTRL_lane0_1_string = "JAL ";
      BranchPlugin_BranchCtrlEnum_JALR : _zz_toplevel_execute_ctrl1_down_BranchPlugin_BRANCH_CTRL_lane0_1_string = "JALR";
      default : _zz_toplevel_execute_ctrl1_down_BranchPlugin_BRANCH_CTRL_lane0_1_string = "????";
    endcase
  end
  always @(*) begin
    case(_zz_toplevel_execute_ctrl1_down_BranchPlugin_BRANCH_CTRL_lane0_2)
      BranchPlugin_BranchCtrlEnum_B : _zz_toplevel_execute_ctrl1_down_BranchPlugin_BRANCH_CTRL_lane0_2_string = "B   ";
      BranchPlugin_BranchCtrlEnum_JAL : _zz_toplevel_execute_ctrl1_down_BranchPlugin_BRANCH_CTRL_lane0_2_string = "JAL ";
      BranchPlugin_BranchCtrlEnum_JALR : _zz_toplevel_execute_ctrl1_down_BranchPlugin_BRANCH_CTRL_lane0_2_string = "JALR";
      default : _zz_toplevel_execute_ctrl1_down_BranchPlugin_BRANCH_CTRL_lane0_2_string = "????";
    endcase
  end
  always @(*) begin
    case(_zz_toplevel_execute_ctrl1_down_early0_EnvPlugin_OP_lane0_1)
      EnvPluginOp_ECALL : _zz_toplevel_execute_ctrl1_down_early0_EnvPlugin_OP_lane0_1_string = "ECALL     ";
      EnvPluginOp_EBREAK : _zz_toplevel_execute_ctrl1_down_early0_EnvPlugin_OP_lane0_1_string = "EBREAK    ";
      EnvPluginOp_PRIV_RET : _zz_toplevel_execute_ctrl1_down_early0_EnvPlugin_OP_lane0_1_string = "PRIV_RET  ";
      EnvPluginOp_FENCE_I : _zz_toplevel_execute_ctrl1_down_early0_EnvPlugin_OP_lane0_1_string = "FENCE_I   ";
      EnvPluginOp_SFENCE_VMA : _zz_toplevel_execute_ctrl1_down_early0_EnvPlugin_OP_lane0_1_string = "SFENCE_VMA";
      EnvPluginOp_WFI : _zz_toplevel_execute_ctrl1_down_early0_EnvPlugin_OP_lane0_1_string = "WFI       ";
      default : _zz_toplevel_execute_ctrl1_down_early0_EnvPlugin_OP_lane0_1_string = "??????????";
    endcase
  end
  always @(*) begin
    case(_zz_toplevel_execute_ctrl1_down_early0_EnvPlugin_OP_lane0_2)
      EnvPluginOp_ECALL : _zz_toplevel_execute_ctrl1_down_early0_EnvPlugin_OP_lane0_2_string = "ECALL     ";
      EnvPluginOp_EBREAK : _zz_toplevel_execute_ctrl1_down_early0_EnvPlugin_OP_lane0_2_string = "EBREAK    ";
      EnvPluginOp_PRIV_RET : _zz_toplevel_execute_ctrl1_down_early0_EnvPlugin_OP_lane0_2_string = "PRIV_RET  ";
      EnvPluginOp_FENCE_I : _zz_toplevel_execute_ctrl1_down_early0_EnvPlugin_OP_lane0_2_string = "FENCE_I   ";
      EnvPluginOp_SFENCE_VMA : _zz_toplevel_execute_ctrl1_down_early0_EnvPlugin_OP_lane0_2_string = "SFENCE_VMA";
      EnvPluginOp_WFI : _zz_toplevel_execute_ctrl1_down_early0_EnvPlugin_OP_lane0_2_string = "WFI       ";
      default : _zz_toplevel_execute_ctrl1_down_early0_EnvPlugin_OP_lane0_2_string = "??????????";
    endcase
  end
  always @(*) begin
    case(_zz_toplevel_execute_ctrl1_down_early0_EnvPlugin_OP_lane0_3)
      EnvPluginOp_ECALL : _zz_toplevel_execute_ctrl1_down_early0_EnvPlugin_OP_lane0_3_string = "ECALL     ";
      EnvPluginOp_EBREAK : _zz_toplevel_execute_ctrl1_down_early0_EnvPlugin_OP_lane0_3_string = "EBREAK    ";
      EnvPluginOp_PRIV_RET : _zz_toplevel_execute_ctrl1_down_early0_EnvPlugin_OP_lane0_3_string = "PRIV_RET  ";
      EnvPluginOp_FENCE_I : _zz_toplevel_execute_ctrl1_down_early0_EnvPlugin_OP_lane0_3_string = "FENCE_I   ";
      EnvPluginOp_SFENCE_VMA : _zz_toplevel_execute_ctrl1_down_early0_EnvPlugin_OP_lane0_3_string = "SFENCE_VMA";
      EnvPluginOp_WFI : _zz_toplevel_execute_ctrl1_down_early0_EnvPlugin_OP_lane0_3_string = "WFI       ";
      default : _zz_toplevel_execute_ctrl1_down_early0_EnvPlugin_OP_lane0_3_string = "??????????";
    endcase
  end
  always @(*) begin
    case(_zz_toplevel_execute_ctrl1_down_late0_IntAluPlugin_ALU_BITWISE_CTRL_lane0_1)
      IntAluPlugin_AluBitwiseCtrlEnum_XOR_1 : _zz_toplevel_execute_ctrl1_down_late0_IntAluPlugin_ALU_BITWISE_CTRL_lane0_1_string = "XOR_1";
      IntAluPlugin_AluBitwiseCtrlEnum_OR_1 : _zz_toplevel_execute_ctrl1_down_late0_IntAluPlugin_ALU_BITWISE_CTRL_lane0_1_string = "OR_1 ";
      IntAluPlugin_AluBitwiseCtrlEnum_AND_1 : _zz_toplevel_execute_ctrl1_down_late0_IntAluPlugin_ALU_BITWISE_CTRL_lane0_1_string = "AND_1";
      IntAluPlugin_AluBitwiseCtrlEnum_ZERO : _zz_toplevel_execute_ctrl1_down_late0_IntAluPlugin_ALU_BITWISE_CTRL_lane0_1_string = "ZERO ";
      default : _zz_toplevel_execute_ctrl1_down_late0_IntAluPlugin_ALU_BITWISE_CTRL_lane0_1_string = "?????";
    endcase
  end
  always @(*) begin
    case(_zz_toplevel_execute_ctrl1_down_late0_IntAluPlugin_ALU_BITWISE_CTRL_lane0_2)
      IntAluPlugin_AluBitwiseCtrlEnum_XOR_1 : _zz_toplevel_execute_ctrl1_down_late0_IntAluPlugin_ALU_BITWISE_CTRL_lane0_2_string = "XOR_1";
      IntAluPlugin_AluBitwiseCtrlEnum_OR_1 : _zz_toplevel_execute_ctrl1_down_late0_IntAluPlugin_ALU_BITWISE_CTRL_lane0_2_string = "OR_1 ";
      IntAluPlugin_AluBitwiseCtrlEnum_AND_1 : _zz_toplevel_execute_ctrl1_down_late0_IntAluPlugin_ALU_BITWISE_CTRL_lane0_2_string = "AND_1";
      IntAluPlugin_AluBitwiseCtrlEnum_ZERO : _zz_toplevel_execute_ctrl1_down_late0_IntAluPlugin_ALU_BITWISE_CTRL_lane0_2_string = "ZERO ";
      default : _zz_toplevel_execute_ctrl1_down_late0_IntAluPlugin_ALU_BITWISE_CTRL_lane0_2_string = "?????";
    endcase
  end
  always @(*) begin
    case(_zz_toplevel_execute_ctrl1_down_late0_IntAluPlugin_ALU_BITWISE_CTRL_lane0_3)
      IntAluPlugin_AluBitwiseCtrlEnum_XOR_1 : _zz_toplevel_execute_ctrl1_down_late0_IntAluPlugin_ALU_BITWISE_CTRL_lane0_3_string = "XOR_1";
      IntAluPlugin_AluBitwiseCtrlEnum_OR_1 : _zz_toplevel_execute_ctrl1_down_late0_IntAluPlugin_ALU_BITWISE_CTRL_lane0_3_string = "OR_1 ";
      IntAluPlugin_AluBitwiseCtrlEnum_AND_1 : _zz_toplevel_execute_ctrl1_down_late0_IntAluPlugin_ALU_BITWISE_CTRL_lane0_3_string = "AND_1";
      IntAluPlugin_AluBitwiseCtrlEnum_ZERO : _zz_toplevel_execute_ctrl1_down_late0_IntAluPlugin_ALU_BITWISE_CTRL_lane0_3_string = "ZERO ";
      default : _zz_toplevel_execute_ctrl1_down_late0_IntAluPlugin_ALU_BITWISE_CTRL_lane0_3_string = "?????";
    endcase
  end
  always @(*) begin
    case(_zz_toplevel_execute_ctrl1_down_early1_IntAluPlugin_ALU_BITWISE_CTRL_lane1)
      IntAluPlugin_AluBitwiseCtrlEnum_XOR_1 : _zz_toplevel_execute_ctrl1_down_early1_IntAluPlugin_ALU_BITWISE_CTRL_lane1_string = "XOR_1";
      IntAluPlugin_AluBitwiseCtrlEnum_OR_1 : _zz_toplevel_execute_ctrl1_down_early1_IntAluPlugin_ALU_BITWISE_CTRL_lane1_string = "OR_1 ";
      IntAluPlugin_AluBitwiseCtrlEnum_AND_1 : _zz_toplevel_execute_ctrl1_down_early1_IntAluPlugin_ALU_BITWISE_CTRL_lane1_string = "AND_1";
      IntAluPlugin_AluBitwiseCtrlEnum_ZERO : _zz_toplevel_execute_ctrl1_down_early1_IntAluPlugin_ALU_BITWISE_CTRL_lane1_string = "ZERO ";
      default : _zz_toplevel_execute_ctrl1_down_early1_IntAluPlugin_ALU_BITWISE_CTRL_lane1_string = "?????";
    endcase
  end
  always @(*) begin
    case(_zz_toplevel_execute_ctrl1_down_early1_IntAluPlugin_ALU_BITWISE_CTRL_lane1_1)
      IntAluPlugin_AluBitwiseCtrlEnum_XOR_1 : _zz_toplevel_execute_ctrl1_down_early1_IntAluPlugin_ALU_BITWISE_CTRL_lane1_1_string = "XOR_1";
      IntAluPlugin_AluBitwiseCtrlEnum_OR_1 : _zz_toplevel_execute_ctrl1_down_early1_IntAluPlugin_ALU_BITWISE_CTRL_lane1_1_string = "OR_1 ";
      IntAluPlugin_AluBitwiseCtrlEnum_AND_1 : _zz_toplevel_execute_ctrl1_down_early1_IntAluPlugin_ALU_BITWISE_CTRL_lane1_1_string = "AND_1";
      IntAluPlugin_AluBitwiseCtrlEnum_ZERO : _zz_toplevel_execute_ctrl1_down_early1_IntAluPlugin_ALU_BITWISE_CTRL_lane1_1_string = "ZERO ";
      default : _zz_toplevel_execute_ctrl1_down_early1_IntAluPlugin_ALU_BITWISE_CTRL_lane1_1_string = "?????";
    endcase
  end
  always @(*) begin
    case(_zz_toplevel_execute_ctrl1_down_early1_IntAluPlugin_ALU_BITWISE_CTRL_lane1_2)
      IntAluPlugin_AluBitwiseCtrlEnum_XOR_1 : _zz_toplevel_execute_ctrl1_down_early1_IntAluPlugin_ALU_BITWISE_CTRL_lane1_2_string = "XOR_1";
      IntAluPlugin_AluBitwiseCtrlEnum_OR_1 : _zz_toplevel_execute_ctrl1_down_early1_IntAluPlugin_ALU_BITWISE_CTRL_lane1_2_string = "OR_1 ";
      IntAluPlugin_AluBitwiseCtrlEnum_AND_1 : _zz_toplevel_execute_ctrl1_down_early1_IntAluPlugin_ALU_BITWISE_CTRL_lane1_2_string = "AND_1";
      IntAluPlugin_AluBitwiseCtrlEnum_ZERO : _zz_toplevel_execute_ctrl1_down_early1_IntAluPlugin_ALU_BITWISE_CTRL_lane1_2_string = "ZERO ";
      default : _zz_toplevel_execute_ctrl1_down_early1_IntAluPlugin_ALU_BITWISE_CTRL_lane1_2_string = "?????";
    endcase
  end
  always @(*) begin
    case(_zz_toplevel_execute_ctrl1_down_BranchPlugin_BRANCH_CTRL_lane1)
      BranchPlugin_BranchCtrlEnum_B : _zz_toplevel_execute_ctrl1_down_BranchPlugin_BRANCH_CTRL_lane1_string = "B   ";
      BranchPlugin_BranchCtrlEnum_JAL : _zz_toplevel_execute_ctrl1_down_BranchPlugin_BRANCH_CTRL_lane1_string = "JAL ";
      BranchPlugin_BranchCtrlEnum_JALR : _zz_toplevel_execute_ctrl1_down_BranchPlugin_BRANCH_CTRL_lane1_string = "JALR";
      default : _zz_toplevel_execute_ctrl1_down_BranchPlugin_BRANCH_CTRL_lane1_string = "????";
    endcase
  end
  always @(*) begin
    case(_zz_toplevel_execute_ctrl1_down_BranchPlugin_BRANCH_CTRL_lane1_1)
      BranchPlugin_BranchCtrlEnum_B : _zz_toplevel_execute_ctrl1_down_BranchPlugin_BRANCH_CTRL_lane1_1_string = "B   ";
      BranchPlugin_BranchCtrlEnum_JAL : _zz_toplevel_execute_ctrl1_down_BranchPlugin_BRANCH_CTRL_lane1_1_string = "JAL ";
      BranchPlugin_BranchCtrlEnum_JALR : _zz_toplevel_execute_ctrl1_down_BranchPlugin_BRANCH_CTRL_lane1_1_string = "JALR";
      default : _zz_toplevel_execute_ctrl1_down_BranchPlugin_BRANCH_CTRL_lane1_1_string = "????";
    endcase
  end
  always @(*) begin
    case(_zz_toplevel_execute_ctrl1_down_BranchPlugin_BRANCH_CTRL_lane1_2)
      BranchPlugin_BranchCtrlEnum_B : _zz_toplevel_execute_ctrl1_down_BranchPlugin_BRANCH_CTRL_lane1_2_string = "B   ";
      BranchPlugin_BranchCtrlEnum_JAL : _zz_toplevel_execute_ctrl1_down_BranchPlugin_BRANCH_CTRL_lane1_2_string = "JAL ";
      BranchPlugin_BranchCtrlEnum_JALR : _zz_toplevel_execute_ctrl1_down_BranchPlugin_BRANCH_CTRL_lane1_2_string = "JALR";
      default : _zz_toplevel_execute_ctrl1_down_BranchPlugin_BRANCH_CTRL_lane1_2_string = "????";
    endcase
  end
  always @(*) begin
    case(_zz_toplevel_execute_ctrl1_down_late1_IntAluPlugin_ALU_BITWISE_CTRL_lane1_2)
      IntAluPlugin_AluBitwiseCtrlEnum_XOR_1 : _zz_toplevel_execute_ctrl1_down_late1_IntAluPlugin_ALU_BITWISE_CTRL_lane1_2_string = "XOR_1";
      IntAluPlugin_AluBitwiseCtrlEnum_OR_1 : _zz_toplevel_execute_ctrl1_down_late1_IntAluPlugin_ALU_BITWISE_CTRL_lane1_2_string = "OR_1 ";
      IntAluPlugin_AluBitwiseCtrlEnum_AND_1 : _zz_toplevel_execute_ctrl1_down_late1_IntAluPlugin_ALU_BITWISE_CTRL_lane1_2_string = "AND_1";
      IntAluPlugin_AluBitwiseCtrlEnum_ZERO : _zz_toplevel_execute_ctrl1_down_late1_IntAluPlugin_ALU_BITWISE_CTRL_lane1_2_string = "ZERO ";
      default : _zz_toplevel_execute_ctrl1_down_late1_IntAluPlugin_ALU_BITWISE_CTRL_lane1_2_string = "?????";
    endcase
  end
  always @(*) begin
    case(_zz_toplevel_execute_ctrl1_down_late1_IntAluPlugin_ALU_BITWISE_CTRL_lane1_3)
      IntAluPlugin_AluBitwiseCtrlEnum_XOR_1 : _zz_toplevel_execute_ctrl1_down_late1_IntAluPlugin_ALU_BITWISE_CTRL_lane1_3_string = "XOR_1";
      IntAluPlugin_AluBitwiseCtrlEnum_OR_1 : _zz_toplevel_execute_ctrl1_down_late1_IntAluPlugin_ALU_BITWISE_CTRL_lane1_3_string = "OR_1 ";
      IntAluPlugin_AluBitwiseCtrlEnum_AND_1 : _zz_toplevel_execute_ctrl1_down_late1_IntAluPlugin_ALU_BITWISE_CTRL_lane1_3_string = "AND_1";
      IntAluPlugin_AluBitwiseCtrlEnum_ZERO : _zz_toplevel_execute_ctrl1_down_late1_IntAluPlugin_ALU_BITWISE_CTRL_lane1_3_string = "ZERO ";
      default : _zz_toplevel_execute_ctrl1_down_late1_IntAluPlugin_ALU_BITWISE_CTRL_lane1_3_string = "?????";
    endcase
  end
  always @(*) begin
    case(_zz_toplevel_execute_ctrl1_down_late1_IntAluPlugin_ALU_BITWISE_CTRL_lane1_4)
      IntAluPlugin_AluBitwiseCtrlEnum_XOR_1 : _zz_toplevel_execute_ctrl1_down_late1_IntAluPlugin_ALU_BITWISE_CTRL_lane1_4_string = "XOR_1";
      IntAluPlugin_AluBitwiseCtrlEnum_OR_1 : _zz_toplevel_execute_ctrl1_down_late1_IntAluPlugin_ALU_BITWISE_CTRL_lane1_4_string = "OR_1 ";
      IntAluPlugin_AluBitwiseCtrlEnum_AND_1 : _zz_toplevel_execute_ctrl1_down_late1_IntAluPlugin_ALU_BITWISE_CTRL_lane1_4_string = "AND_1";
      IntAluPlugin_AluBitwiseCtrlEnum_ZERO : _zz_toplevel_execute_ctrl1_down_late1_IntAluPlugin_ALU_BITWISE_CTRL_lane1_4_string = "ZERO ";
      default : _zz_toplevel_execute_ctrl1_down_late1_IntAluPlugin_ALU_BITWISE_CTRL_lane1_4_string = "?????";
    endcase
  end
  always @(*) begin
    case(LsuPlugin_logic_flusher_stateReg)
      LsuPlugin_logic_flusher_enumDef_IDLE : LsuPlugin_logic_flusher_stateReg_string = "IDLE      ";
      LsuPlugin_logic_flusher_enumDef_CMD : LsuPlugin_logic_flusher_stateReg_string = "CMD       ";
      LsuPlugin_logic_flusher_enumDef_COMPLETION : LsuPlugin_logic_flusher_stateReg_string = "COMPLETION";
      default : LsuPlugin_logic_flusher_stateReg_string = "??????????";
    endcase
  end
  always @(*) begin
    case(LsuPlugin_logic_flusher_stateNext)
      LsuPlugin_logic_flusher_enumDef_IDLE : LsuPlugin_logic_flusher_stateNext_string = "IDLE      ";
      LsuPlugin_logic_flusher_enumDef_CMD : LsuPlugin_logic_flusher_stateNext_string = "CMD       ";
      LsuPlugin_logic_flusher_enumDef_COMPLETION : LsuPlugin_logic_flusher_stateNext_string = "COMPLETION";
      default : LsuPlugin_logic_flusher_stateNext_string = "??????????";
    endcase
  end
  always @(*) begin
    case(TrapPlugin_logic_harts_0_trap_fsm_stateReg)
      TrapPlugin_logic_harts_0_trap_fsm_enumDef_RESET : TrapPlugin_logic_harts_0_trap_fsm_stateReg_string = "RESET      ";
      TrapPlugin_logic_harts_0_trap_fsm_enumDef_RUNNING : TrapPlugin_logic_harts_0_trap_fsm_stateReg_string = "RUNNING    ";
      TrapPlugin_logic_harts_0_trap_fsm_enumDef_PROCESS_1 : TrapPlugin_logic_harts_0_trap_fsm_stateReg_string = "PROCESS_1  ";
      TrapPlugin_logic_harts_0_trap_fsm_enumDef_TRAP_EPC : TrapPlugin_logic_harts_0_trap_fsm_stateReg_string = "TRAP_EPC   ";
      TrapPlugin_logic_harts_0_trap_fsm_enumDef_TRAP_TVAL : TrapPlugin_logic_harts_0_trap_fsm_stateReg_string = "TRAP_TVAL  ";
      TrapPlugin_logic_harts_0_trap_fsm_enumDef_TRAP_TVEC : TrapPlugin_logic_harts_0_trap_fsm_stateReg_string = "TRAP_TVEC  ";
      TrapPlugin_logic_harts_0_trap_fsm_enumDef_TRAP_APPLY : TrapPlugin_logic_harts_0_trap_fsm_stateReg_string = "TRAP_APPLY ";
      TrapPlugin_logic_harts_0_trap_fsm_enumDef_XRET_EPC : TrapPlugin_logic_harts_0_trap_fsm_stateReg_string = "XRET_EPC   ";
      TrapPlugin_logic_harts_0_trap_fsm_enumDef_XRET_APPLY : TrapPlugin_logic_harts_0_trap_fsm_stateReg_string = "XRET_APPLY ";
      TrapPlugin_logic_harts_0_trap_fsm_enumDef_ATS_RSP : TrapPlugin_logic_harts_0_trap_fsm_stateReg_string = "ATS_RSP    ";
      TrapPlugin_logic_harts_0_trap_fsm_enumDef_JUMP : TrapPlugin_logic_harts_0_trap_fsm_stateReg_string = "JUMP       ";
      TrapPlugin_logic_harts_0_trap_fsm_enumDef_LSU_FLUSH : TrapPlugin_logic_harts_0_trap_fsm_stateReg_string = "LSU_FLUSH  ";
      TrapPlugin_logic_harts_0_trap_fsm_enumDef_FETCH_FLUSH : TrapPlugin_logic_harts_0_trap_fsm_stateReg_string = "FETCH_FLUSH";
      default : TrapPlugin_logic_harts_0_trap_fsm_stateReg_string = "???????????";
    endcase
  end
  always @(*) begin
    case(TrapPlugin_logic_harts_0_trap_fsm_stateNext)
      TrapPlugin_logic_harts_0_trap_fsm_enumDef_RESET : TrapPlugin_logic_harts_0_trap_fsm_stateNext_string = "RESET      ";
      TrapPlugin_logic_harts_0_trap_fsm_enumDef_RUNNING : TrapPlugin_logic_harts_0_trap_fsm_stateNext_string = "RUNNING    ";
      TrapPlugin_logic_harts_0_trap_fsm_enumDef_PROCESS_1 : TrapPlugin_logic_harts_0_trap_fsm_stateNext_string = "PROCESS_1  ";
      TrapPlugin_logic_harts_0_trap_fsm_enumDef_TRAP_EPC : TrapPlugin_logic_harts_0_trap_fsm_stateNext_string = "TRAP_EPC   ";
      TrapPlugin_logic_harts_0_trap_fsm_enumDef_TRAP_TVAL : TrapPlugin_logic_harts_0_trap_fsm_stateNext_string = "TRAP_TVAL  ";
      TrapPlugin_logic_harts_0_trap_fsm_enumDef_TRAP_TVEC : TrapPlugin_logic_harts_0_trap_fsm_stateNext_string = "TRAP_TVEC  ";
      TrapPlugin_logic_harts_0_trap_fsm_enumDef_TRAP_APPLY : TrapPlugin_logic_harts_0_trap_fsm_stateNext_string = "TRAP_APPLY ";
      TrapPlugin_logic_harts_0_trap_fsm_enumDef_XRET_EPC : TrapPlugin_logic_harts_0_trap_fsm_stateNext_string = "XRET_EPC   ";
      TrapPlugin_logic_harts_0_trap_fsm_enumDef_XRET_APPLY : TrapPlugin_logic_harts_0_trap_fsm_stateNext_string = "XRET_APPLY ";
      TrapPlugin_logic_harts_0_trap_fsm_enumDef_ATS_RSP : TrapPlugin_logic_harts_0_trap_fsm_stateNext_string = "ATS_RSP    ";
      TrapPlugin_logic_harts_0_trap_fsm_enumDef_JUMP : TrapPlugin_logic_harts_0_trap_fsm_stateNext_string = "JUMP       ";
      TrapPlugin_logic_harts_0_trap_fsm_enumDef_LSU_FLUSH : TrapPlugin_logic_harts_0_trap_fsm_stateNext_string = "LSU_FLUSH  ";
      TrapPlugin_logic_harts_0_trap_fsm_enumDef_FETCH_FLUSH : TrapPlugin_logic_harts_0_trap_fsm_stateNext_string = "FETCH_FLUSH";
      default : TrapPlugin_logic_harts_0_trap_fsm_stateNext_string = "???????????";
    endcase
  end
  always @(*) begin
    case(MmuPlugin_logic_refill_stateReg)
      MmuPlugin_logic_refill_enumDef_BOOT : MmuPlugin_logic_refill_stateReg_string = "BOOT ";
      MmuPlugin_logic_refill_enumDef_IDLE : MmuPlugin_logic_refill_stateReg_string = "IDLE ";
      MmuPlugin_logic_refill_enumDef_CMD_0 : MmuPlugin_logic_refill_stateReg_string = "CMD_0";
      MmuPlugin_logic_refill_enumDef_CMD_1 : MmuPlugin_logic_refill_stateReg_string = "CMD_1";
      MmuPlugin_logic_refill_enumDef_RSP_0 : MmuPlugin_logic_refill_stateReg_string = "RSP_0";
      MmuPlugin_logic_refill_enumDef_RSP_1 : MmuPlugin_logic_refill_stateReg_string = "RSP_1";
      default : MmuPlugin_logic_refill_stateReg_string = "?????";
    endcase
  end
  always @(*) begin
    case(MmuPlugin_logic_refill_stateNext)
      MmuPlugin_logic_refill_enumDef_BOOT : MmuPlugin_logic_refill_stateNext_string = "BOOT ";
      MmuPlugin_logic_refill_enumDef_IDLE : MmuPlugin_logic_refill_stateNext_string = "IDLE ";
      MmuPlugin_logic_refill_enumDef_CMD_0 : MmuPlugin_logic_refill_stateNext_string = "CMD_0";
      MmuPlugin_logic_refill_enumDef_CMD_1 : MmuPlugin_logic_refill_stateNext_string = "CMD_1";
      MmuPlugin_logic_refill_enumDef_RSP_0 : MmuPlugin_logic_refill_stateNext_string = "RSP_0";
      MmuPlugin_logic_refill_enumDef_RSP_1 : MmuPlugin_logic_refill_stateNext_string = "RSP_1";
      default : MmuPlugin_logic_refill_stateNext_string = "?????";
    endcase
  end
  always @(*) begin
    case(CsrAccessPlugin_logic_fsm_stateReg)
      CsrAccessPlugin_logic_fsm_enumDef_IDLE : CsrAccessPlugin_logic_fsm_stateReg_string = "IDLE      ";
      CsrAccessPlugin_logic_fsm_enumDef_READ : CsrAccessPlugin_logic_fsm_stateReg_string = "READ      ";
      CsrAccessPlugin_logic_fsm_enumDef_WRITE : CsrAccessPlugin_logic_fsm_stateReg_string = "WRITE     ";
      CsrAccessPlugin_logic_fsm_enumDef_COMPLETION : CsrAccessPlugin_logic_fsm_stateReg_string = "COMPLETION";
      default : CsrAccessPlugin_logic_fsm_stateReg_string = "??????????";
    endcase
  end
  always @(*) begin
    case(CsrAccessPlugin_logic_fsm_stateNext)
      CsrAccessPlugin_logic_fsm_enumDef_IDLE : CsrAccessPlugin_logic_fsm_stateNext_string = "IDLE      ";
      CsrAccessPlugin_logic_fsm_enumDef_READ : CsrAccessPlugin_logic_fsm_stateNext_string = "READ      ";
      CsrAccessPlugin_logic_fsm_enumDef_WRITE : CsrAccessPlugin_logic_fsm_stateNext_string = "WRITE     ";
      CsrAccessPlugin_logic_fsm_enumDef_COMPLETION : CsrAccessPlugin_logic_fsm_stateNext_string = "COMPLETION";
      default : CsrAccessPlugin_logic_fsm_stateNext_string = "??????????";
    endcase
  end
  `endif

  always @(*) begin
    BtbPlugin_logic_ras_ptr_pop_aheadValue = BtbPlugin_logic_ras_ptr_pop;
    BtbPlugin_logic_ras_ptr_pop_aheadValue = (_zz_BtbPlugin_logic_ras_ptr_pop_aheadValue - _zz_BtbPlugin_logic_ras_ptr_pop_aheadValue_3);
  end

  assign toplevel_execute_ctrl4_down_RD_ENABLE_lane1 = toplevel_execute_ctrl4_RD_ENABLE_lane1_bypass;
  always @(*) begin
    toplevel_execute_ctrl4_RD_ENABLE_lane1_bypass = toplevel_execute_ctrl4_up_RD_ENABLE_lane1;
    if(when_ExecuteLanePlugin_l300_9) begin
      toplevel_execute_ctrl4_RD_ENABLE_lane1_bypass = 1'b0;
    end
  end

  assign toplevel_execute_ctrl4_down_LANE_SEL_lane1 = toplevel_execute_ctrl4_LANE_SEL_lane1_bypass;
  always @(*) begin
    toplevel_execute_ctrl4_LANE_SEL_lane1_bypass = toplevel_execute_ctrl4_up_LANE_SEL_lane1;
    if(when_ExecuteLanePlugin_l300_9) begin
      toplevel_execute_ctrl4_LANE_SEL_lane1_bypass = 1'b0;
    end
  end

  assign toplevel_execute_ctrl3_down_RD_ENABLE_lane1 = toplevel_execute_ctrl3_RD_ENABLE_lane1_bypass;
  always @(*) begin
    toplevel_execute_ctrl3_RD_ENABLE_lane1_bypass = toplevel_execute_ctrl3_up_RD_ENABLE_lane1;
    if(when_ExecuteLanePlugin_l300_8) begin
      toplevel_execute_ctrl3_RD_ENABLE_lane1_bypass = 1'b0;
    end
  end

  assign toplevel_execute_ctrl3_down_LANE_SEL_lane1 = toplevel_execute_ctrl3_LANE_SEL_lane1_bypass;
  always @(*) begin
    toplevel_execute_ctrl3_LANE_SEL_lane1_bypass = toplevel_execute_ctrl3_up_LANE_SEL_lane1;
    if(when_ExecuteLanePlugin_l300_8) begin
      toplevel_execute_ctrl3_LANE_SEL_lane1_bypass = 1'b0;
    end
  end

  assign toplevel_execute_ctrl2_down_RD_ENABLE_lane1 = toplevel_execute_ctrl2_RD_ENABLE_lane1_bypass;
  always @(*) begin
    toplevel_execute_ctrl2_RD_ENABLE_lane1_bypass = toplevel_execute_ctrl2_up_RD_ENABLE_lane1;
    if(when_ExecuteLanePlugin_l300_7) begin
      toplevel_execute_ctrl2_RD_ENABLE_lane1_bypass = 1'b0;
    end
  end

  assign toplevel_execute_ctrl2_down_LANE_SEL_lane1 = toplevel_execute_ctrl2_LANE_SEL_lane1_bypass;
  always @(*) begin
    toplevel_execute_ctrl2_LANE_SEL_lane1_bypass = toplevel_execute_ctrl2_up_LANE_SEL_lane1;
    if(when_ExecuteLanePlugin_l300_7) begin
      toplevel_execute_ctrl2_LANE_SEL_lane1_bypass = 1'b0;
    end
  end

  assign toplevel_execute_ctrl1_down_RD_ENABLE_lane1 = toplevel_execute_ctrl1_RD_ENABLE_lane1_bypass;
  always @(*) begin
    toplevel_execute_ctrl1_RD_ENABLE_lane1_bypass = toplevel_execute_ctrl1_up_RD_ENABLE_lane1;
    if(when_ExecuteLanePlugin_l300_6) begin
      toplevel_execute_ctrl1_RD_ENABLE_lane1_bypass = 1'b0;
    end
  end

  assign toplevel_execute_ctrl1_down_LANE_SEL_lane1 = toplevel_execute_ctrl1_LANE_SEL_lane1_bypass;
  always @(*) begin
    toplevel_execute_ctrl1_LANE_SEL_lane1_bypass = toplevel_execute_ctrl1_up_LANE_SEL_lane1;
    if(when_ExecuteLanePlugin_l300_6) begin
      toplevel_execute_ctrl1_LANE_SEL_lane1_bypass = 1'b0;
    end
  end

  assign toplevel_execute_ctrl0_down_RD_ENABLE_lane1 = toplevel_execute_ctrl0_RD_ENABLE_lane1_bypass;
  always @(*) begin
    toplevel_execute_ctrl0_RD_ENABLE_lane1_bypass = toplevel_execute_ctrl0_up_RD_ENABLE_lane1;
    if(when_ExecuteLanePlugin_l300_5) begin
      toplevel_execute_ctrl0_RD_ENABLE_lane1_bypass = 1'b0;
    end
  end

  assign toplevel_execute_ctrl0_down_LANE_SEL_lane1 = toplevel_execute_ctrl0_LANE_SEL_lane1_bypass;
  always @(*) begin
    toplevel_execute_ctrl0_LANE_SEL_lane1_bypass = toplevel_execute_ctrl0_up_LANE_SEL_lane1;
    if(when_ExecuteLanePlugin_l300_5) begin
      toplevel_execute_ctrl0_LANE_SEL_lane1_bypass = 1'b0;
    end
  end

  assign toplevel_execute_ctrl3_down_integer_RS2_lane1 = toplevel_execute_ctrl3_integer_RS2_lane1_bypass;
  assign toplevel_execute_ctrl2_down_integer_RS2_lane1 = toplevel_execute_ctrl2_integer_RS2_lane1_bypass;
  assign toplevel_execute_ctrl3_down_integer_RS1_lane1 = toplevel_execute_ctrl3_integer_RS1_lane1_bypass;
  assign toplevel_execute_ctrl2_down_integer_RS1_lane1 = toplevel_execute_ctrl2_integer_RS1_lane1_bypass;
  assign toplevel_execute_ctrl4_down_RD_ENABLE_lane0 = toplevel_execute_ctrl4_RD_ENABLE_lane0_bypass;
  always @(*) begin
    toplevel_execute_ctrl4_RD_ENABLE_lane0_bypass = toplevel_execute_ctrl4_up_RD_ENABLE_lane0;
    if(when_ExecuteLanePlugin_l300_4) begin
      toplevel_execute_ctrl4_RD_ENABLE_lane0_bypass = 1'b0;
    end
  end

  assign toplevel_execute_ctrl4_down_LANE_SEL_lane0 = toplevel_execute_ctrl4_LANE_SEL_lane0_bypass;
  always @(*) begin
    toplevel_execute_ctrl4_LANE_SEL_lane0_bypass = toplevel_execute_ctrl4_up_LANE_SEL_lane0;
    if(when_ExecuteLanePlugin_l300_4) begin
      toplevel_execute_ctrl4_LANE_SEL_lane0_bypass = 1'b0;
    end
  end

  assign toplevel_execute_ctrl3_down_RD_ENABLE_lane0 = toplevel_execute_ctrl3_RD_ENABLE_lane0_bypass;
  always @(*) begin
    toplevel_execute_ctrl3_RD_ENABLE_lane0_bypass = toplevel_execute_ctrl3_up_RD_ENABLE_lane0;
    if(when_ExecuteLanePlugin_l300_3) begin
      toplevel_execute_ctrl3_RD_ENABLE_lane0_bypass = 1'b0;
    end
  end

  assign toplevel_execute_ctrl3_down_LANE_SEL_lane0 = toplevel_execute_ctrl3_LANE_SEL_lane0_bypass;
  always @(*) begin
    toplevel_execute_ctrl3_LANE_SEL_lane0_bypass = toplevel_execute_ctrl3_up_LANE_SEL_lane0;
    if(when_ExecuteLanePlugin_l300_3) begin
      toplevel_execute_ctrl3_LANE_SEL_lane0_bypass = 1'b0;
    end
  end

  assign toplevel_execute_ctrl2_down_RD_ENABLE_lane0 = toplevel_execute_ctrl2_RD_ENABLE_lane0_bypass;
  always @(*) begin
    toplevel_execute_ctrl2_RD_ENABLE_lane0_bypass = toplevel_execute_ctrl2_up_RD_ENABLE_lane0;
    if(when_ExecuteLanePlugin_l300_2) begin
      toplevel_execute_ctrl2_RD_ENABLE_lane0_bypass = 1'b0;
    end
  end

  assign toplevel_execute_ctrl2_down_LANE_SEL_lane0 = toplevel_execute_ctrl2_LANE_SEL_lane0_bypass;
  always @(*) begin
    toplevel_execute_ctrl2_LANE_SEL_lane0_bypass = toplevel_execute_ctrl2_up_LANE_SEL_lane0;
    if(when_ExecuteLanePlugin_l300_2) begin
      toplevel_execute_ctrl2_LANE_SEL_lane0_bypass = 1'b0;
    end
  end

  assign toplevel_execute_ctrl1_down_RD_ENABLE_lane0 = toplevel_execute_ctrl1_RD_ENABLE_lane0_bypass;
  always @(*) begin
    toplevel_execute_ctrl1_RD_ENABLE_lane0_bypass = toplevel_execute_ctrl1_up_RD_ENABLE_lane0;
    if(when_ExecuteLanePlugin_l300_1) begin
      toplevel_execute_ctrl1_RD_ENABLE_lane0_bypass = 1'b0;
    end
  end

  assign toplevel_execute_ctrl1_down_LANE_SEL_lane0 = toplevel_execute_ctrl1_LANE_SEL_lane0_bypass;
  always @(*) begin
    toplevel_execute_ctrl1_LANE_SEL_lane0_bypass = toplevel_execute_ctrl1_up_LANE_SEL_lane0;
    if(when_ExecuteLanePlugin_l300_1) begin
      toplevel_execute_ctrl1_LANE_SEL_lane0_bypass = 1'b0;
    end
  end

  assign toplevel_execute_ctrl0_down_RD_ENABLE_lane0 = toplevel_execute_ctrl0_RD_ENABLE_lane0_bypass;
  always @(*) begin
    toplevel_execute_ctrl0_RD_ENABLE_lane0_bypass = toplevel_execute_ctrl0_up_RD_ENABLE_lane0;
    if(when_ExecuteLanePlugin_l300) begin
      toplevel_execute_ctrl0_RD_ENABLE_lane0_bypass = 1'b0;
    end
  end

  assign toplevel_execute_ctrl0_down_LANE_SEL_lane0 = toplevel_execute_ctrl0_LANE_SEL_lane0_bypass;
  always @(*) begin
    toplevel_execute_ctrl0_LANE_SEL_lane0_bypass = toplevel_execute_ctrl0_up_LANE_SEL_lane0;
    if(when_ExecuteLanePlugin_l300) begin
      toplevel_execute_ctrl0_LANE_SEL_lane0_bypass = 1'b0;
    end
  end

  assign toplevel_execute_ctrl3_down_integer_RS2_lane0 = toplevel_execute_ctrl3_integer_RS2_lane0_bypass;
  assign toplevel_execute_ctrl2_down_integer_RS2_lane0 = toplevel_execute_ctrl2_integer_RS2_lane0_bypass;
  assign toplevel_execute_ctrl3_down_integer_RS1_lane0 = toplevel_execute_ctrl3_integer_RS1_lane0_bypass;
  assign toplevel_execute_ctrl2_down_integer_RS1_lane0 = toplevel_execute_ctrl2_integer_RS1_lane0_bypass;
  always @(*) begin
    _zz_2 = 1'b0;
    if(CsrRamPlugin_logic_writeLogic_port_valid) begin
      _zz_2 = 1'b1;
    end
  end

  assign toplevel_execute_ctrl4_down_COMMIT_lane0 = toplevel_execute_ctrl4_COMMIT_lane0_bypass;
  always @(*) begin
    toplevel_execute_ctrl4_COMMIT_lane0_bypass = toplevel_execute_ctrl4_up_COMMIT_lane0;
    if(when_LsuPlugin_l723) begin
      if(LsuPlugin_logic_onCtrl_lsuTrap) begin
        toplevel_execute_ctrl4_COMMIT_lane0_bypass = 1'b0;
      end
    end
  end

  assign toplevel_execute_ctrl4_down_TRAP_lane0 = toplevel_execute_ctrl4_TRAP_lane0_bypass;
  always @(*) begin
    toplevel_execute_ctrl4_TRAP_lane0_bypass = toplevel_execute_ctrl4_up_TRAP_lane0;
    if(when_LsuPlugin_l723) begin
      if(LsuPlugin_logic_onCtrl_lsuTrap) begin
        toplevel_execute_ctrl4_TRAP_lane0_bypass = 1'b1;
      end
    end
  end

  assign toplevel_execute_ctrl4_down_LsuL1_SEL_lane0 = toplevel_execute_ctrl4_LsuL1_SEL_lane0_bypass;
  always @(*) begin
    toplevel_execute_ctrl4_LsuL1_SEL_lane0_bypass = toplevel_execute_ctrl4_up_LsuL1_SEL_lane0;
    if(when_LsuPlugin_l449_1) begin
      toplevel_execute_ctrl4_LsuL1_SEL_lane0_bypass = 1'b0;
    end
  end

  assign toplevel_execute_ctrl3_down_LsuL1_SEL_lane0 = toplevel_execute_ctrl3_LsuL1_SEL_lane0_bypass;
  always @(*) begin
    toplevel_execute_ctrl3_LsuL1_SEL_lane0_bypass = toplevel_execute_ctrl3_up_LsuL1_SEL_lane0;
    if(when_LsuPlugin_l449) begin
      toplevel_execute_ctrl3_LsuL1_SEL_lane0_bypass = 1'b0;
    end
  end

  assign toplevel_execute_ctrl3_down_LsuL1Plugin_logic_SHARED_lane0_plru_0 = toplevel_execute_ctrl3_LsuL1Plugin_logic_SHARED_lane0_bypass_plru_0;
  assign toplevel_execute_ctrl3_down_LsuL1Plugin_logic_SHARED_lane0_dirty = toplevel_execute_ctrl3_LsuL1Plugin_logic_SHARED_lane0_bypass_dirty;
  always @(*) begin
    _zz_3 = 1'b0;
    if(LsuL1Plugin_logic_writeback_read_slotReadLast_valid) begin
      _zz_3 = 1'b1;
    end
  end

  always @(*) begin
    _zz_4 = 1'b0;
    if(LsuL1Plugin_logic_shared_write_valid) begin
      _zz_4 = 1'b1;
    end
  end

  assign toplevel_decode_ctrls_1_down_LANE_SEL_1 = toplevel_decode_ctrls_1_LANE_SEL_1_bypass;
  always @(*) begin
    toplevel_decode_ctrls_1_LANE_SEL_1_bypass = toplevel_decode_ctrls_1_up_LANE_SEL_1;
    if(decode_logic_flushes_1_onLanes_1_doIt) begin
      toplevel_decode_ctrls_1_LANE_SEL_1_bypass = 1'b0;
    end
  end

  assign toplevel_decode_ctrls_1_down_LANE_SEL_0 = toplevel_decode_ctrls_1_LANE_SEL_0_bypass;
  always @(*) begin
    toplevel_decode_ctrls_1_LANE_SEL_0_bypass = toplevel_decode_ctrls_1_up_LANE_SEL_0;
    if(decode_logic_flushes_1_onLanes_0_doIt) begin
      toplevel_decode_ctrls_1_LANE_SEL_0_bypass = 1'b0;
    end
  end

  assign toplevel_decode_ctrls_0_down_LANE_SEL_1 = toplevel_decode_ctrls_0_LANE_SEL_1_bypass;
  always @(*) begin
    toplevel_decode_ctrls_0_LANE_SEL_1_bypass = toplevel_decode_ctrls_0_up_LANE_SEL_1;
    if(decode_logic_flushes_0_onLanes_1_doIt) begin
      toplevel_decode_ctrls_0_LANE_SEL_1_bypass = 1'b0;
    end
  end

  assign toplevel_decode_ctrls_0_down_LANE_SEL_0 = toplevel_decode_ctrls_0_LANE_SEL_0_bypass;
  always @(*) begin
    toplevel_decode_ctrls_0_LANE_SEL_0_bypass = toplevel_decode_ctrls_0_up_LANE_SEL_0;
    if(decode_logic_flushes_0_onLanes_0_doIt) begin
      toplevel_decode_ctrls_0_LANE_SEL_0_bypass = 1'b0;
    end
  end

  assign toplevel_execute_ctrl4_down_lane1_integer_WriteBackPlugin_logic_DATA_lane1 = toplevel_execute_ctrl4_lane1_integer_WriteBackPlugin_logic_DATA_lane1_bypass;
  assign toplevel_execute_ctrl3_down_lane1_integer_WriteBackPlugin_logic_DATA_lane1 = toplevel_execute_ctrl3_lane1_integer_WriteBackPlugin_logic_DATA_lane1_bypass;
  assign toplevel_execute_ctrl2_down_lane1_integer_WriteBackPlugin_logic_DATA_lane1 = toplevel_execute_ctrl2_lane1_integer_WriteBackPlugin_logic_DATA_lane1_bypass;
  assign toplevel_execute_ctrl4_down_lane0_integer_WriteBackPlugin_logic_DATA_lane0 = toplevel_execute_ctrl4_lane0_integer_WriteBackPlugin_logic_DATA_lane0_bypass;
  assign toplevel_execute_ctrl3_down_lane0_integer_WriteBackPlugin_logic_DATA_lane0 = toplevel_execute_ctrl3_lane0_integer_WriteBackPlugin_logic_DATA_lane0_bypass;
  assign toplevel_execute_ctrl2_down_lane0_integer_WriteBackPlugin_logic_DATA_lane0 = toplevel_execute_ctrl2_lane0_integer_WriteBackPlugin_logic_DATA_lane0_bypass;
  assign toplevel_decode_ctrls_1_down_TRAP_1 = toplevel_decode_ctrls_1_TRAP_1_bypass;
  always @(*) begin
    toplevel_decode_ctrls_1_TRAP_1_bypass = toplevel_decode_ctrls_1_up_TRAP_1;
    if(when_DecoderPlugin_l216_1) begin
      toplevel_decode_ctrls_1_TRAP_1_bypass = 1'b1;
    end
  end

  assign toplevel_decode_ctrls_1_down_TRAP_0 = toplevel_decode_ctrls_1_TRAP_0_bypass;
  always @(*) begin
    toplevel_decode_ctrls_1_TRAP_0_bypass = toplevel_decode_ctrls_1_up_TRAP_0;
    if(when_DecoderPlugin_l216) begin
      toplevel_decode_ctrls_1_TRAP_0_bypass = 1'b1;
    end
  end

  assign toplevel_execute_ctrl4_down_COMPLETED_lane0 = toplevel_execute_ctrl4_COMPLETED_lane0_bypass;
  assign toplevel_execute_ctrl3_down_COMPLETED_lane0 = toplevel_execute_ctrl3_COMPLETED_lane0_bypass;
  assign toplevel_execute_ctrl2_down_COMPLETED_lane0 = toplevel_execute_ctrl2_COMPLETED_lane0_bypass;
  assign toplevel_execute_ctrl4_down_COMPLETED_lane1 = toplevel_execute_ctrl4_COMPLETED_lane1_bypass;
  assign toplevel_execute_ctrl3_down_COMPLETED_lane1 = toplevel_execute_ctrl3_COMPLETED_lane1_bypass;
  assign toplevel_execute_ctrl2_down_COMPLETED_lane1 = toplevel_execute_ctrl2_COMPLETED_lane1_bypass;
  always @(*) begin
    late1_BranchPlugin_logic_jumpLogic_history_fromFetch_shifter_4 = late1_BranchPlugin_logic_jumpLogic_history_fromFetch_shifter_3;
    if(when_BranchPlugin_l210_3) begin
      late1_BranchPlugin_logic_jumpLogic_history_fromFetch_shifter_4 = _zz_late1_BranchPlugin_logic_jumpLogic_history_fromFetch_shifter_4[11 : 0];
    end
  end

  always @(*) begin
    late1_BranchPlugin_logic_jumpLogic_history_fromFetch_shifter_3 = late1_BranchPlugin_logic_jumpLogic_history_fromFetch_shifter_2;
    if(when_BranchPlugin_l206_11) begin
      late1_BranchPlugin_logic_jumpLogic_history_fromFetch_shifter_3 = _zz_late1_BranchPlugin_logic_jumpLogic_history_fromFetch_shifter_3[11 : 0];
    end
  end

  always @(*) begin
    late1_BranchPlugin_logic_jumpLogic_history_fromFetch_shifter_2 = late1_BranchPlugin_logic_jumpLogic_history_fromFetch_shifter_1;
    if(when_BranchPlugin_l206_10) begin
      late1_BranchPlugin_logic_jumpLogic_history_fromFetch_shifter_2 = _zz_late1_BranchPlugin_logic_jumpLogic_history_fromFetch_shifter_2[11 : 0];
    end
  end

  always @(*) begin
    late1_BranchPlugin_logic_jumpLogic_history_fromFetch_shifter_1 = late1_BranchPlugin_logic_jumpLogic_history_fromFetch_shifter;
    if(when_BranchPlugin_l206_9) begin
      late1_BranchPlugin_logic_jumpLogic_history_fromFetch_shifter_1 = _zz_late1_BranchPlugin_logic_jumpLogic_history_fromFetch_shifter_1[11 : 0];
    end
  end

  always @(*) begin
    late0_BranchPlugin_logic_jumpLogic_history_fromFetch_shifter_4 = late0_BranchPlugin_logic_jumpLogic_history_fromFetch_shifter_3;
    if(when_BranchPlugin_l210_2) begin
      late0_BranchPlugin_logic_jumpLogic_history_fromFetch_shifter_4 = _zz_late0_BranchPlugin_logic_jumpLogic_history_fromFetch_shifter_4[11 : 0];
    end
  end

  always @(*) begin
    late0_BranchPlugin_logic_jumpLogic_history_fromFetch_shifter_3 = late0_BranchPlugin_logic_jumpLogic_history_fromFetch_shifter_2;
    if(when_BranchPlugin_l206_8) begin
      late0_BranchPlugin_logic_jumpLogic_history_fromFetch_shifter_3 = _zz_late0_BranchPlugin_logic_jumpLogic_history_fromFetch_shifter_3[11 : 0];
    end
  end

  always @(*) begin
    late0_BranchPlugin_logic_jumpLogic_history_fromFetch_shifter_2 = late0_BranchPlugin_logic_jumpLogic_history_fromFetch_shifter_1;
    if(when_BranchPlugin_l206_7) begin
      late0_BranchPlugin_logic_jumpLogic_history_fromFetch_shifter_2 = _zz_late0_BranchPlugin_logic_jumpLogic_history_fromFetch_shifter_2[11 : 0];
    end
  end

  always @(*) begin
    late0_BranchPlugin_logic_jumpLogic_history_fromFetch_shifter_1 = late0_BranchPlugin_logic_jumpLogic_history_fromFetch_shifter;
    if(when_BranchPlugin_l206_6) begin
      late0_BranchPlugin_logic_jumpLogic_history_fromFetch_shifter_1 = _zz_late0_BranchPlugin_logic_jumpLogic_history_fromFetch_shifter_1[11 : 0];
    end
  end

  always @(*) begin
    early1_BranchPlugin_logic_jumpLogic_history_fromFetch_shifter_4 = early1_BranchPlugin_logic_jumpLogic_history_fromFetch_shifter_3;
    if(when_BranchPlugin_l210_1) begin
      early1_BranchPlugin_logic_jumpLogic_history_fromFetch_shifter_4 = _zz_early1_BranchPlugin_logic_jumpLogic_history_fromFetch_shifter_4[11 : 0];
    end
  end

  always @(*) begin
    early1_BranchPlugin_logic_jumpLogic_history_fromFetch_shifter_3 = early1_BranchPlugin_logic_jumpLogic_history_fromFetch_shifter_2;
    if(when_BranchPlugin_l206_5) begin
      early1_BranchPlugin_logic_jumpLogic_history_fromFetch_shifter_3 = _zz_early1_BranchPlugin_logic_jumpLogic_history_fromFetch_shifter_3[11 : 0];
    end
  end

  always @(*) begin
    early1_BranchPlugin_logic_jumpLogic_history_fromFetch_shifter_2 = early1_BranchPlugin_logic_jumpLogic_history_fromFetch_shifter_1;
    if(when_BranchPlugin_l206_4) begin
      early1_BranchPlugin_logic_jumpLogic_history_fromFetch_shifter_2 = _zz_early1_BranchPlugin_logic_jumpLogic_history_fromFetch_shifter_2[11 : 0];
    end
  end

  always @(*) begin
    early1_BranchPlugin_logic_jumpLogic_history_fromFetch_shifter_1 = early1_BranchPlugin_logic_jumpLogic_history_fromFetch_shifter;
    if(when_BranchPlugin_l206_3) begin
      early1_BranchPlugin_logic_jumpLogic_history_fromFetch_shifter_1 = _zz_early1_BranchPlugin_logic_jumpLogic_history_fromFetch_shifter_1[11 : 0];
    end
  end

  assign toplevel_execute_ctrl2_down_COMMIT_lane0 = toplevel_execute_ctrl2_COMMIT_lane0_bypass;
  always @(*) begin
    toplevel_execute_ctrl2_COMMIT_lane0_bypass = toplevel_execute_ctrl2_up_COMMIT_lane0;
    if(when_EnvPlugin_l116) begin
      if(when_EnvPlugin_l120) begin
        toplevel_execute_ctrl2_COMMIT_lane0_bypass = 1'b0;
      end
    end
    case(CsrAccessPlugin_logic_fsm_stateReg)
      CsrAccessPlugin_logic_fsm_enumDef_READ : begin
      end
      CsrAccessPlugin_logic_fsm_enumDef_WRITE : begin
      end
      CsrAccessPlugin_logic_fsm_enumDef_COMPLETION : begin
      end
      default : begin
        if(CsrAccessPlugin_logic_fsm_inject_onDecodeDo) begin
          if(CsrAccessPlugin_logic_fsm_inject_sampled) begin
            if(CsrAccessPlugin_logic_fsm_inject_trapReg) begin
              toplevel_execute_ctrl2_COMMIT_lane0_bypass = 1'b0;
            end
          end
        end
      end
    endcase
  end

  assign toplevel_execute_ctrl2_down_TRAP_lane0 = toplevel_execute_ctrl2_TRAP_lane0_bypass;
  always @(*) begin
    toplevel_execute_ctrl2_TRAP_lane0_bypass = toplevel_execute_ctrl2_up_TRAP_lane0;
    if(when_EnvPlugin_l116) begin
      toplevel_execute_ctrl2_TRAP_lane0_bypass = 1'b1;
    end
    if(CsrAccessPlugin_logic_fsm_inject_flushReg) begin
      toplevel_execute_ctrl2_TRAP_lane0_bypass = 1'b1;
    end
    case(CsrAccessPlugin_logic_fsm_stateReg)
      CsrAccessPlugin_logic_fsm_enumDef_READ : begin
      end
      CsrAccessPlugin_logic_fsm_enumDef_WRITE : begin
      end
      CsrAccessPlugin_logic_fsm_enumDef_COMPLETION : begin
      end
      default : begin
        if(CsrAccessPlugin_logic_fsm_inject_onDecodeDo) begin
          if(CsrAccessPlugin_logic_fsm_inject_sampled) begin
            if(CsrAccessPlugin_logic_fsm_inject_trapReg) begin
              toplevel_execute_ctrl2_TRAP_lane0_bypass = 1'b1;
            end else begin
              if(CsrAccessPlugin_logic_fsm_inject_busTrapReg) begin
                toplevel_execute_ctrl2_TRAP_lane0_bypass = 1'b1;
              end
            end
          end
        end
      end
    endcase
  end

  always @(*) begin
    early0_BranchPlugin_logic_jumpLogic_history_fromFetch_shifter_4 = early0_BranchPlugin_logic_jumpLogic_history_fromFetch_shifter_3;
    if(when_BranchPlugin_l210) begin
      early0_BranchPlugin_logic_jumpLogic_history_fromFetch_shifter_4 = _zz_early0_BranchPlugin_logic_jumpLogic_history_fromFetch_shifter_4[11 : 0];
    end
  end

  always @(*) begin
    early0_BranchPlugin_logic_jumpLogic_history_fromFetch_shifter_3 = early0_BranchPlugin_logic_jumpLogic_history_fromFetch_shifter_2;
    if(when_BranchPlugin_l206_2) begin
      early0_BranchPlugin_logic_jumpLogic_history_fromFetch_shifter_3 = _zz_early0_BranchPlugin_logic_jumpLogic_history_fromFetch_shifter_3[11 : 0];
    end
  end

  always @(*) begin
    early0_BranchPlugin_logic_jumpLogic_history_fromFetch_shifter_2 = early0_BranchPlugin_logic_jumpLogic_history_fromFetch_shifter_1;
    if(when_BranchPlugin_l206_1) begin
      early0_BranchPlugin_logic_jumpLogic_history_fromFetch_shifter_2 = _zz_early0_BranchPlugin_logic_jumpLogic_history_fromFetch_shifter_2[11 : 0];
    end
  end

  always @(*) begin
    early0_BranchPlugin_logic_jumpLogic_history_fromFetch_shifter_1 = early0_BranchPlugin_logic_jumpLogic_history_fromFetch_shifter;
    if(when_BranchPlugin_l206) begin
      early0_BranchPlugin_logic_jumpLogic_history_fromFetch_shifter_1 = _zz_early0_BranchPlugin_logic_jumpLogic_history_fromFetch_shifter_1[11 : 0];
    end
  end

  always @(*) begin
    _zz_5 = 1'b0;
    if(BtbPlugin_logic_ras_write_valid) begin
      _zz_5 = 1'b1;
    end
  end

  always @(*) begin
    _zz_6 = 1'b0;
    if(GSharePlugin_logic_mem_write_valid) begin
      _zz_6 = 1'b1;
    end
  end

  always @(*) begin
    _zz_fetch_logic_ctrls_0_haltRequest_FetchL1Plugin_l233 = 1'b0;
    if(when_FetchL1Plugin_l232) begin
      _zz_fetch_logic_ctrls_0_haltRequest_FetchL1Plugin_l233 = 1'b1;
    end
  end

  always @(*) begin
    _zz_7 = 1'b0;
    if(FetchL1Plugin_logic_plru_write_valid) begin
      _zz_7 = 1'b1;
    end
  end

  always @(*) begin
    _zz_8 = 1'b0;
    if(FetchL1Plugin_logic_banks_1_write_valid) begin
      _zz_8 = 1'b1;
    end
  end

  always @(*) begin
    _zz_9 = 1'b0;
    if(FetchL1Plugin_logic_banks_0_write_valid) begin
      _zz_9 = 1'b1;
    end
  end

  assign AlignerPlugin_api_singleFetch = 1'b0;
  assign AlignerPlugin_api_haltIt = 1'b0;
  always @(*) begin
    DispatchPlugin_api_haltDispatch = 1'b0;
    if(LsuPlugin_logic_onCtrl_hartRegulation_valid) begin
      DispatchPlugin_api_haltDispatch = 1'b1;
    end
  end

  assign CsrRamPlugin_api_holdRead = 1'b0;
  assign CsrRamPlugin_api_holdWrite = 1'b0;
  always @(*) begin
    TrapPlugin_api_harts_0_redo = 1'b0;
    case(TrapPlugin_logic_harts_0_trap_fsm_stateReg)
      TrapPlugin_logic_harts_0_trap_fsm_enumDef_RUNNING : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_enumDef_PROCESS_1 : begin
        if(!when_TrapPlugin_l393) begin
          case(TrapPlugin_logic_harts_0_trap_pending_state_code)
            4'b0000 : begin
            end
            4'b0001 : begin
            end
            4'b0010 : begin
            end
            4'b0100 : begin
              TrapPlugin_api_harts_0_redo = 1'b1;
            end
            4'b0101 : begin
            end
            4'b1000 : begin
            end
            4'b0110 : begin
            end
            4'b0111 : begin
            end
            default : begin
            end
          endcase
        end
      end
      TrapPlugin_logic_harts_0_trap_fsm_enumDef_TRAP_EPC : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_enumDef_TRAP_TVAL : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_enumDef_TRAP_TVEC : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_enumDef_TRAP_APPLY : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_enumDef_XRET_EPC : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_enumDef_XRET_APPLY : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_enumDef_ATS_RSP : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_enumDef_JUMP : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_enumDef_LSU_FLUSH : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_enumDef_FETCH_FLUSH : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    TrapPlugin_api_harts_0_askWake = 1'b0;
    if(when_TrapPlugin_l214) begin
      TrapPlugin_api_harts_0_askWake = 1'b1;
    end
  end

  always @(*) begin
    TrapPlugin_api_harts_0_rvTrap = 1'b0;
    case(TrapPlugin_logic_harts_0_trap_fsm_stateReg)
      TrapPlugin_logic_harts_0_trap_fsm_enumDef_RUNNING : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_enumDef_PROCESS_1 : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_enumDef_TRAP_EPC : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_enumDef_TRAP_TVAL : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_enumDef_TRAP_TVEC : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_enumDef_TRAP_APPLY : begin
        TrapPlugin_api_harts_0_rvTrap = 1'b1;
      end
      TrapPlugin_logic_harts_0_trap_fsm_enumDef_XRET_EPC : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_enumDef_XRET_APPLY : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_enumDef_ATS_RSP : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_enumDef_JUMP : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_enumDef_LSU_FLUSH : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_enumDef_FETCH_FLUSH : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    DecoderPlugin_logic_forgetPort_valid = 1'b0;
    if(DecoderPlugin_logic_laneLogic_0_fixer_doIt) begin
      DecoderPlugin_logic_forgetPort_valid = 1'b1;
    end
    if(DecoderPlugin_logic_laneLogic_1_fixer_doIt) begin
      DecoderPlugin_logic_forgetPort_valid = 1'b1;
    end
  end

  always @(*) begin
    DecoderPlugin_logic_forgetPort_payload_pcOnLastSlice = 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
    if(DecoderPlugin_logic_laneLogic_0_fixer_doIt) begin
      DecoderPlugin_logic_forgetPort_payload_pcOnLastSlice = (toplevel_decode_ctrls_1_down_PC_0 + _zz_DecoderPlugin_logic_forgetPort_payload_pcOnLastSlice);
    end
    if(DecoderPlugin_logic_laneLogic_1_fixer_doIt) begin
      DecoderPlugin_logic_forgetPort_payload_pcOnLastSlice = (toplevel_decode_ctrls_1_down_PC_1 + _zz_DecoderPlugin_logic_forgetPort_payload_pcOnLastSlice_3);
    end
  end

  always @(*) begin
    case(toplevel_execute_ctrl2_down_early0_IntAluPlugin_ALU_BITWISE_CTRL_lane0)
      IntAluPlugin_AluBitwiseCtrlEnum_AND_1 : begin
        early0_IntAluPlugin_logic_alu_bitwise = (toplevel_execute_ctrl2_down_early0_SrcPlugin_SRC1_lane0 & toplevel_execute_ctrl2_down_early0_SrcPlugin_SRC2_lane0);
      end
      IntAluPlugin_AluBitwiseCtrlEnum_OR_1 : begin
        early0_IntAluPlugin_logic_alu_bitwise = (toplevel_execute_ctrl2_down_early0_SrcPlugin_SRC1_lane0 | toplevel_execute_ctrl2_down_early0_SrcPlugin_SRC2_lane0);
      end
      IntAluPlugin_AluBitwiseCtrlEnum_XOR_1 : begin
        early0_IntAluPlugin_logic_alu_bitwise = (toplevel_execute_ctrl2_down_early0_SrcPlugin_SRC1_lane0 ^ toplevel_execute_ctrl2_down_early0_SrcPlugin_SRC2_lane0);
      end
      default : begin
        early0_IntAluPlugin_logic_alu_bitwise = 32'h0;
      end
    endcase
  end

  assign early0_IntAluPlugin_logic_alu_result = (_zz_early0_IntAluPlugin_logic_alu_result | _zz_early0_IntAluPlugin_logic_alu_result_2);
  assign toplevel_execute_ctrl2_down_early0_IntAluPlugin_ALU_RESULT_lane0 = early0_IntAluPlugin_logic_alu_result;
  assign early0_IntAluPlugin_logic_wb_valid = toplevel_execute_ctrl2_down_early0_IntAluPlugin_SEL_lane0;
  assign early0_IntAluPlugin_logic_wb_payload = toplevel_execute_ctrl2_down_early0_IntAluPlugin_ALU_RESULT_lane0;
  assign early0_BarrelShifterPlugin_logic_shift_amplitude = _zz_early0_BarrelShifterPlugin_logic_shift_amplitude;
  assign early0_BarrelShifterPlugin_logic_shift_reversed = (toplevel_execute_ctrl2_down_BarrelShifterPlugin_LEFT_lane0 ? _zz_early0_BarrelShifterPlugin_logic_shift_reversed : toplevel_execute_ctrl2_down_early0_SrcPlugin_SRC1_lane0);
  assign early0_BarrelShifterPlugin_logic_shift_shifted = _zz_early0_BarrelShifterPlugin_logic_shift_shifted[31:0];
  assign early0_BarrelShifterPlugin_logic_shift_patched = (toplevel_execute_ctrl2_down_BarrelShifterPlugin_LEFT_lane0 ? _zz_early0_BarrelShifterPlugin_logic_shift_patched : early0_BarrelShifterPlugin_logic_shift_shifted);
  assign toplevel_execute_ctrl2_down_early0_BarrelShifterPlugin_SHIFT_RESULT_lane0 = early0_BarrelShifterPlugin_logic_shift_patched;
  assign early0_BarrelShifterPlugin_logic_wb_valid = toplevel_execute_ctrl3_down_early0_BarrelShifterPlugin_SEL_lane0;
  assign early0_BarrelShifterPlugin_logic_wb_payload = toplevel_execute_ctrl3_down_early0_BarrelShifterPlugin_SHIFT_RESULT_lane0;
  always @(*) begin
    LsuL1_ackUnlock = 1'b0;
    if(LsuPlugin_logic_onCtrl_io_cmdSent) begin
      LsuL1_ackUnlock = 1'b1;
    end
  end

  assign toplevel_execute_ctrl2_down_MUL_SRC1_lane0 = _zz_toplevel_execute_ctrl2_down_MUL_SRC1_lane0;
  assign toplevel_execute_ctrl2_down_MUL_SRC2_lane0 = _zz_toplevel_execute_ctrl2_down_MUL_SRC2_lane0;
  assign toplevel_execute_ctrl3_down_early0_MulPlugin_logic_mul_VALUES_0_lane0 = (toplevel_execute_ctrl3_down_MUL_SRC1_lane0[16 : 0] * toplevel_execute_ctrl3_down_MUL_SRC2_lane0[16 : 0]);
  assign toplevel_execute_ctrl3_down_early0_MulPlugin_logic_mul_VALUES_1_lane0 = _zz_toplevel_execute_ctrl3_down_early0_MulPlugin_logic_mul_VALUES_1_lane0;
  assign toplevel_execute_ctrl3_down_early0_MulPlugin_logic_mul_VALUES_2_lane0 = _zz_toplevel_execute_ctrl3_down_early0_MulPlugin_logic_mul_VALUES_2_lane0;
  assign toplevel_execute_ctrl3_down_early0_MulPlugin_logic_mul_VALUES_3_lane0 = _zz_toplevel_execute_ctrl3_down_early0_MulPlugin_logic_mul_VALUES_3_lane0;
  always @(*) begin
    _zz_toplevel_execute_ctrl3_down_early0_MulPlugin_logic_steps_0_adders_0_lane0 = 61'h0;
    _zz_toplevel_execute_ctrl3_down_early0_MulPlugin_logic_steps_0_adders_0_lane0[33 : 0] = toplevel_execute_ctrl3_down_early0_MulPlugin_logic_mul_VALUES_0_lane0[33 : 0];
    _zz_toplevel_execute_ctrl3_down_early0_MulPlugin_logic_steps_0_adders_0_lane0[60 : 34] = toplevel_execute_ctrl3_down_early0_MulPlugin_logic_mul_VALUES_3_lane0[26 : 0];
  end

  always @(*) begin
    _zz_toplevel_execute_ctrl3_down_early0_MulPlugin_logic_steps_0_adders_0_lane0_1 = 61'h0;
    _zz_toplevel_execute_ctrl3_down_early0_MulPlugin_logic_steps_0_adders_0_lane0_1[60 : 17] = toplevel_execute_ctrl3_down_early0_MulPlugin_logic_mul_VALUES_1_lane0[43 : 0];
  end

  always @(*) begin
    _zz_toplevel_execute_ctrl3_down_early0_MulPlugin_logic_steps_0_adders_0_lane0_2 = 61'h0;
    _zz_toplevel_execute_ctrl3_down_early0_MulPlugin_logic_steps_0_adders_0_lane0_2[60 : 17] = toplevel_execute_ctrl3_down_early0_MulPlugin_logic_mul_VALUES_2_lane0[43 : 0];
  end

  always @(*) begin
    _zz_toplevel_execute_ctrl3_down_early0_MulPlugin_logic_steps_0_adders_1_lane0 = 3'b000;
    _zz_toplevel_execute_ctrl3_down_early0_MulPlugin_logic_steps_0_adders_1_lane0[2 : 0] = toplevel_execute_ctrl3_down_early0_MulPlugin_logic_mul_VALUES_3_lane0[29 : 27];
  end

  always @(*) begin
    _zz_toplevel_execute_ctrl3_down_early0_MulPlugin_logic_steps_0_adders_1_lane0_1 = 3'b000;
    _zz_toplevel_execute_ctrl3_down_early0_MulPlugin_logic_steps_0_adders_1_lane0_1[2 : 0] = toplevel_execute_ctrl3_down_early0_MulPlugin_logic_mul_VALUES_1_lane0[46 : 44];
  end

  always @(*) begin
    _zz_toplevel_execute_ctrl3_down_early0_MulPlugin_logic_steps_0_adders_1_lane0_2 = 3'b000;
    _zz_toplevel_execute_ctrl3_down_early0_MulPlugin_logic_steps_0_adders_1_lane0_2[2 : 0] = toplevel_execute_ctrl3_down_early0_MulPlugin_logic_mul_VALUES_2_lane0[46 : 44];
  end

  assign toplevel_execute_ctrl3_down_early0_MulPlugin_logic_steps_0_adders_0_lane0 = (_zz_toplevel_execute_ctrl3_down_early0_MulPlugin_logic_steps_0_adders_0_lane0_3 + _zz_toplevel_execute_ctrl3_down_early0_MulPlugin_logic_steps_0_adders_0_lane0_6);
  assign toplevel_execute_ctrl3_down_early0_MulPlugin_logic_steps_0_adders_1_lane0 = (_zz_toplevel_execute_ctrl3_down_early0_MulPlugin_logic_steps_0_adders_1_lane0_3 + _zz_toplevel_execute_ctrl3_down_early0_MulPlugin_logic_steps_0_adders_1_lane0_6);
  always @(*) begin
    _zz_toplevel_execute_ctrl4_down_early0_MulPlugin_logic_steps_1_adders_0_lane0 = 66'h0;
    _zz_toplevel_execute_ctrl4_down_early0_MulPlugin_logic_steps_1_adders_0_lane0[62 : 0] = toplevel_execute_ctrl4_down_early0_MulPlugin_logic_steps_0_adders_0_lane0[62 : 0];
  end

  always @(*) begin
    _zz_toplevel_execute_ctrl4_down_early0_MulPlugin_logic_steps_1_adders_0_lane0_1 = 66'h0;
    _zz_toplevel_execute_ctrl4_down_early0_MulPlugin_logic_steps_1_adders_0_lane0_1[65 : 61] = toplevel_execute_ctrl4_down_early0_MulPlugin_logic_steps_0_adders_1_lane0[4 : 0];
  end

  assign toplevel_execute_ctrl4_down_early0_MulPlugin_logic_steps_1_adders_0_lane0 = (_zz_toplevel_execute_ctrl4_down_early0_MulPlugin_logic_steps_1_adders_0_lane0 + _zz_toplevel_execute_ctrl4_down_early0_MulPlugin_logic_steps_1_adders_0_lane0_1);
  assign when_MulPlugin_l195 = ((toplevel_execute_ctrl4_up_LANE_SEL_lane0 && (! toplevel_execute_ctrl4_down_isReady)) && (! toplevel_execute_lane0_ctrls_4_upIsCancel));
  assign early0_MulPlugin_logic_formatBus_valid = toplevel_execute_ctrl4_down_early0_MulPlugin_SEL_lane0;
  assign early0_MulPlugin_logic_formatBus_payload = (toplevel_execute_ctrl4_down_MulPlugin_HIGH_lane0 ? early0_MulPlugin_logic_writeback_buffer_data : toplevel_execute_ctrl4_down_early0_MulPlugin_logic_steps_1_adders_0_lane0[31 : 0]);
  assign toplevel_execute_ctrl2_down_RsUnsignedPlugin_RS1_FORMATED_lane0 = toplevel_execute_ctrl2_up_integer_RS1_lane0;
  assign toplevel_execute_ctrl2_down_RsUnsignedPlugin_RS2_FORMATED_lane0 = toplevel_execute_ctrl2_up_integer_RS2_lane0;
  assign toplevel_execute_ctrl2_down_RsUnsignedPlugin_RS1_REVERT_lane0 = (toplevel_execute_ctrl2_down_RsUnsignedPlugin_RS1_SIGNED_lane0 && toplevel_execute_ctrl2_down_RsUnsignedPlugin_RS1_FORMATED_lane0[31]);
  assign toplevel_execute_ctrl2_down_RsUnsignedPlugin_RS2_REVERT_lane0 = (toplevel_execute_ctrl2_down_RsUnsignedPlugin_RS2_SIGNED_lane0 && toplevel_execute_ctrl2_down_RsUnsignedPlugin_RS2_FORMATED_lane0[31]);
  assign toplevel_execute_ctrl2_down_RsUnsignedPlugin_RS1_UNSIGNED_lane0 = ((toplevel_execute_ctrl2_down_RsUnsignedPlugin_RS1_REVERT_lane0 ? (~ toplevel_execute_ctrl2_down_RsUnsignedPlugin_RS1_FORMATED_lane0) : toplevel_execute_ctrl2_down_RsUnsignedPlugin_RS1_FORMATED_lane0) + _zz_toplevel_execute_ctrl2_down_RsUnsignedPlugin_RS1_UNSIGNED_lane0);
  assign toplevel_execute_ctrl2_down_RsUnsignedPlugin_RS2_UNSIGNED_lane0 = ((toplevel_execute_ctrl2_down_RsUnsignedPlugin_RS2_REVERT_lane0 ? (~ toplevel_execute_ctrl2_down_RsUnsignedPlugin_RS2_FORMATED_lane0) : toplevel_execute_ctrl2_down_RsUnsignedPlugin_RS2_FORMATED_lane0) + _zz_toplevel_execute_ctrl2_down_RsUnsignedPlugin_RS2_UNSIGNED_lane0);
  assign early0_DivPlugin_logic_processing_div_io_cmd_fire = (early0_DivPlugin_logic_processing_div_io_cmd_valid && early0_DivPlugin_logic_processing_div_io_cmd_ready);
  assign early0_DivPlugin_logic_processing_request = (toplevel_execute_ctrl2_up_LANE_SEL_lane0 && toplevel_execute_ctrl2_down_early0_DivPlugin_SEL_lane0);
  assign early0_DivPlugin_logic_processing_a = toplevel_execute_ctrl2_down_RsUnsignedPlugin_RS1_UNSIGNED_lane0;
  assign early0_DivPlugin_logic_processing_b = toplevel_execute_ctrl2_down_RsUnsignedPlugin_RS2_UNSIGNED_lane0;
  always @(*) begin
    early0_DivPlugin_logic_processing_div_io_cmd_valid = (early0_DivPlugin_logic_processing_request && (! early0_DivPlugin_logic_processing_cmdSent));
    if(when_DivPlugin_l118) begin
      early0_DivPlugin_logic_processing_div_io_cmd_valid = 1'b0;
    end
  end

  assign when_DivPlugin_l118 = (! early0_DivPlugin_logic_processing_relaxer_hadRequest);
  assign early0_DivPlugin_logic_processing_freeze = ((early0_DivPlugin_logic_processing_request && (! early0_DivPlugin_logic_processing_div_io_rsp_valid)) && (! early0_DivPlugin_logic_processing_unscheduleRequest));
  assign early0_DivPlugin_logic_processing_selected = (toplevel_execute_ctrl2_down_DivPlugin_REM_lane0 ? early0_DivPlugin_logic_processing_div_io_rsp_payload_remain : early0_DivPlugin_logic_processing_div_io_rsp_payload_result);
  assign _zz_toplevel_execute_ctrl2_down_DivPlugin_DIV_RESULT_lane0 = early0_DivPlugin_logic_processing_selected;
  assign toplevel_execute_ctrl2_down_DivPlugin_DIV_RESULT_lane0 = _zz_toplevel_execute_ctrl2_down_DivPlugin_DIV_RESULT_lane0_1;
  assign early0_DivPlugin_logic_formatBus_valid = toplevel_execute_ctrl3_down_early0_DivPlugin_SEL_lane0;
  assign early0_DivPlugin_logic_formatBus_payload = toplevel_execute_ctrl3_down_DivPlugin_DIV_RESULT_lane0;
  always @(*) begin
    case(toplevel_execute_ctrl4_down_late0_IntAluPlugin_ALU_BITWISE_CTRL_lane0)
      IntAluPlugin_AluBitwiseCtrlEnum_AND_1 : begin
        late0_IntAluPlugin_logic_alu_bitwise = (toplevel_execute_ctrl4_down_late0_SrcPlugin_SRC1_lane0 & toplevel_execute_ctrl4_down_late0_SrcPlugin_SRC2_lane0);
      end
      IntAluPlugin_AluBitwiseCtrlEnum_OR_1 : begin
        late0_IntAluPlugin_logic_alu_bitwise = (toplevel_execute_ctrl4_down_late0_SrcPlugin_SRC1_lane0 | toplevel_execute_ctrl4_down_late0_SrcPlugin_SRC2_lane0);
      end
      IntAluPlugin_AluBitwiseCtrlEnum_XOR_1 : begin
        late0_IntAluPlugin_logic_alu_bitwise = (toplevel_execute_ctrl4_down_late0_SrcPlugin_SRC1_lane0 ^ toplevel_execute_ctrl4_down_late0_SrcPlugin_SRC2_lane0);
      end
      default : begin
        late0_IntAluPlugin_logic_alu_bitwise = 32'h0;
      end
    endcase
  end

  assign late0_IntAluPlugin_logic_alu_result = (_zz_late0_IntAluPlugin_logic_alu_result | _zz_late0_IntAluPlugin_logic_alu_result_2);
  assign toplevel_execute_ctrl4_down_late0_IntAluPlugin_ALU_RESULT_lane0 = late0_IntAluPlugin_logic_alu_result;
  assign late0_IntAluPlugin_logic_wb_valid = toplevel_execute_ctrl4_down_late0_IntAluPlugin_SEL_lane0;
  assign late0_IntAluPlugin_logic_wb_payload = toplevel_execute_ctrl4_down_late0_IntAluPlugin_ALU_RESULT_lane0;
  assign late0_BarrelShifterPlugin_logic_shift_amplitude = _zz_late0_BarrelShifterPlugin_logic_shift_amplitude;
  assign late0_BarrelShifterPlugin_logic_shift_reversed = (toplevel_execute_ctrl4_down_BarrelShifterPlugin_LEFT_lane0 ? _zz_late0_BarrelShifterPlugin_logic_shift_reversed : toplevel_execute_ctrl4_down_late0_SrcPlugin_SRC1_lane0);
  assign late0_BarrelShifterPlugin_logic_shift_shifted = _zz_late0_BarrelShifterPlugin_logic_shift_shifted[31:0];
  assign late0_BarrelShifterPlugin_logic_shift_patched = (toplevel_execute_ctrl4_down_BarrelShifterPlugin_LEFT_lane0 ? _zz_late0_BarrelShifterPlugin_logic_shift_patched : late0_BarrelShifterPlugin_logic_shift_shifted);
  assign toplevel_execute_ctrl4_down_late0_BarrelShifterPlugin_SHIFT_RESULT_lane0 = late0_BarrelShifterPlugin_logic_shift_patched;
  assign late0_BarrelShifterPlugin_logic_wb_valid = toplevel_execute_ctrl4_down_late0_BarrelShifterPlugin_SEL_lane0;
  assign late0_BarrelShifterPlugin_logic_wb_payload = toplevel_execute_ctrl4_down_late0_BarrelShifterPlugin_SHIFT_RESULT_lane0;
  always @(*) begin
    case(toplevel_execute_ctrl2_down_early1_IntAluPlugin_ALU_BITWISE_CTRL_lane1)
      IntAluPlugin_AluBitwiseCtrlEnum_AND_1 : begin
        early1_IntAluPlugin_logic_alu_bitwise = (toplevel_execute_ctrl2_down_early1_SrcPlugin_SRC1_lane1 & toplevel_execute_ctrl2_down_early1_SrcPlugin_SRC2_lane1);
      end
      IntAluPlugin_AluBitwiseCtrlEnum_OR_1 : begin
        early1_IntAluPlugin_logic_alu_bitwise = (toplevel_execute_ctrl2_down_early1_SrcPlugin_SRC1_lane1 | toplevel_execute_ctrl2_down_early1_SrcPlugin_SRC2_lane1);
      end
      IntAluPlugin_AluBitwiseCtrlEnum_XOR_1 : begin
        early1_IntAluPlugin_logic_alu_bitwise = (toplevel_execute_ctrl2_down_early1_SrcPlugin_SRC1_lane1 ^ toplevel_execute_ctrl2_down_early1_SrcPlugin_SRC2_lane1);
      end
      default : begin
        early1_IntAluPlugin_logic_alu_bitwise = 32'h0;
      end
    endcase
  end

  assign early1_IntAluPlugin_logic_alu_result = (_zz_early1_IntAluPlugin_logic_alu_result | _zz_early1_IntAluPlugin_logic_alu_result_2);
  assign toplevel_execute_ctrl2_down_early1_IntAluPlugin_ALU_RESULT_lane1 = early1_IntAluPlugin_logic_alu_result;
  assign early1_IntAluPlugin_logic_wb_valid = toplevel_execute_ctrl2_down_early1_IntAluPlugin_SEL_lane1;
  assign early1_IntAluPlugin_logic_wb_payload = toplevel_execute_ctrl2_down_early1_IntAluPlugin_ALU_RESULT_lane1;
  assign early1_BarrelShifterPlugin_logic_shift_amplitude = _zz_early1_BarrelShifterPlugin_logic_shift_amplitude;
  assign early1_BarrelShifterPlugin_logic_shift_reversed = (toplevel_execute_ctrl2_down_BarrelShifterPlugin_LEFT_lane1 ? _zz_early1_BarrelShifterPlugin_logic_shift_reversed : toplevel_execute_ctrl2_down_early1_SrcPlugin_SRC1_lane1);
  assign early1_BarrelShifterPlugin_logic_shift_shifted = _zz_early1_BarrelShifterPlugin_logic_shift_shifted[31:0];
  assign early1_BarrelShifterPlugin_logic_shift_patched = (toplevel_execute_ctrl2_down_BarrelShifterPlugin_LEFT_lane1 ? _zz_early1_BarrelShifterPlugin_logic_shift_patched : early1_BarrelShifterPlugin_logic_shift_shifted);
  assign toplevel_execute_ctrl2_down_early1_BarrelShifterPlugin_SHIFT_RESULT_lane1 = early1_BarrelShifterPlugin_logic_shift_patched;
  assign early1_BarrelShifterPlugin_logic_wb_valid = toplevel_execute_ctrl3_down_early1_BarrelShifterPlugin_SEL_lane1;
  assign early1_BarrelShifterPlugin_logic_wb_payload = toplevel_execute_ctrl3_down_early1_BarrelShifterPlugin_SHIFT_RESULT_lane1;
  always @(*) begin
    case(toplevel_execute_ctrl4_down_late1_IntAluPlugin_ALU_BITWISE_CTRL_lane1)
      IntAluPlugin_AluBitwiseCtrlEnum_AND_1 : begin
        late1_IntAluPlugin_logic_alu_bitwise = (toplevel_execute_ctrl4_down_late1_SrcPlugin_SRC1_lane1 & toplevel_execute_ctrl4_down_late1_SrcPlugin_SRC2_lane1);
      end
      IntAluPlugin_AluBitwiseCtrlEnum_OR_1 : begin
        late1_IntAluPlugin_logic_alu_bitwise = (toplevel_execute_ctrl4_down_late1_SrcPlugin_SRC1_lane1 | toplevel_execute_ctrl4_down_late1_SrcPlugin_SRC2_lane1);
      end
      IntAluPlugin_AluBitwiseCtrlEnum_XOR_1 : begin
        late1_IntAluPlugin_logic_alu_bitwise = (toplevel_execute_ctrl4_down_late1_SrcPlugin_SRC1_lane1 ^ toplevel_execute_ctrl4_down_late1_SrcPlugin_SRC2_lane1);
      end
      default : begin
        late1_IntAluPlugin_logic_alu_bitwise = 32'h0;
      end
    endcase
  end

  assign late1_IntAluPlugin_logic_alu_result = (_zz_late1_IntAluPlugin_logic_alu_result | _zz_late1_IntAluPlugin_logic_alu_result_2);
  assign toplevel_execute_ctrl4_down_late1_IntAluPlugin_ALU_RESULT_lane1 = late1_IntAluPlugin_logic_alu_result;
  assign late1_IntAluPlugin_logic_wb_valid = toplevel_execute_ctrl4_down_late1_IntAluPlugin_SEL_lane1;
  assign late1_IntAluPlugin_logic_wb_payload = toplevel_execute_ctrl4_down_late1_IntAluPlugin_ALU_RESULT_lane1;
  assign late1_BarrelShifterPlugin_logic_shift_amplitude = _zz_late1_BarrelShifterPlugin_logic_shift_amplitude;
  assign late1_BarrelShifterPlugin_logic_shift_reversed = (toplevel_execute_ctrl4_down_BarrelShifterPlugin_LEFT_lane1 ? _zz_late1_BarrelShifterPlugin_logic_shift_reversed : toplevel_execute_ctrl4_down_late1_SrcPlugin_SRC1_lane1);
  assign late1_BarrelShifterPlugin_logic_shift_shifted = _zz_late1_BarrelShifterPlugin_logic_shift_shifted[31:0];
  assign late1_BarrelShifterPlugin_logic_shift_patched = (toplevel_execute_ctrl4_down_BarrelShifterPlugin_LEFT_lane1 ? _zz_late1_BarrelShifterPlugin_logic_shift_patched : late1_BarrelShifterPlugin_logic_shift_shifted);
  assign toplevel_execute_ctrl4_down_late1_BarrelShifterPlugin_SHIFT_RESULT_lane1 = late1_BarrelShifterPlugin_logic_shift_patched;
  assign late1_BarrelShifterPlugin_logic_wb_valid = toplevel_execute_ctrl4_down_late1_BarrelShifterPlugin_SEL_lane1;
  assign late1_BarrelShifterPlugin_logic_wb_payload = toplevel_execute_ctrl4_down_late1_BarrelShifterPlugin_SHIFT_RESULT_lane1;
  assign WhiteboxerPlugin_logic_fetch_fire = fetch_logic_ctrls_0_down_isFiring;
  assign PrivilegedPlugin_api_harts_0_allowInterrupts = 1'b1;
  assign PrivilegedPlugin_api_harts_0_allowException = 1'b1;
  assign PrivilegedPlugin_api_harts_0_allowEbreakException = 1'b1;
  assign PrivilegedPlugin_api_harts_0_fpuEnable = 1'b0;
  always @(*) begin
    case(toplevel_execute_ctrl2_down_BranchPlugin_BRANCH_CTRL_lane0)
      BranchPlugin_BranchCtrlEnum_JALR : begin
        early0_BranchPlugin_pcCalc_target_a = toplevel_execute_ctrl2_down_early0_SrcPlugin_SRC1_lane0;
      end
      default : begin
        early0_BranchPlugin_pcCalc_target_a = toplevel_execute_ctrl2_down_PC_lane0;
      end
    endcase
  end

  always @(*) begin
    case(toplevel_execute_ctrl2_down_BranchPlugin_BRANCH_CTRL_lane0)
      BranchPlugin_BranchCtrlEnum_JAL : begin
        early0_BranchPlugin_pcCalc_target_b = {{11{_zz_early0_BranchPlugin_pcCalc_target_b[20]}}, _zz_early0_BranchPlugin_pcCalc_target_b};
      end
      BranchPlugin_BranchCtrlEnum_JALR : begin
        early0_BranchPlugin_pcCalc_target_b = {{20{_zz_early0_BranchPlugin_pcCalc_target_b_1[11]}}, _zz_early0_BranchPlugin_pcCalc_target_b_1};
      end
      default : begin
        early0_BranchPlugin_pcCalc_target_b = {{19{_zz_early0_BranchPlugin_pcCalc_target_b_2[12]}}, _zz_early0_BranchPlugin_pcCalc_target_b_2};
      end
    endcase
  end

  assign early0_BranchPlugin_pcCalc_slices = ({1'b0,toplevel_execute_ctrl2_down_Decode_INSTRUCTION_SLICE_COUNT_lane0} + {1'b0,1'b1});
  always @(*) begin
    toplevel_execute_ctrl2_down_early0_BranchPlugin_pcCalc_PC_TRUE_lane0 = _zz_toplevel_execute_ctrl2_down_early0_BranchPlugin_pcCalc_PC_TRUE_lane0;
    toplevel_execute_ctrl2_down_early0_BranchPlugin_pcCalc_PC_TRUE_lane0[0] = 1'b0;
  end

  assign toplevel_execute_ctrl2_down_early0_BranchPlugin_pcCalc_PC_FALSE_lane0 = (toplevel_execute_ctrl2_down_PC_lane0 + _zz_toplevel_execute_ctrl2_down_early0_BranchPlugin_pcCalc_PC_FALSE_lane0);
  assign toplevel_execute_ctrl2_down_early0_BranchPlugin_pcCalc_PC_LAST_SLICE_lane0 = (toplevel_execute_ctrl2_down_PC_lane0 + _zz_toplevel_execute_ctrl2_down_early0_BranchPlugin_pcCalc_PC_LAST_SLICE_lane0);
  always @(*) begin
    case(toplevel_execute_ctrl2_down_BranchPlugin_BRANCH_CTRL_lane1)
      BranchPlugin_BranchCtrlEnum_JALR : begin
        early1_BranchPlugin_pcCalc_target_a = toplevel_execute_ctrl2_down_early1_SrcPlugin_SRC1_lane1;
      end
      default : begin
        early1_BranchPlugin_pcCalc_target_a = toplevel_execute_ctrl2_down_PC_lane1;
      end
    endcase
  end

  always @(*) begin
    case(toplevel_execute_ctrl2_down_BranchPlugin_BRANCH_CTRL_lane1)
      BranchPlugin_BranchCtrlEnum_JAL : begin
        early1_BranchPlugin_pcCalc_target_b = {{11{_zz_early1_BranchPlugin_pcCalc_target_b[20]}}, _zz_early1_BranchPlugin_pcCalc_target_b};
      end
      BranchPlugin_BranchCtrlEnum_JALR : begin
        early1_BranchPlugin_pcCalc_target_b = {{20{_zz_early1_BranchPlugin_pcCalc_target_b_1[11]}}, _zz_early1_BranchPlugin_pcCalc_target_b_1};
      end
      default : begin
        early1_BranchPlugin_pcCalc_target_b = {{19{_zz_early1_BranchPlugin_pcCalc_target_b_2[12]}}, _zz_early1_BranchPlugin_pcCalc_target_b_2};
      end
    endcase
  end

  assign early1_BranchPlugin_pcCalc_slices = ({1'b0,toplevel_execute_ctrl2_down_Decode_INSTRUCTION_SLICE_COUNT_lane1} + {1'b0,1'b1});
  always @(*) begin
    toplevel_execute_ctrl2_down_early1_BranchPlugin_pcCalc_PC_TRUE_lane1 = _zz_toplevel_execute_ctrl2_down_early1_BranchPlugin_pcCalc_PC_TRUE_lane1;
    toplevel_execute_ctrl2_down_early1_BranchPlugin_pcCalc_PC_TRUE_lane1[0] = 1'b0;
  end

  assign toplevel_execute_ctrl2_down_early1_BranchPlugin_pcCalc_PC_FALSE_lane1 = (toplevel_execute_ctrl2_down_PC_lane1 + _zz_toplevel_execute_ctrl2_down_early1_BranchPlugin_pcCalc_PC_FALSE_lane1);
  assign toplevel_execute_ctrl2_down_early1_BranchPlugin_pcCalc_PC_LAST_SLICE_lane1 = (toplevel_execute_ctrl2_down_PC_lane1 + _zz_toplevel_execute_ctrl2_down_early1_BranchPlugin_pcCalc_PC_LAST_SLICE_lane1);
  assign AlignerPlugin_logic_maskGen_frontMasks_0 = 4'b1111;
  assign AlignerPlugin_logic_maskGen_frontMasks_1 = 4'b1110;
  assign AlignerPlugin_logic_maskGen_frontMasks_2 = 4'b1100;
  assign AlignerPlugin_logic_maskGen_frontMasks_3 = 4'b1000;
  assign AlignerPlugin_logic_maskGen_backMasks_0 = 4'b0001;
  assign AlignerPlugin_logic_maskGen_backMasks_1 = 4'b0011;
  assign AlignerPlugin_logic_maskGen_backMasks_2 = 4'b0111;
  assign AlignerPlugin_logic_maskGen_backMasks_3 = 4'b1111;
  assign fetch_logic_ctrls_2_down_AlignerPlugin_logic_FETCH_MASK = (_zz_fetch_logic_ctrls_2_down_AlignerPlugin_logic_FETCH_MASK & ((! fetch_logic_ctrls_2_down_Prediction_WORD_JUMPED) ? 4'b1111 : _zz_fetch_logic_ctrls_2_down_AlignerPlugin_logic_FETCH_MASK_2));
  assign fetch_logic_ctrls_2_down_AlignerPlugin_logic_FETCH_LAST = ((fetch_logic_ctrls_2_up_isValid && fetch_logic_ctrls_2_down_Prediction_WORD_JUMPED) ? _zz_fetch_logic_ctrls_2_down_AlignerPlugin_logic_FETCH_LAST : 4'b0000);
  assign AlignerPlugin_logic_slicesInstructions_0 = {AlignerPlugin_logic_slices_data_1,AlignerPlugin_logic_slices_data_0};
  assign AlignerPlugin_logic_slicesInstructions_1 = {AlignerPlugin_logic_slices_data_2,AlignerPlugin_logic_slices_data_1};
  assign AlignerPlugin_logic_slicesInstructions_2 = {AlignerPlugin_logic_slices_data_3,AlignerPlugin_logic_slices_data_2};
  assign AlignerPlugin_logic_slicesInstructions_3 = {AlignerPlugin_logic_slices_data_4,AlignerPlugin_logic_slices_data_3};
  assign AlignerPlugin_logic_slicesInstructions_4 = {AlignerPlugin_logic_slices_data_5,AlignerPlugin_logic_slices_data_4};
  assign AlignerPlugin_logic_slicesInstructions_5 = {AlignerPlugin_logic_slices_data_6,AlignerPlugin_logic_slices_data_5};
  assign AlignerPlugin_logic_slicesInstructions_6 = {AlignerPlugin_logic_slices_data_7,AlignerPlugin_logic_slices_data_6};
  assign AlignerPlugin_logic_slicesInstructions_7 = {16'd0, AlignerPlugin_logic_slices_data_7};
  always @(*) begin
    AlignerPlugin_logic_scanners_0_usageMask = 8'h0;
    AlignerPlugin_logic_scanners_0_usageMask[0] = AlignerPlugin_logic_scanners_0_checker_0_required;
    AlignerPlugin_logic_scanners_0_usageMask[1] = AlignerPlugin_logic_scanners_0_checker_1_required;
  end

  assign AlignerPlugin_logic_scanners_0_checker_0_required = 1'b1;
  assign AlignerPlugin_logic_scanners_0_checker_0_last = (AlignerPlugin_logic_slices_data_0[1 : 0] != 2'b11);
  assign AlignerPlugin_logic_scanners_0_checker_0_redo = ((AlignerPlugin_logic_scanners_0_checker_0_required && AlignerPlugin_logic_slices_last[0]) && (! AlignerPlugin_logic_scanners_0_checker_0_last));
  assign AlignerPlugin_logic_scanners_0_checker_0_present = AlignerPlugin_logic_slices_mask[0];
  assign AlignerPlugin_logic_scanners_0_checker_0_valid = AlignerPlugin_logic_scanners_0_checker_0_present;
  assign AlignerPlugin_logic_scanners_0_checker_1_required = (AlignerPlugin_logic_slices_data_0[1 : 0] == 2'b11);
  assign AlignerPlugin_logic_scanners_0_checker_1_last = (AlignerPlugin_logic_slices_data_0[1 : 0] == 2'b11);
  assign AlignerPlugin_logic_scanners_0_checker_1_redo = ((AlignerPlugin_logic_scanners_0_checker_1_required && AlignerPlugin_logic_slices_last[1]) && (! AlignerPlugin_logic_scanners_0_checker_1_last));
  assign AlignerPlugin_logic_scanners_0_checker_1_present = AlignerPlugin_logic_slices_mask[1];
  assign AlignerPlugin_logic_scanners_0_checker_1_valid = (AlignerPlugin_logic_scanners_0_checker_1_present || (! AlignerPlugin_logic_scanners_0_checker_1_required));
  assign AlignerPlugin_logic_scanners_0_redo = (|{AlignerPlugin_logic_scanners_0_checker_1_redo,AlignerPlugin_logic_scanners_0_checker_0_redo});
  assign AlignerPlugin_logic_scanners_0_valid = (AlignerPlugin_logic_scanners_0_checker_0_valid && ((&AlignerPlugin_logic_scanners_0_checker_1_valid) || (|{AlignerPlugin_logic_scanners_0_checker_1_redo,AlignerPlugin_logic_scanners_0_checker_0_redo})));
  always @(*) begin
    AlignerPlugin_logic_scanners_1_usageMask = 8'h0;
    AlignerPlugin_logic_scanners_1_usageMask[1] = AlignerPlugin_logic_scanners_1_checker_0_required;
    AlignerPlugin_logic_scanners_1_usageMask[2] = AlignerPlugin_logic_scanners_1_checker_1_required;
  end

  assign AlignerPlugin_logic_scanners_1_checker_0_required = 1'b1;
  assign AlignerPlugin_logic_scanners_1_checker_0_last = (AlignerPlugin_logic_slices_data_1[1 : 0] != 2'b11);
  assign AlignerPlugin_logic_scanners_1_checker_0_redo = ((AlignerPlugin_logic_scanners_1_checker_0_required && AlignerPlugin_logic_slices_last[1]) && (! AlignerPlugin_logic_scanners_1_checker_0_last));
  assign AlignerPlugin_logic_scanners_1_checker_0_present = AlignerPlugin_logic_slices_mask[1];
  assign AlignerPlugin_logic_scanners_1_checker_0_valid = AlignerPlugin_logic_scanners_1_checker_0_present;
  assign AlignerPlugin_logic_scanners_1_checker_1_required = (AlignerPlugin_logic_slices_data_1[1 : 0] == 2'b11);
  assign AlignerPlugin_logic_scanners_1_checker_1_last = (AlignerPlugin_logic_slices_data_1[1 : 0] == 2'b11);
  assign AlignerPlugin_logic_scanners_1_checker_1_redo = ((AlignerPlugin_logic_scanners_1_checker_1_required && AlignerPlugin_logic_slices_last[2]) && (! AlignerPlugin_logic_scanners_1_checker_1_last));
  assign AlignerPlugin_logic_scanners_1_checker_1_present = AlignerPlugin_logic_slices_mask[2];
  assign AlignerPlugin_logic_scanners_1_checker_1_valid = (AlignerPlugin_logic_scanners_1_checker_1_present || (! AlignerPlugin_logic_scanners_1_checker_1_required));
  assign AlignerPlugin_logic_scanners_1_redo = (|{AlignerPlugin_logic_scanners_1_checker_1_redo,AlignerPlugin_logic_scanners_1_checker_0_redo});
  assign AlignerPlugin_logic_scanners_1_valid = (AlignerPlugin_logic_scanners_1_checker_0_valid && ((&AlignerPlugin_logic_scanners_1_checker_1_valid) || (|{AlignerPlugin_logic_scanners_1_checker_1_redo,AlignerPlugin_logic_scanners_1_checker_0_redo})));
  always @(*) begin
    AlignerPlugin_logic_scanners_2_usageMask = 8'h0;
    AlignerPlugin_logic_scanners_2_usageMask[2] = AlignerPlugin_logic_scanners_2_checker_0_required;
    AlignerPlugin_logic_scanners_2_usageMask[3] = AlignerPlugin_logic_scanners_2_checker_1_required;
  end

  assign AlignerPlugin_logic_scanners_2_checker_0_required = 1'b1;
  assign AlignerPlugin_logic_scanners_2_checker_0_last = (AlignerPlugin_logic_slices_data_2[1 : 0] != 2'b11);
  assign AlignerPlugin_logic_scanners_2_checker_0_redo = ((AlignerPlugin_logic_scanners_2_checker_0_required && AlignerPlugin_logic_slices_last[2]) && (! AlignerPlugin_logic_scanners_2_checker_0_last));
  assign AlignerPlugin_logic_scanners_2_checker_0_present = AlignerPlugin_logic_slices_mask[2];
  assign AlignerPlugin_logic_scanners_2_checker_0_valid = AlignerPlugin_logic_scanners_2_checker_0_present;
  assign AlignerPlugin_logic_scanners_2_checker_1_required = (AlignerPlugin_logic_slices_data_2[1 : 0] == 2'b11);
  assign AlignerPlugin_logic_scanners_2_checker_1_last = (AlignerPlugin_logic_slices_data_2[1 : 0] == 2'b11);
  assign AlignerPlugin_logic_scanners_2_checker_1_redo = ((AlignerPlugin_logic_scanners_2_checker_1_required && AlignerPlugin_logic_slices_last[3]) && (! AlignerPlugin_logic_scanners_2_checker_1_last));
  assign AlignerPlugin_logic_scanners_2_checker_1_present = AlignerPlugin_logic_slices_mask[3];
  assign AlignerPlugin_logic_scanners_2_checker_1_valid = (AlignerPlugin_logic_scanners_2_checker_1_present || (! AlignerPlugin_logic_scanners_2_checker_1_required));
  assign AlignerPlugin_logic_scanners_2_redo = (|{AlignerPlugin_logic_scanners_2_checker_1_redo,AlignerPlugin_logic_scanners_2_checker_0_redo});
  assign AlignerPlugin_logic_scanners_2_valid = (AlignerPlugin_logic_scanners_2_checker_0_valid && ((&AlignerPlugin_logic_scanners_2_checker_1_valid) || (|{AlignerPlugin_logic_scanners_2_checker_1_redo,AlignerPlugin_logic_scanners_2_checker_0_redo})));
  always @(*) begin
    AlignerPlugin_logic_scanners_3_usageMask = 8'h0;
    AlignerPlugin_logic_scanners_3_usageMask[3] = AlignerPlugin_logic_scanners_3_checker_0_required;
    AlignerPlugin_logic_scanners_3_usageMask[4] = AlignerPlugin_logic_scanners_3_checker_1_required;
  end

  assign AlignerPlugin_logic_scanners_3_checker_0_required = 1'b1;
  assign AlignerPlugin_logic_scanners_3_checker_0_last = (AlignerPlugin_logic_slices_data_3[1 : 0] != 2'b11);
  assign AlignerPlugin_logic_scanners_3_checker_0_redo = ((AlignerPlugin_logic_scanners_3_checker_0_required && AlignerPlugin_logic_slices_last[3]) && (! AlignerPlugin_logic_scanners_3_checker_0_last));
  assign AlignerPlugin_logic_scanners_3_checker_0_present = AlignerPlugin_logic_slices_mask[3];
  assign AlignerPlugin_logic_scanners_3_checker_0_valid = AlignerPlugin_logic_scanners_3_checker_0_present;
  assign AlignerPlugin_logic_scanners_3_checker_1_required = (AlignerPlugin_logic_slices_data_3[1 : 0] == 2'b11);
  assign AlignerPlugin_logic_scanners_3_checker_1_last = (AlignerPlugin_logic_slices_data_3[1 : 0] == 2'b11);
  assign AlignerPlugin_logic_scanners_3_checker_1_redo = ((AlignerPlugin_logic_scanners_3_checker_1_required && AlignerPlugin_logic_slices_last[4]) && (! AlignerPlugin_logic_scanners_3_checker_1_last));
  assign AlignerPlugin_logic_scanners_3_checker_1_present = AlignerPlugin_logic_slices_mask[4];
  assign AlignerPlugin_logic_scanners_3_checker_1_valid = (AlignerPlugin_logic_scanners_3_checker_1_present || (! AlignerPlugin_logic_scanners_3_checker_1_required));
  assign AlignerPlugin_logic_scanners_3_redo = (|{AlignerPlugin_logic_scanners_3_checker_1_redo,AlignerPlugin_logic_scanners_3_checker_0_redo});
  assign AlignerPlugin_logic_scanners_3_valid = (AlignerPlugin_logic_scanners_3_checker_0_valid && ((&AlignerPlugin_logic_scanners_3_checker_1_valid) || (|{AlignerPlugin_logic_scanners_3_checker_1_redo,AlignerPlugin_logic_scanners_3_checker_0_redo})));
  always @(*) begin
    AlignerPlugin_logic_scanners_4_usageMask = 8'h0;
    AlignerPlugin_logic_scanners_4_usageMask[4] = AlignerPlugin_logic_scanners_4_checker_0_required;
    AlignerPlugin_logic_scanners_4_usageMask[5] = AlignerPlugin_logic_scanners_4_checker_1_required;
  end

  assign AlignerPlugin_logic_scanners_4_checker_0_required = 1'b1;
  assign AlignerPlugin_logic_scanners_4_checker_0_last = (AlignerPlugin_logic_slices_data_4[1 : 0] != 2'b11);
  assign AlignerPlugin_logic_scanners_4_checker_0_redo = ((AlignerPlugin_logic_scanners_4_checker_0_required && AlignerPlugin_logic_slices_last[4]) && (! AlignerPlugin_logic_scanners_4_checker_0_last));
  assign AlignerPlugin_logic_scanners_4_checker_0_present = AlignerPlugin_logic_slices_mask[4];
  assign AlignerPlugin_logic_scanners_4_checker_0_valid = AlignerPlugin_logic_scanners_4_checker_0_present;
  assign AlignerPlugin_logic_scanners_4_checker_1_required = (AlignerPlugin_logic_slices_data_4[1 : 0] == 2'b11);
  assign AlignerPlugin_logic_scanners_4_checker_1_last = (AlignerPlugin_logic_slices_data_4[1 : 0] == 2'b11);
  assign AlignerPlugin_logic_scanners_4_checker_1_redo = ((AlignerPlugin_logic_scanners_4_checker_1_required && AlignerPlugin_logic_slices_last[5]) && (! AlignerPlugin_logic_scanners_4_checker_1_last));
  assign AlignerPlugin_logic_scanners_4_checker_1_present = AlignerPlugin_logic_slices_mask[5];
  assign AlignerPlugin_logic_scanners_4_checker_1_valid = (AlignerPlugin_logic_scanners_4_checker_1_present || (! AlignerPlugin_logic_scanners_4_checker_1_required));
  assign AlignerPlugin_logic_scanners_4_redo = (|{AlignerPlugin_logic_scanners_4_checker_1_redo,AlignerPlugin_logic_scanners_4_checker_0_redo});
  assign AlignerPlugin_logic_scanners_4_valid = (AlignerPlugin_logic_scanners_4_checker_0_valid && ((&AlignerPlugin_logic_scanners_4_checker_1_valid) || (|{AlignerPlugin_logic_scanners_4_checker_1_redo,AlignerPlugin_logic_scanners_4_checker_0_redo})));
  always @(*) begin
    AlignerPlugin_logic_scanners_5_usageMask = 8'h0;
    AlignerPlugin_logic_scanners_5_usageMask[5] = AlignerPlugin_logic_scanners_5_checker_0_required;
    AlignerPlugin_logic_scanners_5_usageMask[6] = AlignerPlugin_logic_scanners_5_checker_1_required;
  end

  assign AlignerPlugin_logic_scanners_5_checker_0_required = 1'b1;
  assign AlignerPlugin_logic_scanners_5_checker_0_last = (AlignerPlugin_logic_slices_data_5[1 : 0] != 2'b11);
  assign AlignerPlugin_logic_scanners_5_checker_0_redo = ((AlignerPlugin_logic_scanners_5_checker_0_required && AlignerPlugin_logic_slices_last[5]) && (! AlignerPlugin_logic_scanners_5_checker_0_last));
  assign AlignerPlugin_logic_scanners_5_checker_0_present = AlignerPlugin_logic_slices_mask[5];
  assign AlignerPlugin_logic_scanners_5_checker_0_valid = AlignerPlugin_logic_scanners_5_checker_0_present;
  assign AlignerPlugin_logic_scanners_5_checker_1_required = (AlignerPlugin_logic_slices_data_5[1 : 0] == 2'b11);
  assign AlignerPlugin_logic_scanners_5_checker_1_last = (AlignerPlugin_logic_slices_data_5[1 : 0] == 2'b11);
  assign AlignerPlugin_logic_scanners_5_checker_1_redo = ((AlignerPlugin_logic_scanners_5_checker_1_required && AlignerPlugin_logic_slices_last[6]) && (! AlignerPlugin_logic_scanners_5_checker_1_last));
  assign AlignerPlugin_logic_scanners_5_checker_1_present = AlignerPlugin_logic_slices_mask[6];
  assign AlignerPlugin_logic_scanners_5_checker_1_valid = (AlignerPlugin_logic_scanners_5_checker_1_present || (! AlignerPlugin_logic_scanners_5_checker_1_required));
  assign AlignerPlugin_logic_scanners_5_redo = (|{AlignerPlugin_logic_scanners_5_checker_1_redo,AlignerPlugin_logic_scanners_5_checker_0_redo});
  assign AlignerPlugin_logic_scanners_5_valid = (AlignerPlugin_logic_scanners_5_checker_0_valid && ((&AlignerPlugin_logic_scanners_5_checker_1_valid) || (|{AlignerPlugin_logic_scanners_5_checker_1_redo,AlignerPlugin_logic_scanners_5_checker_0_redo})));
  always @(*) begin
    AlignerPlugin_logic_scanners_6_usageMask = 8'h0;
    AlignerPlugin_logic_scanners_6_usageMask[6] = AlignerPlugin_logic_scanners_6_checker_0_required;
    AlignerPlugin_logic_scanners_6_usageMask[7] = AlignerPlugin_logic_scanners_6_checker_1_required;
  end

  assign AlignerPlugin_logic_scanners_6_checker_0_required = 1'b1;
  assign AlignerPlugin_logic_scanners_6_checker_0_last = (AlignerPlugin_logic_slices_data_6[1 : 0] != 2'b11);
  assign AlignerPlugin_logic_scanners_6_checker_0_redo = ((AlignerPlugin_logic_scanners_6_checker_0_required && AlignerPlugin_logic_slices_last[6]) && (! AlignerPlugin_logic_scanners_6_checker_0_last));
  assign AlignerPlugin_logic_scanners_6_checker_0_present = AlignerPlugin_logic_slices_mask[6];
  assign AlignerPlugin_logic_scanners_6_checker_0_valid = AlignerPlugin_logic_scanners_6_checker_0_present;
  assign AlignerPlugin_logic_scanners_6_checker_1_required = (AlignerPlugin_logic_slices_data_6[1 : 0] == 2'b11);
  assign AlignerPlugin_logic_scanners_6_checker_1_last = (AlignerPlugin_logic_slices_data_6[1 : 0] == 2'b11);
  assign AlignerPlugin_logic_scanners_6_checker_1_redo = ((AlignerPlugin_logic_scanners_6_checker_1_required && AlignerPlugin_logic_slices_last[7]) && (! AlignerPlugin_logic_scanners_6_checker_1_last));
  assign AlignerPlugin_logic_scanners_6_checker_1_present = AlignerPlugin_logic_slices_mask[7];
  assign AlignerPlugin_logic_scanners_6_checker_1_valid = (AlignerPlugin_logic_scanners_6_checker_1_present || (! AlignerPlugin_logic_scanners_6_checker_1_required));
  assign AlignerPlugin_logic_scanners_6_redo = (|{AlignerPlugin_logic_scanners_6_checker_1_redo,AlignerPlugin_logic_scanners_6_checker_0_redo});
  assign AlignerPlugin_logic_scanners_6_valid = (AlignerPlugin_logic_scanners_6_checker_0_valid && ((&AlignerPlugin_logic_scanners_6_checker_1_valid) || (|{AlignerPlugin_logic_scanners_6_checker_1_redo,AlignerPlugin_logic_scanners_6_checker_0_redo})));
  always @(*) begin
    AlignerPlugin_logic_scanners_7_usageMask = 8'h0;
    AlignerPlugin_logic_scanners_7_usageMask[7] = AlignerPlugin_logic_scanners_7_checker_0_required;
  end

  assign AlignerPlugin_logic_scanners_7_checker_0_required = 1'b1;
  assign AlignerPlugin_logic_scanners_7_checker_0_last = (AlignerPlugin_logic_slices_data_7[1 : 0] != 2'b11);
  assign AlignerPlugin_logic_scanners_7_checker_0_redo = ((AlignerPlugin_logic_scanners_7_checker_0_required && AlignerPlugin_logic_slices_last[7]) && (! AlignerPlugin_logic_scanners_7_checker_0_last));
  assign AlignerPlugin_logic_scanners_7_checker_0_present = AlignerPlugin_logic_slices_mask[7];
  assign AlignerPlugin_logic_scanners_7_checker_0_valid = AlignerPlugin_logic_scanners_7_checker_0_present;
  assign AlignerPlugin_logic_scanners_7_checker_1_required = (AlignerPlugin_logic_slices_data_7[1 : 0] == 2'b11);
  assign AlignerPlugin_logic_scanners_7_checker_1_last = (AlignerPlugin_logic_slices_data_7[1 : 0] == 2'b11);
  assign AlignerPlugin_logic_scanners_7_checker_1_redo = 1'b0;
  assign AlignerPlugin_logic_scanners_7_checker_1_present = 1'b0;
  assign AlignerPlugin_logic_scanners_7_checker_1_valid = (AlignerPlugin_logic_scanners_7_checker_1_present || (! AlignerPlugin_logic_scanners_7_checker_1_required));
  assign AlignerPlugin_logic_scanners_7_redo = (|{AlignerPlugin_logic_scanners_7_checker_1_redo,AlignerPlugin_logic_scanners_7_checker_0_redo});
  assign AlignerPlugin_logic_scanners_7_valid = (AlignerPlugin_logic_scanners_7_checker_0_valid && ((&AlignerPlugin_logic_scanners_7_checker_1_valid) || (|{AlignerPlugin_logic_scanners_7_checker_1_redo,AlignerPlugin_logic_scanners_7_checker_0_redo})));
  assign AlignerPlugin_logic_usedMask_0 = 8'h0;
  assign AlignerPlugin_logic_extractors_0_first = 1'b1;
  assign AlignerPlugin_logic_extractors_0_usableMask = {(AlignerPlugin_logic_scanners_7_valid && (! AlignerPlugin_logic_usedMask_0[7])),{(AlignerPlugin_logic_scanners_6_valid && (! AlignerPlugin_logic_usedMask_0[6])),{(AlignerPlugin_logic_scanners_5_valid && (! AlignerPlugin_logic_usedMask_0[5])),{(AlignerPlugin_logic_scanners_4_valid && (! _zz_AlignerPlugin_logic_extractors_0_usableMask)),{(AlignerPlugin_logic_scanners_3_valid && _zz_AlignerPlugin_logic_extractors_0_usableMask_1),{_zz_AlignerPlugin_logic_extractors_0_usableMask_2,{_zz_AlignerPlugin_logic_extractors_0_usableMask_3,_zz_AlignerPlugin_logic_extractors_0_usableMask_4}}}}}}};
  assign _zz_AlignerPlugin_logic_extractors_0_usableMask_bools_0 = AlignerPlugin_logic_extractors_0_usableMask;
  assign AlignerPlugin_logic_extractors_0_usableMask_bools_0 = _zz_AlignerPlugin_logic_extractors_0_usableMask_bools_0[0];
  assign AlignerPlugin_logic_extractors_0_usableMask_bools_1 = _zz_AlignerPlugin_logic_extractors_0_usableMask_bools_0[1];
  assign AlignerPlugin_logic_extractors_0_usableMask_bools_2 = _zz_AlignerPlugin_logic_extractors_0_usableMask_bools_0[2];
  assign AlignerPlugin_logic_extractors_0_usableMask_bools_3 = _zz_AlignerPlugin_logic_extractors_0_usableMask_bools_0[3];
  assign AlignerPlugin_logic_extractors_0_usableMask_bools_4 = _zz_AlignerPlugin_logic_extractors_0_usableMask_bools_0[4];
  assign AlignerPlugin_logic_extractors_0_usableMask_bools_5 = _zz_AlignerPlugin_logic_extractors_0_usableMask_bools_0[5];
  assign AlignerPlugin_logic_extractors_0_usableMask_bools_6 = _zz_AlignerPlugin_logic_extractors_0_usableMask_bools_0[6];
  assign AlignerPlugin_logic_extractors_0_usableMask_bools_7 = _zz_AlignerPlugin_logic_extractors_0_usableMask_bools_0[7];
  always @(*) begin
    _zz_AlignerPlugin_logic_extractors_0_slicesOh[0] = (AlignerPlugin_logic_extractors_0_usableMask_bools_0 && (! 1'b0));
    _zz_AlignerPlugin_logic_extractors_0_slicesOh[1] = (AlignerPlugin_logic_extractors_0_usableMask_bools_1 && (! AlignerPlugin_logic_extractors_0_usableMask_bools_0));
    _zz_AlignerPlugin_logic_extractors_0_slicesOh[2] = (AlignerPlugin_logic_extractors_0_usableMask_bools_2 && (! AlignerPlugin_logic_extractors_0_usableMask_range_0_to_1));
    _zz_AlignerPlugin_logic_extractors_0_slicesOh[3] = (AlignerPlugin_logic_extractors_0_usableMask_bools_3 && (! AlignerPlugin_logic_extractors_0_usableMask_range_0_to_2));
    _zz_AlignerPlugin_logic_extractors_0_slicesOh[4] = (AlignerPlugin_logic_extractors_0_usableMask_bools_4 && (! AlignerPlugin_logic_extractors_0_usableMask_range_0_to_3));
    _zz_AlignerPlugin_logic_extractors_0_slicesOh[5] = (AlignerPlugin_logic_extractors_0_usableMask_bools_5 && (! (AlignerPlugin_logic_extractors_0_usableMask_bools_4 || AlignerPlugin_logic_extractors_0_usableMask_range_0_to_3)));
    _zz_AlignerPlugin_logic_extractors_0_slicesOh[6] = (AlignerPlugin_logic_extractors_0_usableMask_bools_6 && (! (AlignerPlugin_logic_extractors_0_usableMask_range_4_to_5 || AlignerPlugin_logic_extractors_0_usableMask_range_0_to_3)));
    _zz_AlignerPlugin_logic_extractors_0_slicesOh[7] = (AlignerPlugin_logic_extractors_0_usableMask_bools_7 && (! (AlignerPlugin_logic_extractors_0_usableMask_range_4_to_6 || AlignerPlugin_logic_extractors_0_usableMask_range_0_to_3)));
  end

  assign AlignerPlugin_logic_extractors_0_usableMask_range_0_to_1 = (|{AlignerPlugin_logic_extractors_0_usableMask_bools_1,AlignerPlugin_logic_extractors_0_usableMask_bools_0});
  assign AlignerPlugin_logic_extractors_0_usableMask_range_0_to_2 = (|{AlignerPlugin_logic_extractors_0_usableMask_bools_2,{AlignerPlugin_logic_extractors_0_usableMask_bools_1,AlignerPlugin_logic_extractors_0_usableMask_bools_0}});
  assign AlignerPlugin_logic_extractors_0_usableMask_range_0_to_3 = (|{AlignerPlugin_logic_extractors_0_usableMask_bools_3,{AlignerPlugin_logic_extractors_0_usableMask_bools_2,{AlignerPlugin_logic_extractors_0_usableMask_bools_1,AlignerPlugin_logic_extractors_0_usableMask_bools_0}}});
  assign AlignerPlugin_logic_extractors_0_usableMask_range_4_to_5 = (|{AlignerPlugin_logic_extractors_0_usableMask_bools_5,AlignerPlugin_logic_extractors_0_usableMask_bools_4});
  assign AlignerPlugin_logic_extractors_0_usableMask_range_4_to_6 = (|{AlignerPlugin_logic_extractors_0_usableMask_bools_6,{AlignerPlugin_logic_extractors_0_usableMask_bools_5,AlignerPlugin_logic_extractors_0_usableMask_bools_4}});
  assign AlignerPlugin_logic_extractors_0_slicesOh = _zz_AlignerPlugin_logic_extractors_0_slicesOh;
  assign _zz_AlignerPlugin_logic_extractors_0_redo = AlignerPlugin_logic_extractors_0_slicesOh[0];
  assign _zz_AlignerPlugin_logic_extractors_0_redo_1 = AlignerPlugin_logic_extractors_0_slicesOh[1];
  assign _zz_AlignerPlugin_logic_extractors_0_redo_2 = AlignerPlugin_logic_extractors_0_slicesOh[2];
  assign _zz_AlignerPlugin_logic_extractors_0_redo_3 = AlignerPlugin_logic_extractors_0_slicesOh[3];
  assign _zz_AlignerPlugin_logic_extractors_0_redo_4 = AlignerPlugin_logic_extractors_0_slicesOh[4];
  assign _zz_AlignerPlugin_logic_extractors_0_redo_5 = AlignerPlugin_logic_extractors_0_slicesOh[5];
  assign _zz_AlignerPlugin_logic_extractors_0_redo_6 = AlignerPlugin_logic_extractors_0_slicesOh[6];
  assign _zz_AlignerPlugin_logic_extractors_0_redo_7 = AlignerPlugin_logic_extractors_0_slicesOh[7];
  always @(*) begin
    AlignerPlugin_logic_extractors_0_redo = _zz_AlignerPlugin_logic_extractors_0_redo_8[0];
    if(when_AlignerPlugin_l163) begin
      AlignerPlugin_logic_extractors_0_redo = 1'b0;
    end
  end

  assign AlignerPlugin_logic_extractors_0_localMask = ((((_zz_AlignerPlugin_logic_extractors_0_redo ? {_zz_AlignerPlugin_logic_extractors_0_localMask,_zz_AlignerPlugin_logic_extractors_0_localMask_1} : 2'b00) | (_zz_AlignerPlugin_logic_extractors_0_redo_1 ? {_zz_AlignerPlugin_logic_extractors_0_localMask_2,_zz_AlignerPlugin_logic_extractors_0_localMask_3} : 2'b00)) | ((_zz_AlignerPlugin_logic_extractors_0_redo_2 ? {_zz_AlignerPlugin_logic_extractors_0_localMask_4,_zz_AlignerPlugin_logic_extractors_0_localMask_5} : 2'b00) | (_zz_AlignerPlugin_logic_extractors_0_redo_3 ? {_zz_AlignerPlugin_logic_extractors_0_localMask_6,_zz_AlignerPlugin_logic_extractors_0_localMask_7} : 2'b00))) | (((_zz_AlignerPlugin_logic_extractors_0_redo_4 ? {_zz_AlignerPlugin_logic_extractors_0_localMask_8,_zz_AlignerPlugin_logic_extractors_0_localMask_9} : 2'b00) | (_zz_AlignerPlugin_logic_extractors_0_redo_5 ? {_zz_AlignerPlugin_logic_extractors_0_localMask_10,_zz_AlignerPlugin_logic_extractors_0_localMask_11} : 2'b00)) | ((_zz_AlignerPlugin_logic_extractors_0_redo_6 ? {_zz_AlignerPlugin_logic_extractors_0_localMask_12,_zz_AlignerPlugin_logic_extractors_0_localMask_13} : 2'b00) | (_zz_AlignerPlugin_logic_extractors_0_redo_7 ? {_zz_AlignerPlugin_logic_extractors_0_localMask_14,_zz_AlignerPlugin_logic_extractors_0_localMask_15} : 2'b00))));
  assign AlignerPlugin_logic_extractors_0_usageMask = ((((_zz_AlignerPlugin_logic_extractors_0_redo ? AlignerPlugin_logic_scanners_0_usageMask : 8'h0) | (_zz_AlignerPlugin_logic_extractors_0_redo_1 ? AlignerPlugin_logic_scanners_1_usageMask : 8'h0)) | ((_zz_AlignerPlugin_logic_extractors_0_redo_2 ? AlignerPlugin_logic_scanners_2_usageMask : 8'h0) | (_zz_AlignerPlugin_logic_extractors_0_redo_3 ? AlignerPlugin_logic_scanners_3_usageMask : 8'h0))) | (((_zz_AlignerPlugin_logic_extractors_0_redo_4 ? AlignerPlugin_logic_scanners_4_usageMask : 8'h0) | (_zz_AlignerPlugin_logic_extractors_0_redo_5 ? AlignerPlugin_logic_scanners_5_usageMask : 8'h0)) | ((_zz_AlignerPlugin_logic_extractors_0_redo_6 ? AlignerPlugin_logic_scanners_6_usageMask : 8'h0) | (_zz_AlignerPlugin_logic_extractors_0_redo_7 ? AlignerPlugin_logic_scanners_7_usageMask : 8'h0))));
  assign AlignerPlugin_logic_usedMask_1 = (AlignerPlugin_logic_usedMask_0 | AlignerPlugin_logic_extractors_0_usageMask);
  always @(*) begin
    AlignerPlugin_logic_extractors_0_valid = (|AlignerPlugin_logic_extractors_0_slicesOh);
    if(when_AlignerPlugin_l163) begin
      AlignerPlugin_logic_extractors_0_valid = 1'b0;
    end
    if(when_AlignerPlugin_l243) begin
      if(when_AlignerPlugin_l244) begin
        AlignerPlugin_logic_extractors_0_valid = 1'b0;
      end
    end
  end

  assign when_AlignerPlugin_l163 = (AlignerPlugin_api_haltIt || (AlignerPlugin_api_singleFetch && (! AlignerPlugin_logic_extractors_0_first)));
  assign AlignerPlugin_logic_extractors_1_first = 1'b0;
  assign AlignerPlugin_logic_extractors_1_usableMask = {(AlignerPlugin_logic_scanners_7_valid && (! AlignerPlugin_logic_usedMask_1[7])),{(AlignerPlugin_logic_scanners_6_valid && (! AlignerPlugin_logic_usedMask_1[6])),{(AlignerPlugin_logic_scanners_5_valid && (! AlignerPlugin_logic_usedMask_1[5])),{(AlignerPlugin_logic_scanners_4_valid && (! _zz_AlignerPlugin_logic_extractors_1_usableMask)),{(AlignerPlugin_logic_scanners_3_valid && _zz_AlignerPlugin_logic_extractors_1_usableMask_1),{_zz_AlignerPlugin_logic_extractors_1_usableMask_2,_zz_AlignerPlugin_logic_extractors_1_usableMask_3}}}}}};
  assign _zz_AlignerPlugin_logic_extractors_1_usableMask_bools_0 = AlignerPlugin_logic_extractors_1_usableMask;
  assign AlignerPlugin_logic_extractors_1_usableMask_bools_0 = _zz_AlignerPlugin_logic_extractors_1_usableMask_bools_0[0];
  assign AlignerPlugin_logic_extractors_1_usableMask_bools_1 = _zz_AlignerPlugin_logic_extractors_1_usableMask_bools_0[1];
  assign AlignerPlugin_logic_extractors_1_usableMask_bools_2 = _zz_AlignerPlugin_logic_extractors_1_usableMask_bools_0[2];
  assign AlignerPlugin_logic_extractors_1_usableMask_bools_3 = _zz_AlignerPlugin_logic_extractors_1_usableMask_bools_0[3];
  assign AlignerPlugin_logic_extractors_1_usableMask_bools_4 = _zz_AlignerPlugin_logic_extractors_1_usableMask_bools_0[4];
  assign AlignerPlugin_logic_extractors_1_usableMask_bools_5 = _zz_AlignerPlugin_logic_extractors_1_usableMask_bools_0[5];
  assign AlignerPlugin_logic_extractors_1_usableMask_bools_6 = _zz_AlignerPlugin_logic_extractors_1_usableMask_bools_0[6];
  always @(*) begin
    _zz_AlignerPlugin_logic_extractors_1_slicesOh[0] = (AlignerPlugin_logic_extractors_1_usableMask_bools_0 && (! 1'b0));
    _zz_AlignerPlugin_logic_extractors_1_slicesOh[1] = (AlignerPlugin_logic_extractors_1_usableMask_bools_1 && (! AlignerPlugin_logic_extractors_1_usableMask_bools_0));
    _zz_AlignerPlugin_logic_extractors_1_slicesOh[2] = (AlignerPlugin_logic_extractors_1_usableMask_bools_2 && (! AlignerPlugin_logic_extractors_1_usableMask_range_0_to_1));
    _zz_AlignerPlugin_logic_extractors_1_slicesOh[3] = (AlignerPlugin_logic_extractors_1_usableMask_bools_3 && (! AlignerPlugin_logic_extractors_1_usableMask_range_0_to_2));
    _zz_AlignerPlugin_logic_extractors_1_slicesOh[4] = (AlignerPlugin_logic_extractors_1_usableMask_bools_4 && (! AlignerPlugin_logic_extractors_1_usableMask_range_0_to_3));
    _zz_AlignerPlugin_logic_extractors_1_slicesOh[5] = (AlignerPlugin_logic_extractors_1_usableMask_bools_5 && (! (AlignerPlugin_logic_extractors_1_usableMask_bools_4 || AlignerPlugin_logic_extractors_1_usableMask_range_0_to_3)));
    _zz_AlignerPlugin_logic_extractors_1_slicesOh[6] = (AlignerPlugin_logic_extractors_1_usableMask_bools_6 && (! (AlignerPlugin_logic_extractors_1_usableMask_range_4_to_5 || AlignerPlugin_logic_extractors_1_usableMask_range_0_to_3)));
  end

  assign AlignerPlugin_logic_extractors_1_usableMask_range_0_to_1 = (|{AlignerPlugin_logic_extractors_1_usableMask_bools_1,AlignerPlugin_logic_extractors_1_usableMask_bools_0});
  assign AlignerPlugin_logic_extractors_1_usableMask_range_0_to_2 = (|{AlignerPlugin_logic_extractors_1_usableMask_bools_2,{AlignerPlugin_logic_extractors_1_usableMask_bools_1,AlignerPlugin_logic_extractors_1_usableMask_bools_0}});
  assign AlignerPlugin_logic_extractors_1_usableMask_range_0_to_3 = (|{AlignerPlugin_logic_extractors_1_usableMask_bools_3,{AlignerPlugin_logic_extractors_1_usableMask_bools_2,{AlignerPlugin_logic_extractors_1_usableMask_bools_1,AlignerPlugin_logic_extractors_1_usableMask_bools_0}}});
  assign AlignerPlugin_logic_extractors_1_usableMask_range_4_to_5 = (|{AlignerPlugin_logic_extractors_1_usableMask_bools_5,AlignerPlugin_logic_extractors_1_usableMask_bools_4});
  assign AlignerPlugin_logic_extractors_1_slicesOh = _zz_AlignerPlugin_logic_extractors_1_slicesOh;
  assign _zz_AlignerPlugin_logic_extractors_1_redo = AlignerPlugin_logic_extractors_1_slicesOh[0];
  assign _zz_AlignerPlugin_logic_extractors_1_redo_1 = AlignerPlugin_logic_extractors_1_slicesOh[1];
  assign _zz_AlignerPlugin_logic_extractors_1_redo_2 = AlignerPlugin_logic_extractors_1_slicesOh[2];
  assign _zz_AlignerPlugin_logic_extractors_1_redo_3 = AlignerPlugin_logic_extractors_1_slicesOh[3];
  assign _zz_AlignerPlugin_logic_extractors_1_redo_4 = AlignerPlugin_logic_extractors_1_slicesOh[4];
  assign _zz_AlignerPlugin_logic_extractors_1_redo_5 = AlignerPlugin_logic_extractors_1_slicesOh[5];
  assign _zz_AlignerPlugin_logic_extractors_1_redo_6 = AlignerPlugin_logic_extractors_1_slicesOh[6];
  always @(*) begin
    AlignerPlugin_logic_extractors_1_redo = _zz_AlignerPlugin_logic_extractors_1_redo_7[0];
    if(when_AlignerPlugin_l163_1) begin
      AlignerPlugin_logic_extractors_1_redo = 1'b0;
    end
  end

  assign AlignerPlugin_logic_extractors_1_localMask = ((((_zz_AlignerPlugin_logic_extractors_1_redo ? {_zz_AlignerPlugin_logic_extractors_1_localMask,_zz_AlignerPlugin_logic_extractors_1_localMask_1} : 2'b00) | (_zz_AlignerPlugin_logic_extractors_1_redo_1 ? {_zz_AlignerPlugin_logic_extractors_1_localMask_2,_zz_AlignerPlugin_logic_extractors_1_localMask_3} : 2'b00)) | ((_zz_AlignerPlugin_logic_extractors_1_redo_2 ? {_zz_AlignerPlugin_logic_extractors_1_localMask_4,_zz_AlignerPlugin_logic_extractors_1_localMask_5} : 2'b00) | (_zz_AlignerPlugin_logic_extractors_1_redo_3 ? {_zz_AlignerPlugin_logic_extractors_1_localMask_6,_zz_AlignerPlugin_logic_extractors_1_localMask_7} : 2'b00))) | (((_zz_AlignerPlugin_logic_extractors_1_redo_4 ? {_zz_AlignerPlugin_logic_extractors_1_localMask_8,_zz_AlignerPlugin_logic_extractors_1_localMask_9} : 2'b00) | (_zz_AlignerPlugin_logic_extractors_1_redo_5 ? {_zz_AlignerPlugin_logic_extractors_1_localMask_10,_zz_AlignerPlugin_logic_extractors_1_localMask_11} : 2'b00)) | (_zz_AlignerPlugin_logic_extractors_1_redo_6 ? {AlignerPlugin_logic_scanners_7_checker_1_required,AlignerPlugin_logic_scanners_7_checker_0_required} : 2'b00)));
  assign AlignerPlugin_logic_extractors_1_usageMask = ((((_zz_AlignerPlugin_logic_extractors_1_redo ? AlignerPlugin_logic_scanners_1_usageMask : 8'h0) | (_zz_AlignerPlugin_logic_extractors_1_redo_1 ? AlignerPlugin_logic_scanners_2_usageMask : 8'h0)) | ((_zz_AlignerPlugin_logic_extractors_1_redo_2 ? AlignerPlugin_logic_scanners_3_usageMask : 8'h0) | (_zz_AlignerPlugin_logic_extractors_1_redo_3 ? AlignerPlugin_logic_scanners_4_usageMask : 8'h0))) | (((_zz_AlignerPlugin_logic_extractors_1_redo_4 ? AlignerPlugin_logic_scanners_5_usageMask : 8'h0) | (_zz_AlignerPlugin_logic_extractors_1_redo_5 ? AlignerPlugin_logic_scanners_6_usageMask : 8'h0)) | (_zz_AlignerPlugin_logic_extractors_1_redo_6 ? AlignerPlugin_logic_scanners_7_usageMask : 8'h0)));
  assign AlignerPlugin_logic_usedMask_2 = (AlignerPlugin_logic_usedMask_1 | AlignerPlugin_logic_extractors_1_usageMask);
  always @(*) begin
    AlignerPlugin_logic_extractors_1_valid = (|AlignerPlugin_logic_extractors_1_slicesOh);
    if(when_AlignerPlugin_l163_1) begin
      AlignerPlugin_logic_extractors_1_valid = 1'b0;
    end
    if(when_AlignerPlugin_l243) begin
      if(when_AlignerPlugin_l244_1) begin
        AlignerPlugin_logic_extractors_1_valid = 1'b0;
      end
    end
  end

  assign when_AlignerPlugin_l163_1 = (AlignerPlugin_api_haltIt || (AlignerPlugin_api_singleFetch && (! AlignerPlugin_logic_extractors_1_first)));
  assign when_AlignerPlugin_l173 = (toplevel_decode_ctrls_0_up_isFiring && 1'b1);
  assign AlignerPlugin_logic_feeder_lanes_0_valid = AlignerPlugin_logic_extractors_0_valid;
  assign toplevel_decode_ctrls_0_up_LANE_SEL_0 = AlignerPlugin_logic_feeder_lanes_0_valid;
  always @(*) begin
    toplevel_decode_ctrls_0_up_Decode_INSTRUCTION_0 = AlignerPlugin_logic_extractors_0_ctx_instruction;
    if(AlignerPlugin_logic_feeder_lanes_0_isRvc) begin
      toplevel_decode_ctrls_0_up_Decode_INSTRUCTION_0 = AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst;
    end
  end

  always @(*) begin
    toplevel_decode_ctrls_0_up_Decode_DECOMPRESSION_FAULT_0 = 1'b0;
    if(AlignerPlugin_logic_feeder_lanes_0_isRvc) begin
      toplevel_decode_ctrls_0_up_Decode_DECOMPRESSION_FAULT_0 = AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_illegal;
    end
  end

  always @(*) begin
    toplevel_decode_ctrls_0_up_Decode_INSTRUCTION_RAW_0 = AlignerPlugin_logic_extractors_0_ctx_instruction;
    if(AlignerPlugin_logic_feeder_lanes_0_isRvc) begin
      toplevel_decode_ctrls_0_up_Decode_INSTRUCTION_RAW_0[31 : 16] = 16'h0;
    end
  end

  assign AlignerPlugin_logic_feeder_lanes_0_isRvc = (AlignerPlugin_logic_extractors_0_ctx_instruction[1 : 0] != 2'b11);
  always @(*) begin
    AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst = 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
    case(switch_Rvc_l52)
      5'h0 : begin
        AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst = {{{{{{{{{2'b00,AlignerPlugin_logic_extractors_0_ctx_instruction[10 : 7]},AlignerPlugin_logic_extractors_0_ctx_instruction[12 : 11]},AlignerPlugin_logic_extractors_0_ctx_instruction[5]},AlignerPlugin_logic_extractors_0_ctx_instruction[6]},2'b00},5'h02},3'b000},_zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_1},7'h13};
      end
      5'h02 : begin
        AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst = {{{{_zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_2,_zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst},3'b010},_zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_1},7'h03};
      end
      5'h05 : begin
        AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst = {{{{{_zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_3[11 : 5],_zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_1},_zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst},3'b011},_zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_3[4 : 0]},7'h27};
      end
      5'h06 : begin
        AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst = {{{{{_zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_2[11 : 5],_zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_1},_zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst},3'b010},_zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_2[4 : 0]},7'h23};
      end
      5'h08 : begin
        AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst = {{{{_zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_5,AlignerPlugin_logic_extractors_0_ctx_instruction[11 : 7]},3'b000},AlignerPlugin_logic_extractors_0_ctx_instruction[11 : 7]},7'h13};
      end
      5'h09 : begin
        AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst = {{{{{_zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_8[20],_zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_8[10 : 1]},_zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_8[11]},_zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_8[19 : 12]},_zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_20},7'h6f};
      end
      5'h0a : begin
        AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst = {{{{_zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_5,5'h0},3'b000},AlignerPlugin_logic_extractors_0_ctx_instruction[11 : 7]},7'h13};
      end
      5'h0b : begin
        AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst = ((AlignerPlugin_logic_extractors_0_ctx_instruction[11 : 7] == 5'h02) ? {{{{{{{{_zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_23,_zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_24},_zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_25},AlignerPlugin_logic_extractors_0_ctx_instruction[6]},4'b0000},AlignerPlugin_logic_extractors_0_ctx_instruction[11 : 7]},3'b000},AlignerPlugin_logic_extractors_0_ctx_instruction[11 : 7]},7'h13} : {{_zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_26[31 : 12],AlignerPlugin_logic_extractors_0_ctx_instruction[11 : 7]},7'h37});
      end
      5'h0c : begin
        AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst = _zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_27;
      end
      5'h0d : begin
        AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst = {{{{{_zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_15[20],_zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_15[10 : 1]},_zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_15[11]},_zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_15[19 : 12]},_zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_19},7'h6f};
      end
      5'h0e : begin
        AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst = {{{{{{{_zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_18[12],_zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_18[10 : 5]},_zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_19},_zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst},3'b000},_zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_18[4 : 1]},_zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_18[11]},7'h63};
      end
      5'h0f : begin
        AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst = {{{{{{{_zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_18[12],_zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_18[10 : 5]},_zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_19},_zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst},3'b001},_zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_18[4 : 1]},_zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_18[11]},7'h63};
      end
      5'h10 : begin
        AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst = {{{{{{6'h0,AlignerPlugin_logic_extractors_0_ctx_instruction[12]},AlignerPlugin_logic_extractors_0_ctx_instruction[6 : 2]},AlignerPlugin_logic_extractors_0_ctx_instruction[11 : 7]},3'b001},AlignerPlugin_logic_extractors_0_ctx_instruction[11 : 7]},7'h13};
      end
      5'h12 : begin
        AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst = {{{{{{{{4'b0000,AlignerPlugin_logic_extractors_0_ctx_instruction[3 : 2]},AlignerPlugin_logic_extractors_0_ctx_instruction[12]},AlignerPlugin_logic_extractors_0_ctx_instruction[6 : 4]},2'b00},_zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_21},3'b010},AlignerPlugin_logic_extractors_0_ctx_instruction[11 : 7]},7'h03};
      end
      5'h14 : begin
        AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst = ((AlignerPlugin_logic_extractors_0_ctx_instruction[12 : 2] == 11'h400) ? 32'h00100073 : ((AlignerPlugin_logic_extractors_0_ctx_instruction[6 : 2] == 5'h0) ? {{{{12'h0,AlignerPlugin_logic_extractors_0_ctx_instruction[11 : 7]},3'b000},(AlignerPlugin_logic_extractors_0_ctx_instruction[12] ? _zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_20 : _zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_19)},7'h67} : {{{{{_zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_31,_zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_32},(_zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_33 ? _zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_34 : _zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_19)},3'b000},AlignerPlugin_logic_extractors_0_ctx_instruction[11 : 7]},7'h33}));
      end
      5'h16 : begin
        AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst = {{{{{_zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_35[11 : 5],AlignerPlugin_logic_extractors_0_ctx_instruction[6 : 2]},_zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_21},3'b010},_zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_36[4 : 0]},7'h23};
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_illegal = 1'b0;
    case(switch_Rvc_l52)
      5'h0 : begin
        if(when_Rvc_l56) begin
          AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_illegal = 1'b1;
        end
      end
      5'h02 : begin
      end
      5'h05 : begin
      end
      5'h06 : begin
      end
      5'h08 : begin
      end
      5'h09 : begin
      end
      5'h0a : begin
      end
      5'h0b : begin
        if(when_Rvc_l77) begin
          AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_illegal = 1'b1;
        end
      end
      5'h0c : begin
      end
      5'h0d : begin
      end
      5'h0e : begin
      end
      5'h0f : begin
      end
      5'h10 : begin
      end
      5'h12 : begin
        if(when_Rvc_l98) begin
          AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_illegal = 1'b1;
        end
      end
      5'h14 : begin
        if(when_Rvc_l111) begin
          AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_illegal = 1'b1;
        end
      end
      5'h16 : begin
      end
      default : begin
        AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_illegal = 1'b1;
      end
    endcase
  end

  assign _zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst = {2'b01,AlignerPlugin_logic_extractors_0_ctx_instruction[9 : 7]};
  assign _zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_1 = {2'b01,AlignerPlugin_logic_extractors_0_ctx_instruction[4 : 2]};
  assign _zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_2 = {{{{5'h0,AlignerPlugin_logic_extractors_0_ctx_instruction[5]},AlignerPlugin_logic_extractors_0_ctx_instruction[12 : 10]},AlignerPlugin_logic_extractors_0_ctx_instruction[6]},2'b00};
  assign _zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_3 = {{{4'b0000,AlignerPlugin_logic_extractors_0_ctx_instruction[6 : 5]},AlignerPlugin_logic_extractors_0_ctx_instruction[12 : 10]},3'b000};
  assign _zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_4 = AlignerPlugin_logic_extractors_0_ctx_instruction[12];
  always @(*) begin
    _zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_5[11] = _zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_4;
    _zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_5[10] = _zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_4;
    _zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_5[9] = _zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_4;
    _zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_5[8] = _zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_4;
    _zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_5[7] = _zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_4;
    _zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_5[6] = _zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_4;
    _zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_5[5] = _zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_4;
    _zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_5[4 : 0] = AlignerPlugin_logic_extractors_0_ctx_instruction[6 : 2];
  end

  assign _zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_6 = AlignerPlugin_logic_extractors_0_ctx_instruction[12];
  always @(*) begin
    _zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_7[9] = _zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_6;
    _zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_7[8] = _zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_6;
    _zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_7[7] = _zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_6;
    _zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_7[6] = _zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_6;
    _zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_7[5] = _zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_6;
    _zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_7[4] = _zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_6;
    _zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_7[3] = _zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_6;
    _zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_7[2] = _zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_6;
    _zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_7[1] = _zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_6;
    _zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_7[0] = _zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_6;
  end

  assign _zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_8 = {{{{{{{{_zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_7,AlignerPlugin_logic_extractors_0_ctx_instruction[8]},AlignerPlugin_logic_extractors_0_ctx_instruction[10 : 9]},AlignerPlugin_logic_extractors_0_ctx_instruction[6]},AlignerPlugin_logic_extractors_0_ctx_instruction[7]},AlignerPlugin_logic_extractors_0_ctx_instruction[2]},AlignerPlugin_logic_extractors_0_ctx_instruction[11]},AlignerPlugin_logic_extractors_0_ctx_instruction[5 : 3]},1'b0};
  assign _zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_9 = AlignerPlugin_logic_extractors_0_ctx_instruction[12];
  always @(*) begin
    _zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_10[14] = _zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_9;
    _zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_10[13] = _zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_9;
    _zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_10[12] = _zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_9;
    _zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_10[11] = _zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_9;
    _zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_10[10] = _zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_9;
    _zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_10[9] = _zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_9;
    _zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_10[8] = _zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_9;
    _zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_10[7] = _zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_9;
    _zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_10[6] = _zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_9;
    _zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_10[5] = _zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_9;
    _zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_10[4] = _zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_9;
    _zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_10[3] = _zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_9;
    _zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_10[2] = _zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_9;
    _zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_10[1] = _zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_9;
    _zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_10[0] = _zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_9;
  end

  assign _zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_11 = AlignerPlugin_logic_extractors_0_ctx_instruction[12];
  always @(*) begin
    _zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_12[2] = _zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_11;
    _zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_12[1] = _zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_11;
    _zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_12[0] = _zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_11;
  end

  assign _zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_13 = AlignerPlugin_logic_extractors_0_ctx_instruction[12];
  always @(*) begin
    _zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_14[9] = _zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_13;
    _zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_14[8] = _zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_13;
    _zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_14[7] = _zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_13;
    _zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_14[6] = _zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_13;
    _zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_14[5] = _zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_13;
    _zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_14[4] = _zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_13;
    _zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_14[3] = _zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_13;
    _zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_14[2] = _zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_13;
    _zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_14[1] = _zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_13;
    _zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_14[0] = _zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_13;
  end

  assign _zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_15 = {{{{{{{{_zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_14,AlignerPlugin_logic_extractors_0_ctx_instruction[8]},AlignerPlugin_logic_extractors_0_ctx_instruction[10 : 9]},AlignerPlugin_logic_extractors_0_ctx_instruction[6]},AlignerPlugin_logic_extractors_0_ctx_instruction[7]},AlignerPlugin_logic_extractors_0_ctx_instruction[2]},AlignerPlugin_logic_extractors_0_ctx_instruction[11]},AlignerPlugin_logic_extractors_0_ctx_instruction[5 : 3]},1'b0};
  assign _zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_16 = AlignerPlugin_logic_extractors_0_ctx_instruction[12];
  always @(*) begin
    _zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_17[4] = _zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_16;
    _zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_17[3] = _zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_16;
    _zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_17[2] = _zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_16;
    _zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_17[1] = _zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_16;
    _zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_17[0] = _zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_16;
  end

  assign _zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_18 = {{{{{_zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_17,AlignerPlugin_logic_extractors_0_ctx_instruction[6 : 5]},AlignerPlugin_logic_extractors_0_ctx_instruction[2]},AlignerPlugin_logic_extractors_0_ctx_instruction[11 : 10]},AlignerPlugin_logic_extractors_0_ctx_instruction[4 : 3]},1'b0};
  assign _zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_19 = 5'h0;
  assign _zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_20 = 5'h01;
  assign _zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_21 = 5'h02;
  assign switch_Rvc_l52 = {AlignerPlugin_logic_extractors_0_ctx_instruction[1 : 0],AlignerPlugin_logic_extractors_0_ctx_instruction[15 : 13]};
  assign when_Rvc_l56 = (AlignerPlugin_logic_extractors_0_ctx_instruction[12 : 5] == 8'h0);
  assign when_Rvc_l77 = ((AlignerPlugin_logic_extractors_0_ctx_instruction[6 : 2] == 5'h0) && (AlignerPlugin_logic_extractors_0_ctx_instruction[12] == 1'b0));
  assign _zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_22 = {{{{_zz__zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst_22,_zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst},3'b101},_zz_AlignerPlugin_logic_feeder_lanes_0_withRvc_dec_inst},7'h13};
  assign when_Rvc_l98 = (AlignerPlugin_logic_extractors_0_ctx_instruction[11 : 7] == 5'h0);
  assign when_Rvc_l111 = (((AlignerPlugin_logic_extractors_0_ctx_instruction[11 : 7] == 5'h0) && (AlignerPlugin_logic_extractors_0_ctx_instruction[6 : 2] == 5'h0)) && (AlignerPlugin_logic_extractors_0_ctx_instruction[12] == 1'b0));
  assign _zz_toplevel_decode_ctrls_0_up_Decode_INSTRUCTION_SLICE_COUNT_0 = AlignerPlugin_logic_extractors_0_localMask;
  assign _zz_toplevel_decode_ctrls_0_up_Decode_INSTRUCTION_SLICE_COUNT_0_1 = {_zz_toplevel_decode_ctrls_0_up_Decode_INSTRUCTION_SLICE_COUNT_0[0],_zz_toplevel_decode_ctrls_0_up_Decode_INSTRUCTION_SLICE_COUNT_0[1]};
  assign _zz_toplevel_decode_ctrls_0_up_Decode_INSTRUCTION_SLICE_COUNT_0_2 = _zz_toplevel_decode_ctrls_0_up_Decode_INSTRUCTION_SLICE_COUNT_0_1[0];
  always @(*) begin
    _zz_toplevel_decode_ctrls_0_up_Decode_INSTRUCTION_SLICE_COUNT_0_3[0] = (_zz_toplevel_decode_ctrls_0_up_Decode_INSTRUCTION_SLICE_COUNT_0_2 && (! 1'b0));
    _zz_toplevel_decode_ctrls_0_up_Decode_INSTRUCTION_SLICE_COUNT_0_3[1] = (_zz_toplevel_decode_ctrls_0_up_Decode_INSTRUCTION_SLICE_COUNT_0_1[1] && (! _zz_toplevel_decode_ctrls_0_up_Decode_INSTRUCTION_SLICE_COUNT_0_2));
  end

  assign _zz_toplevel_decode_ctrls_0_up_Decode_INSTRUCTION_SLICE_COUNT_0_4 = _zz_toplevel_decode_ctrls_0_up_Decode_INSTRUCTION_SLICE_COUNT_0_3;
  assign _zz_toplevel_decode_ctrls_0_up_Decode_INSTRUCTION_SLICE_COUNT_0_5 = _zz__zz_toplevel_decode_ctrls_0_up_Decode_INSTRUCTION_SLICE_COUNT_0_5[1];
  assign toplevel_decode_ctrls_0_up_Decode_INSTRUCTION_SLICE_COUNT_0 = _zz_toplevel_decode_ctrls_0_up_Decode_INSTRUCTION_SLICE_COUNT_0_5;
  assign toplevel_decode_ctrls_0_up_PC_0 = AlignerPlugin_logic_extractors_0_ctx_pc;
  assign toplevel_decode_ctrls_0_up_Decode_DOP_ID_0 = AlignerPlugin_logic_feeder_harts_0_dopId;
  assign toplevel_decode_ctrls_0_up_Fetch_ID_0 = AlignerPlugin_logic_extractors_0_ctx_hm_Fetch_ID;
  assign toplevel_decode_ctrls_0_up_GSharePlugin_GSHARE_COUNTER_0_0 = AlignerPlugin_logic_extractors_0_ctx_hm_GSharePlugin_GSHARE_COUNTER_0;
  assign toplevel_decode_ctrls_0_up_GSharePlugin_GSHARE_COUNTER_0_1 = AlignerPlugin_logic_extractors_0_ctx_hm_GSharePlugin_GSHARE_COUNTER_1;
  assign toplevel_decode_ctrls_0_up_GSharePlugin_GSHARE_COUNTER_0_2 = AlignerPlugin_logic_extractors_0_ctx_hm_GSharePlugin_GSHARE_COUNTER_2;
  assign toplevel_decode_ctrls_0_up_GSharePlugin_GSHARE_COUNTER_0_3 = AlignerPlugin_logic_extractors_0_ctx_hm_GSharePlugin_GSHARE_COUNTER_3;
  assign toplevel_decode_ctrls_0_up_Prediction_BRANCH_HISTORY_0 = AlignerPlugin_logic_extractors_0_ctx_hm_Prediction_BRANCH_HISTORY;
  assign toplevel_decode_ctrls_0_up_Prediction_WORD_SLICES_BRANCH_0 = AlignerPlugin_logic_extractors_0_ctx_hm_Prediction_WORD_SLICES_BRANCH;
  assign toplevel_decode_ctrls_0_up_Prediction_WORD_SLICES_TAKEN_0 = AlignerPlugin_logic_extractors_0_ctx_hm_Prediction_WORD_SLICES_TAKEN;
  assign toplevel_decode_ctrls_0_up_Prediction_WORD_JUMP_PC_0 = AlignerPlugin_logic_extractors_0_ctx_hm_Prediction_WORD_JUMP_PC;
  assign toplevel_decode_ctrls_0_up_Prediction_WORD_JUMPED_0 = AlignerPlugin_logic_extractors_0_ctx_hm_Prediction_WORD_JUMPED;
  assign toplevel_decode_ctrls_0_up_Prediction_WORD_JUMP_SLICE_0 = AlignerPlugin_logic_extractors_0_ctx_hm_Prediction_WORD_JUMP_SLICE;
  assign toplevel_decode_ctrls_0_up_TRAP_0 = AlignerPlugin_logic_extractors_0_ctx_trap;
  assign AlignerPlugin_logic_feeder_lanes_0_onBtb_pcLastSlice = (toplevel_decode_ctrls_0_up_PC_0[2 : 1] + _zz_AlignerPlugin_logic_feeder_lanes_0_onBtb_pcLastSlice);
  assign AlignerPlugin_logic_feeder_lanes_0_onBtb_didPrediction = (toplevel_decode_ctrls_0_up_Prediction_WORD_JUMP_SLICE_0 <= AlignerPlugin_logic_feeder_lanes_0_onBtb_pcLastSlice);
  assign toplevel_decode_ctrls_0_up_Prediction_ALIGNED_JUMPED_0 = (toplevel_decode_ctrls_0_up_Prediction_WORD_JUMPED_0 && AlignerPlugin_logic_feeder_lanes_0_onBtb_didPrediction);
  assign toplevel_decode_ctrls_0_up_Prediction_ALIGNED_JUMPED_PC_0 = toplevel_decode_ctrls_0_up_Prediction_WORD_JUMP_PC_0;
  assign toplevel_decode_ctrls_0_up_Prediction_ALIGNED_SLICES_BRANCH_0 = toplevel_decode_ctrls_0_up_Prediction_WORD_SLICES_BRANCH_0;
  assign toplevel_decode_ctrls_0_up_Prediction_ALIGNED_SLICES_TAKEN_0 = toplevel_decode_ctrls_0_up_Prediction_WORD_SLICES_TAKEN_0;
  assign toplevel_decode_ctrls_0_up_Prediction_ALIGN_REDO_0 = AlignerPlugin_logic_extractors_0_redo;
  assign AlignerPlugin_logic_feeder_lanes_1_valid = AlignerPlugin_logic_extractors_1_valid;
  assign toplevel_decode_ctrls_0_up_LANE_SEL_1 = AlignerPlugin_logic_feeder_lanes_1_valid;
  always @(*) begin
    toplevel_decode_ctrls_0_up_Decode_INSTRUCTION_1 = AlignerPlugin_logic_extractors_1_ctx_instruction;
    if(AlignerPlugin_logic_feeder_lanes_1_isRvc) begin
      toplevel_decode_ctrls_0_up_Decode_INSTRUCTION_1 = AlignerPlugin_logic_feeder_lanes_1_withRvc_dec_inst;
    end
  end

  always @(*) begin
    toplevel_decode_ctrls_0_up_Decode_DECOMPRESSION_FAULT_1 = 1'b0;
    if(AlignerPlugin_logic_feeder_lanes_1_isRvc) begin
      toplevel_decode_ctrls_0_up_Decode_DECOMPRESSION_FAULT_1 = AlignerPlugin_logic_feeder_lanes_1_withRvc_dec_illegal;
    end
  end

  always @(*) begin
    toplevel_decode_ctrls_0_up_Decode_INSTRUCTION_RAW_1 = AlignerPlugin_logic_extractors_1_ctx_instruction;
    if(AlignerPlugin_logic_feeder_lanes_1_isRvc) begin
      toplevel_decode_ctrls_0_up_Decode_INSTRUCTION_RAW_1[31 : 16] = 16'h0;
    end
  end

  assign AlignerPlugin_logic_feeder_lanes_1_isRvc = (AlignerPlugin_logic_extractors_1_ctx_instruction[1 : 0] != 2'b11);
  always @(*) begin
    AlignerPlugin_logic_feeder_lanes_1_withRvc_dec_inst = 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
    case(switch_Rvc_l52_1)
      5'h0 : begin
        AlignerPlugin_logic_feeder_lanes_1_withRvc_dec_inst = {{{{{{{{{2'b00,AlignerPlugin_logic_extractors_1_ctx_instruction[10 : 7]},AlignerPlugin_logic_extractors_1_ctx_instruction[12 : 11]},AlignerPlugin_logic_extractors_1_ctx_instruction[5]},AlignerPlugin_logic_extractors_1_ctx_instruction[6]},2'b00},5'h02},3'b000},_zz_AlignerPlugin_logic_feeder_lanes_1_withRvc_dec_inst_1},7'h13};
      end
      5'h02 : begin
        AlignerPlugin_logic_feeder_lanes_1_withRvc_dec_inst = {{{{_zz_AlignerPlugin_logic_feeder_lanes_1_withRvc_dec_inst_2,_zz_AlignerPlugin_logic_feeder_lanes_1_withRvc_dec_inst},3'b010},_zz_AlignerPlugin_logic_feeder_lanes_1_withRvc_dec_inst_1},7'h03};
      end
      5'h05 : begin
        AlignerPlugin_logic_feeder_lanes_1_withRvc_dec_inst = {{{{{_zz_AlignerPlugin_logic_feeder_lanes_1_withRvc_dec_inst_3[11 : 5],_zz_AlignerPlugin_logic_feeder_lanes_1_withRvc_dec_inst_1},_zz_AlignerPlugin_logic_feeder_lanes_1_withRvc_dec_inst},3'b011},_zz_AlignerPlugin_logic_feeder_lanes_1_withRvc_dec_inst_3[4 : 0]},7'h27};
      end
      5'h06 : begin
        AlignerPlugin_logic_feeder_lanes_1_withRvc_dec_inst = {{{{{_zz_AlignerPlugin_logic_feeder_lanes_1_withRvc_dec_inst_2[11 : 5],_zz_AlignerPlugin_logic_feeder_lanes_1_withRvc_dec_inst_1},_zz_AlignerPlugin_logic_feeder_lanes_1_withRvc_dec_inst},3'b010},_zz_AlignerPlugin_logic_feeder_lanes_1_withRvc_dec_inst_2[4 : 0]},7'h23};
      end
      5'h08 : begin
        AlignerPlugin_logic_feeder_lanes_1_withRvc_dec_inst = {{{{_zz_AlignerPlugin_logic_feeder_lanes_1_withRvc_dec_inst_5,AlignerPlugin_logic_extractors_1_ctx_instruction[11 : 7]},3'b000},AlignerPlugin_logic_extractors_1_ctx_instruction[11 : 7]},7'h13};
      end
      5'h09 : begin
        AlignerPlugin_logic_feeder_lanes_1_withRvc_dec_inst = {{{{{_zz_AlignerPlugin_logic_feeder_lanes_1_withRvc_dec_inst_8[20],_zz_AlignerPlugin_logic_feeder_lanes_1_withRvc_dec_inst_8[10 : 1]},_zz_AlignerPlugin_logic_feeder_lanes_1_withRvc_dec_inst_8[11]},_zz_AlignerPlugin_logic_feeder_lanes_1_withRvc_dec_inst_8[19 : 12]},_zz_AlignerPlugin_logic_feeder_lanes_1_withRvc_dec_inst_20},7'h6f};
      end
      5'h0a : begin
        AlignerPlugin_logic_feeder_lanes_1_withRvc_dec_inst = {{{{_zz_AlignerPlugin_logic_feeder_lanes_1_withRvc_dec_inst_5,5'h0},3'b000},AlignerPlugin_logic_extractors_1_ctx_instruction[11 : 7]},7'h13};
      end
      5'h0b : begin
        AlignerPlugin_logic_feeder_lanes_1_withRvc_dec_inst = ((AlignerPlugin_logic_extractors_1_ctx_instruction[11 : 7] == 5'h02) ? {{{{{{{{_zz_AlignerPlugin_logic_feeder_lanes_1_withRvc_dec_inst_23,_zz_AlignerPlugin_logic_feeder_lanes_1_withRvc_dec_inst_24},_zz_AlignerPlugin_logic_feeder_lanes_1_withRvc_dec_inst_25},AlignerPlugin_logic_extractors_1_ctx_instruction[6]},4'b0000},AlignerPlugin_logic_extractors_1_ctx_instruction[11 : 7]},3'b000},AlignerPlugin_logic_extractors_1_ctx_instruction[11 : 7]},7'h13} : {{_zz_AlignerPlugin_logic_feeder_lanes_1_withRvc_dec_inst_26[31 : 12],AlignerPlugin_logic_extractors_1_ctx_instruction[11 : 7]},7'h37});
      end
      5'h0c : begin
        AlignerPlugin_logic_feeder_lanes_1_withRvc_dec_inst = _zz_AlignerPlugin_logic_feeder_lanes_1_withRvc_dec_inst_27;
      end
      5'h0d : begin
        AlignerPlugin_logic_feeder_lanes_1_withRvc_dec_inst = {{{{{_zz_AlignerPlugin_logic_feeder_lanes_1_withRvc_dec_inst_15[20],_zz_AlignerPlugin_logic_feeder_lanes_1_withRvc_dec_inst_15[10 : 1]},_zz_AlignerPlugin_logic_feeder_lanes_1_withRvc_dec_inst_15[11]},_zz_AlignerPlugin_logic_feeder_lanes_1_withRvc_dec_inst_15[19 : 12]},_zz_AlignerPlugin_logic_feeder_lanes_1_withRvc_dec_inst_19},7'h6f};
      end
      5'h0e : begin
        AlignerPlugin_logic_feeder_lanes_1_withRvc_dec_inst = {{{{{{{_zz_AlignerPlugin_logic_feeder_lanes_1_withRvc_dec_inst_18[12],_zz_AlignerPlugin_logic_feeder_lanes_1_withRvc_dec_inst_18[10 : 5]},_zz_AlignerPlugin_logic_feeder_lanes_1_withRvc_dec_inst_19},_zz_AlignerPlugin_logic_feeder_lanes_1_withRvc_dec_inst},3'b000},_zz_AlignerPlugin_logic_feeder_lanes_1_withRvc_dec_inst_18[4 : 1]},_zz_AlignerPlugin_logic_feeder_lanes_1_withRvc_dec_inst_18[11]},7'h63};
      end
      5'h0f : begin
        AlignerPlugin_logic_feeder_lanes_1_withRvc_dec_inst = {{{{{{{_zz_AlignerPlugin_logic_feeder_lanes_1_withRvc_dec_inst_18[12],_zz_AlignerPlugin_logic_feeder_lanes_1_withRvc_dec_inst_18[10 : 5]},_zz_AlignerPlugin_logic_feeder_lanes_1_withRvc_dec_inst_19},_zz_AlignerPlugin_logic_feeder_lanes_1_withRvc_dec_inst},3'b001},_zz_AlignerPlugin_logic_feeder_lanes_1_withRvc_dec_inst_18[4 : 1]},_zz_AlignerPlugin_logic_feeder_lanes_1_withRvc_dec_inst_18[11]},7'h63};
      end
      5'h10 : begin
        AlignerPlugin_logic_feeder_lanes_1_withRvc_dec_inst = {{{{{{6'h0,AlignerPlugin_logic_extractors_1_ctx_instruction[12]},AlignerPlugin_logic_extractors_1_ctx_instruction[6 : 2]},AlignerPlugin_logic_extractors_1_ctx_instruction[11 : 7]},3'b001},AlignerPlugin_logic_extractors_1_ctx_instruction[11 : 7]},7'h13};
      end
      5'h12 : begin
        AlignerPlugin_logic_feeder_lanes_1_withRvc_dec_inst = {{{{{{{{4'b0000,AlignerPlugin_logic_extractors_1_ctx_instruction[3 : 2]},AlignerPlugin_logic_extractors_1_ctx_instruction[12]},AlignerPlugin_logic_extractors_1_ctx_instruction[6 : 4]},2'b00},_zz_AlignerPlugin_logic_feeder_lanes_1_withRvc_dec_inst_21},3'b010},AlignerPlugin_logic_extractors_1_ctx_instruction[11 : 7]},7'h03};
      end
      5'h14 : begin
        AlignerPlugin_logic_feeder_lanes_1_withRvc_dec_inst = ((AlignerPlugin_logic_extractors_1_ctx_instruction[12 : 2] == 11'h400) ? 32'h00100073 : ((AlignerPlugin_logic_extractors_1_ctx_instruction[6 : 2] == 5'h0) ? {{{{12'h0,AlignerPlugin_logic_extractors_1_ctx_instruction[11 : 7]},3'b000},(AlignerPlugin_logic_extractors_1_ctx_instruction[12] ? _zz_AlignerPlugin_logic_feeder_lanes_1_withRvc_dec_inst_20 : _zz_AlignerPlugin_logic_feeder_lanes_1_withRvc_dec_inst_19)},7'h67} : {{{{{_zz_AlignerPlugin_logic_feeder_lanes_1_withRvc_dec_inst_31,_zz_AlignerPlugin_logic_feeder_lanes_1_withRvc_dec_inst_32},(_zz_AlignerPlugin_logic_feeder_lanes_1_withRvc_dec_inst_33 ? _zz_AlignerPlugin_logic_feeder_lanes_1_withRvc_dec_inst_34 : _zz_AlignerPlugin_logic_feeder_lanes_1_withRvc_dec_inst_19)},3'b000},AlignerPlugin_logic_extractors_1_ctx_instruction[11 : 7]},7'h33}));
      end
      5'h16 : begin
        AlignerPlugin_logic_feeder_lanes_1_withRvc_dec_inst = {{{{{_zz_AlignerPlugin_logic_feeder_lanes_1_withRvc_dec_inst_35[11 : 5],AlignerPlugin_logic_extractors_1_ctx_instruction[6 : 2]},_zz_AlignerPlugin_logic_feeder_lanes_1_withRvc_dec_inst_21},3'b010},_zz_AlignerPlugin_logic_feeder_lanes_1_withRvc_dec_inst_36[4 : 0]},7'h23};
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    AlignerPlugin_logic_feeder_lanes_1_withRvc_dec_illegal = 1'b0;
    case(switch_Rvc_l52_1)
      5'h0 : begin
        if(when_Rvc_l56_1) begin
          AlignerPlugin_logic_feeder_lanes_1_withRvc_dec_illegal = 1'b1;
        end
      end
      5'h02 : begin
      end
      5'h05 : begin
      end
      5'h06 : begin
      end
      5'h08 : begin
      end
      5'h09 : begin
      end
      5'h0a : begin
      end
      5'h0b : begin
        if(when_Rvc_l77_1) begin
          AlignerPlugin_logic_feeder_lanes_1_withRvc_dec_illegal = 1'b1;
        end
      end
      5'h0c : begin
      end
      5'h0d : begin
      end
      5'h0e : begin
      end
      5'h0f : begin
      end
      5'h10 : begin
      end
      5'h12 : begin
        if(when_Rvc_l98_1) begin
          AlignerPlugin_logic_feeder_lanes_1_withRvc_dec_illegal = 1'b1;
        end
      end
      5'h14 : begin
        if(when_Rvc_l111_1) begin
          AlignerPlugin_logic_feeder_lanes_1_withRvc_dec_illegal = 1'b1;
        end
      end
      5'h16 : begin
      end
      default : begin
        AlignerPlugin_logic_feeder_lanes_1_withRvc_dec_illegal = 1'b1;
      end
    endcase
  end

  assign _zz_AlignerPlugin_logic_feeder_lanes_1_withRvc_dec_inst = {2'b01,AlignerPlugin_logic_extractors_1_ctx_instruction[9 : 7]};
  assign _zz_AlignerPlugin_logic_feeder_lanes_1_withRvc_dec_inst_1 = {2'b01,AlignerPlugin_logic_extractors_1_ctx_instruction[4 : 2]};
  assign _zz_AlignerPlugin_logic_feeder_lanes_1_withRvc_dec_inst_2 = {{{{5'h0,AlignerPlugin_logic_extractors_1_ctx_instruction[5]},AlignerPlugin_logic_extractors_1_ctx_instruction[12 : 10]},AlignerPlugin_logic_extractors_1_ctx_instruction[6]},2'b00};
  assign _zz_AlignerPlugin_logic_feeder_lanes_1_withRvc_dec_inst_3 = {{{4'b0000,AlignerPlugin_logic_extractors_1_ctx_instruction[6 : 5]},AlignerPlugin_logic_extractors_1_ctx_instruction[12 : 10]},3'b000};
  assign _zz_AlignerPlugin_logic_feeder_lanes_1_withRvc_dec_inst_4 = AlignerPlugin_logic_extractors_1_ctx_instruction[12];
  always @(*) begin
    _zz_AlignerPlugin_logic_feeder_lanes_1_withRvc_dec_inst_5[11] = _zz_AlignerPlugin_logic_feeder_lanes_1_withRvc_dec_inst_4;
    _zz_AlignerPlugin_logic_feeder_lanes_1_withRvc_dec_inst_5[10] = _zz_AlignerPlugin_logic_feeder_lanes_1_withRvc_dec_inst_4;
    _zz_AlignerPlugin_logic_feeder_lanes_1_withRvc_dec_inst_5[9] = _zz_AlignerPlugin_logic_feeder_lanes_1_withRvc_dec_inst_4;
    _zz_AlignerPlugin_logic_feeder_lanes_1_withRvc_dec_inst_5[8] = _zz_AlignerPlugin_logic_feeder_lanes_1_withRvc_dec_inst_4;
    _zz_AlignerPlugin_logic_feeder_lanes_1_withRvc_dec_inst_5[7] = _zz_AlignerPlugin_logic_feeder_lanes_1_withRvc_dec_inst_4;
    _zz_AlignerPlugin_logic_feeder_lanes_1_withRvc_dec_inst_5[6] = _zz_AlignerPlugin_logic_feeder_lanes_1_withRvc_dec_inst_4;
    _zz_AlignerPlugin_logic_feeder_lanes_1_withRvc_dec_inst_5[5] = _zz_AlignerPlugin_logic_feeder_lanes_1_withRvc_dec_inst_4;
    _zz_AlignerPlugin_logic_feeder_lanes_1_withRvc_dec_inst_5[4 : 0] = AlignerPlugin_logic_extractors_1_ctx_instruction[6 : 2];
  end

  assign _zz_AlignerPlugin_logic_feeder_lanes_1_withRvc_dec_inst_6 = AlignerPlugin_logic_extractors_1_ctx_instruction[12];
  always @(*) begin
    _zz_AlignerPlugin_logic_feeder_lanes_1_withRvc_dec_inst_7[9] = _zz_AlignerPlugin_logic_feeder_lanes_1_withRvc_dec_inst_6;
    _zz_AlignerPlugin_logic_feeder_lanes_1_withRvc_dec_inst_7[8] = _zz_AlignerPlugin_logic_feeder_lanes_1_withRvc_dec_inst_6;
    _zz_AlignerPlugin_logic_feeder_lanes_1_withRvc_dec_inst_7[7] = _zz_AlignerPlugin_logic_feeder_lanes_1_withRvc_dec_inst_6;
    _zz_AlignerPlugin_logic_feeder_lanes_1_withRvc_dec_inst_7[6] = _zz_AlignerPlugin_logic_feeder_lanes_1_withRvc_dec_inst_6;
    _zz_AlignerPlugin_logic_feeder_lanes_1_withRvc_dec_inst_7[5] = _zz_AlignerPlugin_logic_feeder_lanes_1_withRvc_dec_inst_6;
    _zz_AlignerPlugin_logic_feeder_lanes_1_withRvc_dec_inst_7[4] = _zz_AlignerPlugin_logic_feeder_lanes_1_withRvc_dec_inst_6;
    _zz_AlignerPlugin_logic_feeder_lanes_1_withRvc_dec_inst_7[3] = _zz_AlignerPlugin_logic_feeder_lanes_1_withRvc_dec_inst_6;
    _zz_AlignerPlugin_logic_feeder_lanes_1_withRvc_dec_inst_7[2] = _zz_AlignerPlugin_logic_feeder_lanes_1_withRvc_dec_inst_6;
    _zz_AlignerPlugin_logic_feeder_lanes_1_withRvc_dec_inst_7[1] = _zz_AlignerPlugin_logic_feeder_lanes_1_withRvc_dec_inst_6;
    _zz_AlignerPlugin_logic_feeder_lanes_1_withRvc_dec_inst_7[0] = _zz_AlignerPlugin_logic_feeder_lanes_1_withRvc_dec_inst_6;
  end

  assign _zz_AlignerPlugin_logic_feeder_lanes_1_withRvc_dec_inst_8 = {{{{{{{{_zz_AlignerPlugin_logic_feeder_lanes_1_withRvc_dec_inst_7,AlignerPlugin_logic_extractors_1_ctx_instruction[8]},AlignerPlugin_logic_extractors_1_ctx_instruction[10 : 9]},AlignerPlugin_logic_extractors_1_ctx_instruction[6]},AlignerPlugin_logic_extractors_1_ctx_instruction[7]},AlignerPlugin_logic_extractors_1_ctx_instruction[2]},AlignerPlugin_logic_extractors_1_ctx_instruction[11]},AlignerPlugin_logic_extractors_1_ctx_instruction[5 : 3]},1'b0};
  assign _zz_AlignerPlugin_logic_feeder_lanes_1_withRvc_dec_inst_9 = AlignerPlugin_logic_extractors_1_ctx_instruction[12];
  always @(*) begin
    _zz_AlignerPlugin_logic_feeder_lanes_1_withRvc_dec_inst_10[14] = _zz_AlignerPlugin_logic_feeder_lanes_1_withRvc_dec_inst_9;
    _zz_AlignerPlugin_logic_feeder_lanes_1_withRvc_dec_inst_10[13] = _zz_AlignerPlugin_logic_feeder_lanes_1_withRvc_dec_inst_9;
    _zz_AlignerPlugin_logic_feeder_lanes_1_withRvc_dec_inst_10[12] = _zz_AlignerPlugin_logic_feeder_lanes_1_withRvc_dec_inst_9;
    _zz_AlignerPlugin_logic_feeder_lanes_1_withRvc_dec_inst_10[11] = _zz_AlignerPlugin_logic_feeder_lanes_1_withRvc_dec_inst_9;
    _zz_AlignerPlugin_logic_feeder_lanes_1_withRvc_dec_inst_10[10] = _zz_AlignerPlugin_logic_feeder_lanes_1_withRvc_dec_inst_9;
    _zz_AlignerPlugin_logic_feeder_lanes_1_withRvc_dec_inst_10[9] = _zz_AlignerPlugin_logic_feeder_lanes_1_withRvc_dec_inst_9;
    _zz_AlignerPlugin_logic_feeder_lanes_1_withRvc_dec_inst_10[8] = _zz_AlignerPlugin_logic_feeder_lanes_1_withRvc_dec_inst_9;
    _zz_AlignerPlugin_logic_feeder_lanes_1_withRvc_dec_inst_10[7] = _zz_AlignerPlugin_logic_feeder_lanes_1_withRvc_dec_inst_9;
    _zz_AlignerPlugin_logic_feeder_lanes_1_withRvc_dec_inst_10[6] = _zz_AlignerPlugin_logic_feeder_lanes_1_withRvc_dec_inst_9;
    _zz_AlignerPlugin_logic_feeder_lanes_1_withRvc_dec_inst_10[5] = _zz_AlignerPlugin_logic_feeder_lanes_1_withRvc_dec_inst_9;
    _zz_AlignerPlugin_logic_feeder_lanes_1_withRvc_dec_inst_10[4] = _zz_AlignerPlugin_logic_feeder_lanes_1_withRvc_dec_inst_9;
    _zz_AlignerPlugin_logic_feeder_lanes_1_withRvc_dec_inst_10[3] = _zz_AlignerPlugin_logic_feeder_lanes_1_withRvc_dec_inst_9;
    _zz_AlignerPlugin_logic_feeder_lanes_1_withRvc_dec_inst_10[2] = _zz_AlignerPlugin_logic_feeder_lanes_1_withRvc_dec_inst_9;
    _zz_AlignerPlugin_logic_feeder_lanes_1_withRvc_dec_inst_10[1] = _zz_AlignerPlugin_logic_feeder_lanes_1_withRvc_dec_inst_9;
    _zz_AlignerPlugin_logic_feeder_lanes_1_withRvc_dec_inst_10[0] = _zz_AlignerPlugin_logic_feeder_lanes_1_withRvc_dec_inst_9;
  end

  assign _zz_AlignerPlugin_logic_feeder_lanes_1_withRvc_dec_inst_11 = AlignerPlugin_logic_extractors_1_ctx_instruction[12];
  always @(*) begin
    _zz_AlignerPlugin_logic_feeder_lanes_1_withRvc_dec_inst_12[2] = _zz_AlignerPlugin_logic_feeder_lanes_1_withRvc_dec_inst_11;
    _zz_AlignerPlugin_logic_feeder_lanes_1_withRvc_dec_inst_12[1] = _zz_AlignerPlugin_logic_feeder_lanes_1_withRvc_dec_inst_11;
    _zz_AlignerPlugin_logic_feeder_lanes_1_withRvc_dec_inst_12[0] = _zz_AlignerPlugin_logic_feeder_lanes_1_withRvc_dec_inst_11;
  end

  assign _zz_AlignerPlugin_logic_feeder_lanes_1_withRvc_dec_inst_13 = AlignerPlugin_logic_extractors_1_ctx_instruction[12];
  always @(*) begin
    _zz_AlignerPlugin_logic_feeder_lanes_1_withRvc_dec_inst_14[9] = _zz_AlignerPlugin_logic_feeder_lanes_1_withRvc_dec_inst_13;
    _zz_AlignerPlugin_logic_feeder_lanes_1_withRvc_dec_inst_14[8] = _zz_AlignerPlugin_logic_feeder_lanes_1_withRvc_dec_inst_13;
    _zz_AlignerPlugin_logic_feeder_lanes_1_withRvc_dec_inst_14[7] = _zz_AlignerPlugin_logic_feeder_lanes_1_withRvc_dec_inst_13;
    _zz_AlignerPlugin_logic_feeder_lanes_1_withRvc_dec_inst_14[6] = _zz_AlignerPlugin_logic_feeder_lanes_1_withRvc_dec_inst_13;
    _zz_AlignerPlugin_logic_feeder_lanes_1_withRvc_dec_inst_14[5] = _zz_AlignerPlugin_logic_feeder_lanes_1_withRvc_dec_inst_13;
    _zz_AlignerPlugin_logic_feeder_lanes_1_withRvc_dec_inst_14[4] = _zz_AlignerPlugin_logic_feeder_lanes_1_withRvc_dec_inst_13;
    _zz_AlignerPlugin_logic_feeder_lanes_1_withRvc_dec_inst_14[3] = _zz_AlignerPlugin_logic_feeder_lanes_1_withRvc_dec_inst_13;
    _zz_AlignerPlugin_logic_feeder_lanes_1_withRvc_dec_inst_14[2] = _zz_AlignerPlugin_logic_feeder_lanes_1_withRvc_dec_inst_13;
    _zz_AlignerPlugin_logic_feeder_lanes_1_withRvc_dec_inst_14[1] = _zz_AlignerPlugin_logic_feeder_lanes_1_withRvc_dec_inst_13;
    _zz_AlignerPlugin_logic_feeder_lanes_1_withRvc_dec_inst_14[0] = _zz_AlignerPlugin_logic_feeder_lanes_1_withRvc_dec_inst_13;
  end

  assign _zz_AlignerPlugin_logic_feeder_lanes_1_withRvc_dec_inst_15 = {{{{{{{{_zz_AlignerPlugin_logic_feeder_lanes_1_withRvc_dec_inst_14,AlignerPlugin_logic_extractors_1_ctx_instruction[8]},AlignerPlugin_logic_extractors_1_ctx_instruction[10 : 9]},AlignerPlugin_logic_extractors_1_ctx_instruction[6]},AlignerPlugin_logic_extractors_1_ctx_instruction[7]},AlignerPlugin_logic_extractors_1_ctx_instruction[2]},AlignerPlugin_logic_extractors_1_ctx_instruction[11]},AlignerPlugin_logic_extractors_1_ctx_instruction[5 : 3]},1'b0};
  assign _zz_AlignerPlugin_logic_feeder_lanes_1_withRvc_dec_inst_16 = AlignerPlugin_logic_extractors_1_ctx_instruction[12];
  always @(*) begin
    _zz_AlignerPlugin_logic_feeder_lanes_1_withRvc_dec_inst_17[4] = _zz_AlignerPlugin_logic_feeder_lanes_1_withRvc_dec_inst_16;
    _zz_AlignerPlugin_logic_feeder_lanes_1_withRvc_dec_inst_17[3] = _zz_AlignerPlugin_logic_feeder_lanes_1_withRvc_dec_inst_16;
    _zz_AlignerPlugin_logic_feeder_lanes_1_withRvc_dec_inst_17[2] = _zz_AlignerPlugin_logic_feeder_lanes_1_withRvc_dec_inst_16;
    _zz_AlignerPlugin_logic_feeder_lanes_1_withRvc_dec_inst_17[1] = _zz_AlignerPlugin_logic_feeder_lanes_1_withRvc_dec_inst_16;
    _zz_AlignerPlugin_logic_feeder_lanes_1_withRvc_dec_inst_17[0] = _zz_AlignerPlugin_logic_feeder_lanes_1_withRvc_dec_inst_16;
  end

  assign _zz_AlignerPlugin_logic_feeder_lanes_1_withRvc_dec_inst_18 = {{{{{_zz_AlignerPlugin_logic_feeder_lanes_1_withRvc_dec_inst_17,AlignerPlugin_logic_extractors_1_ctx_instruction[6 : 5]},AlignerPlugin_logic_extractors_1_ctx_instruction[2]},AlignerPlugin_logic_extractors_1_ctx_instruction[11 : 10]},AlignerPlugin_logic_extractors_1_ctx_instruction[4 : 3]},1'b0};
  assign _zz_AlignerPlugin_logic_feeder_lanes_1_withRvc_dec_inst_19 = 5'h0;
  assign _zz_AlignerPlugin_logic_feeder_lanes_1_withRvc_dec_inst_20 = 5'h01;
  assign _zz_AlignerPlugin_logic_feeder_lanes_1_withRvc_dec_inst_21 = 5'h02;
  assign switch_Rvc_l52_1 = {AlignerPlugin_logic_extractors_1_ctx_instruction[1 : 0],AlignerPlugin_logic_extractors_1_ctx_instruction[15 : 13]};
  assign when_Rvc_l56_1 = (AlignerPlugin_logic_extractors_1_ctx_instruction[12 : 5] == 8'h0);
  assign when_Rvc_l77_1 = ((AlignerPlugin_logic_extractors_1_ctx_instruction[6 : 2] == 5'h0) && (AlignerPlugin_logic_extractors_1_ctx_instruction[12] == 1'b0));
  assign _zz_AlignerPlugin_logic_feeder_lanes_1_withRvc_dec_inst_22 = {{{{_zz__zz_AlignerPlugin_logic_feeder_lanes_1_withRvc_dec_inst_22,_zz_AlignerPlugin_logic_feeder_lanes_1_withRvc_dec_inst},3'b101},_zz_AlignerPlugin_logic_feeder_lanes_1_withRvc_dec_inst},7'h13};
  assign when_Rvc_l98_1 = (AlignerPlugin_logic_extractors_1_ctx_instruction[11 : 7] == 5'h0);
  assign when_Rvc_l111_1 = (((AlignerPlugin_logic_extractors_1_ctx_instruction[11 : 7] == 5'h0) && (AlignerPlugin_logic_extractors_1_ctx_instruction[6 : 2] == 5'h0)) && (AlignerPlugin_logic_extractors_1_ctx_instruction[12] == 1'b0));
  assign _zz_toplevel_decode_ctrls_0_up_Decode_INSTRUCTION_SLICE_COUNT_1 = AlignerPlugin_logic_extractors_1_localMask;
  assign _zz_toplevel_decode_ctrls_0_up_Decode_INSTRUCTION_SLICE_COUNT_1_1 = {_zz_toplevel_decode_ctrls_0_up_Decode_INSTRUCTION_SLICE_COUNT_1[0],_zz_toplevel_decode_ctrls_0_up_Decode_INSTRUCTION_SLICE_COUNT_1[1]};
  assign _zz_toplevel_decode_ctrls_0_up_Decode_INSTRUCTION_SLICE_COUNT_1_2 = _zz_toplevel_decode_ctrls_0_up_Decode_INSTRUCTION_SLICE_COUNT_1_1[0];
  always @(*) begin
    _zz_toplevel_decode_ctrls_0_up_Decode_INSTRUCTION_SLICE_COUNT_1_3[0] = (_zz_toplevel_decode_ctrls_0_up_Decode_INSTRUCTION_SLICE_COUNT_1_2 && (! 1'b0));
    _zz_toplevel_decode_ctrls_0_up_Decode_INSTRUCTION_SLICE_COUNT_1_3[1] = (_zz_toplevel_decode_ctrls_0_up_Decode_INSTRUCTION_SLICE_COUNT_1_1[1] && (! _zz_toplevel_decode_ctrls_0_up_Decode_INSTRUCTION_SLICE_COUNT_1_2));
  end

  assign _zz_toplevel_decode_ctrls_0_up_Decode_INSTRUCTION_SLICE_COUNT_1_4 = _zz_toplevel_decode_ctrls_0_up_Decode_INSTRUCTION_SLICE_COUNT_1_3;
  assign _zz_toplevel_decode_ctrls_0_up_Decode_INSTRUCTION_SLICE_COUNT_1_5 = _zz__zz_toplevel_decode_ctrls_0_up_Decode_INSTRUCTION_SLICE_COUNT_1_5[1];
  assign toplevel_decode_ctrls_0_up_Decode_INSTRUCTION_SLICE_COUNT_1 = _zz_toplevel_decode_ctrls_0_up_Decode_INSTRUCTION_SLICE_COUNT_1_5;
  assign toplevel_decode_ctrls_0_up_PC_1 = AlignerPlugin_logic_extractors_1_ctx_pc;
  assign toplevel_decode_ctrls_0_up_Decode_DOP_ID_1 = (toplevel_decode_ctrls_0_down_Decode_DOP_ID_0 + _zz_toplevel_decode_ctrls_0_up_Decode_DOP_ID_1);
  assign toplevel_decode_ctrls_0_up_Fetch_ID_1 = AlignerPlugin_logic_extractors_1_ctx_hm_Fetch_ID;
  assign toplevel_decode_ctrls_0_up_GSharePlugin_GSHARE_COUNTER_1_0 = AlignerPlugin_logic_extractors_1_ctx_hm_GSharePlugin_GSHARE_COUNTER_0;
  assign toplevel_decode_ctrls_0_up_GSharePlugin_GSHARE_COUNTER_1_1 = AlignerPlugin_logic_extractors_1_ctx_hm_GSharePlugin_GSHARE_COUNTER_1;
  assign toplevel_decode_ctrls_0_up_GSharePlugin_GSHARE_COUNTER_1_2 = AlignerPlugin_logic_extractors_1_ctx_hm_GSharePlugin_GSHARE_COUNTER_2;
  assign toplevel_decode_ctrls_0_up_GSharePlugin_GSHARE_COUNTER_1_3 = AlignerPlugin_logic_extractors_1_ctx_hm_GSharePlugin_GSHARE_COUNTER_3;
  assign toplevel_decode_ctrls_0_up_Prediction_BRANCH_HISTORY_1 = AlignerPlugin_logic_extractors_1_ctx_hm_Prediction_BRANCH_HISTORY;
  assign toplevel_decode_ctrls_0_up_Prediction_WORD_SLICES_BRANCH_1 = AlignerPlugin_logic_extractors_1_ctx_hm_Prediction_WORD_SLICES_BRANCH;
  assign toplevel_decode_ctrls_0_up_Prediction_WORD_SLICES_TAKEN_1 = AlignerPlugin_logic_extractors_1_ctx_hm_Prediction_WORD_SLICES_TAKEN;
  assign toplevel_decode_ctrls_0_up_Prediction_WORD_JUMP_PC_1 = AlignerPlugin_logic_extractors_1_ctx_hm_Prediction_WORD_JUMP_PC;
  assign toplevel_decode_ctrls_0_up_Prediction_WORD_JUMPED_1 = AlignerPlugin_logic_extractors_1_ctx_hm_Prediction_WORD_JUMPED;
  assign toplevel_decode_ctrls_0_up_Prediction_WORD_JUMP_SLICE_1 = AlignerPlugin_logic_extractors_1_ctx_hm_Prediction_WORD_JUMP_SLICE;
  assign toplevel_decode_ctrls_0_up_TRAP_1 = AlignerPlugin_logic_extractors_1_ctx_trap;
  assign AlignerPlugin_logic_feeder_lanes_1_onBtb_pcLastSlice = (toplevel_decode_ctrls_0_up_PC_1[2 : 1] + _zz_AlignerPlugin_logic_feeder_lanes_1_onBtb_pcLastSlice);
  assign AlignerPlugin_logic_feeder_lanes_1_onBtb_didPrediction = (toplevel_decode_ctrls_0_up_Prediction_WORD_JUMP_SLICE_1 <= AlignerPlugin_logic_feeder_lanes_1_onBtb_pcLastSlice);
  assign toplevel_decode_ctrls_0_up_Prediction_ALIGNED_JUMPED_1 = (toplevel_decode_ctrls_0_up_Prediction_WORD_JUMPED_1 && AlignerPlugin_logic_feeder_lanes_1_onBtb_didPrediction);
  assign toplevel_decode_ctrls_0_up_Prediction_ALIGNED_JUMPED_PC_1 = toplevel_decode_ctrls_0_up_Prediction_WORD_JUMP_PC_1;
  assign toplevel_decode_ctrls_0_up_Prediction_ALIGNED_SLICES_BRANCH_1 = toplevel_decode_ctrls_0_up_Prediction_WORD_SLICES_BRANCH_1;
  assign toplevel_decode_ctrls_0_up_Prediction_ALIGNED_SLICES_TAKEN_1 = toplevel_decode_ctrls_0_up_Prediction_WORD_SLICES_TAKEN_1;
  assign toplevel_decode_ctrls_0_up_Prediction_ALIGN_REDO_1 = AlignerPlugin_logic_extractors_1_redo;
  assign toplevel_decode_ctrls_0_up_valid = (|{AlignerPlugin_logic_feeder_lanes_1_valid,AlignerPlugin_logic_feeder_lanes_0_valid});
  assign _zz_AlignerPlugin_logic_slices_data_0 = {fetch_logic_ctrls_2_down_Fetch_WORD,AlignerPlugin_logic_buffer_data};
  assign AlignerPlugin_logic_slices_data_0 = _zz_AlignerPlugin_logic_slices_data_0[15 : 0];
  assign AlignerPlugin_logic_slices_data_1 = _zz_AlignerPlugin_logic_slices_data_0[31 : 16];
  assign AlignerPlugin_logic_slices_data_2 = _zz_AlignerPlugin_logic_slices_data_0[47 : 32];
  assign AlignerPlugin_logic_slices_data_3 = _zz_AlignerPlugin_logic_slices_data_0[63 : 48];
  assign AlignerPlugin_logic_slices_data_4 = _zz_AlignerPlugin_logic_slices_data_0[79 : 64];
  assign AlignerPlugin_logic_slices_data_5 = _zz_AlignerPlugin_logic_slices_data_0[95 : 80];
  assign AlignerPlugin_logic_slices_data_6 = _zz_AlignerPlugin_logic_slices_data_0[111 : 96];
  assign AlignerPlugin_logic_slices_data_7 = _zz_AlignerPlugin_logic_slices_data_0[127 : 112];
  assign AlignerPlugin_logic_slices_mask = {fetch_logic_ctrls_2_down_AlignerPlugin_logic_FETCH_MASK,AlignerPlugin_logic_buffer_mask};
  assign AlignerPlugin_logic_slices_last = {fetch_logic_ctrls_2_down_AlignerPlugin_logic_FETCH_LAST,AlignerPlugin_logic_buffer_last};
  assign when_AlignerPlugin_l243 = (! fetch_logic_ctrls_2_down_valid);
  assign when_AlignerPlugin_l244 = (AlignerPlugin_logic_extractors_0_usageMask[7 : 4] != 4'b0000);
  assign when_AlignerPlugin_l244_1 = (AlignerPlugin_logic_extractors_1_usageMask[7 : 4] != 4'b0000);
  assign AlignerPlugin_logic_buffer_downFire = (toplevel_decode_ctrls_0_up_isReady || toplevel_decode_ctrls_0_up_isCancel);
  assign AlignerPlugin_logic_buffer_usedMask = ((AlignerPlugin_logic_extractors_0_valid ? AlignerPlugin_logic_extractors_0_usageMask : 8'h0) | (AlignerPlugin_logic_extractors_1_valid ? AlignerPlugin_logic_extractors_1_usageMask : 8'h0));
  assign AlignerPlugin_logic_buffer_haltUp = ((|(AlignerPlugin_logic_buffer_mask & (~ (AlignerPlugin_logic_buffer_downFire ? AlignerPlugin_logic_buffer_usedMask[3 : 0] : 4'b0000)))) || AlignerPlugin_api_haltIt);
  assign fetch_logic_ctrls_2_down_ready = ((! fetch_logic_ctrls_2_down_valid) || (! AlignerPlugin_logic_buffer_haltUp));
  assign when_AlignerPlugin_l259 = ((fetch_logic_ctrls_2_down_isValid && fetch_logic_ctrls_2_down_isReady) && (! fetch_logic_ctrls_2_down_isCancel));
  always @(*) begin
    CsrAccessPlugin_bus_decode_exception = 1'b0;
    if(when_PrivilegedPlugin_l679) begin
      CsrAccessPlugin_bus_decode_exception = 1'b1;
    end
    if(when_CsrAccessPlugin_l155) begin
      if(when_MmuPlugin_l212) begin
        CsrAccessPlugin_bus_decode_exception = 1'b1;
      end
    end
  end

  always @(*) begin
    CsrAccessPlugin_bus_decode_trap = 1'b0;
    if(when_CsrAccessPlugin_l155) begin
      if(!when_MmuPlugin_l212) begin
        CsrAccessPlugin_bus_decode_trap = 1'b1;
      end
    end
    if(when_CsrAccessPlugin_l155_1) begin
      if(CsrAccessPlugin_bus_decode_write) begin
        CsrAccessPlugin_bus_decode_trap = 1'b1;
      end
    end
  end

  always @(*) begin
    CsrAccessPlugin_bus_decode_trapCode = 4'bxxxx;
    if(when_CsrAccessPlugin_l155) begin
      if(!when_MmuPlugin_l212) begin
        CsrAccessPlugin_bus_decode_trapCode = 4'b0110;
      end
    end
    if(when_CsrAccessPlugin_l155_1) begin
      if(CsrAccessPlugin_bus_decode_write) begin
        CsrAccessPlugin_bus_decode_trapCode = 4'b0101;
      end
    end
  end

  always @(*) begin
    CsrAccessPlugin_bus_read_halt = 1'b0;
    if(when_CsrRamPlugin_l77) begin
      CsrAccessPlugin_bus_read_halt = 1'b1;
    end
  end

  always @(*) begin
    CsrAccessPlugin_bus_write_halt = 1'b0;
    if(when_CsrRamPlugin_l88) begin
      CsrAccessPlugin_bus_write_halt = 1'b1;
    end
  end

  assign FetchL1Plugin_logic_banks_0_read_rsp = FetchL1Plugin_logic_banks_0_mem_spinal_port1;
  assign fetch_logic_ctrls_1_down_FetchL1Plugin_logic_BANKS_WORDS_0 = FetchL1Plugin_logic_banks_0_read_rsp;
  assign FetchL1Plugin_logic_banks_1_read_rsp = FetchL1Plugin_logic_banks_1_mem_spinal_port1;
  assign fetch_logic_ctrls_1_down_FetchL1Plugin_logic_BANKS_WORDS_1 = FetchL1Plugin_logic_banks_1_read_rsp;
  always @(*) begin
    FetchL1Plugin_logic_waysWrite_mask = 2'b00;
    if(when_FetchL1Plugin_l220) begin
      FetchL1Plugin_logic_waysWrite_mask = 2'b11;
    end
    if(FetchL1Plugin_logic_invalidate_done) begin
      if(when_FetchL1Plugin_l324) begin
        FetchL1Plugin_logic_waysWrite_mask[FetchL1Plugin_logic_refill_onRsp_wayToAllocate] = 1'b1;
      end
    end
  end

  always @(*) begin
    FetchL1Plugin_logic_waysWrite_address = 6'bxxxxxx;
    if(when_FetchL1Plugin_l220) begin
      FetchL1Plugin_logic_waysWrite_address = FetchL1Plugin_logic_invalidate_counter[5:0];
    end
    if(FetchL1Plugin_logic_invalidate_done) begin
      FetchL1Plugin_logic_waysWrite_address = FetchL1Plugin_logic_refill_onRsp_address[11 : 6];
    end
  end

  always @(*) begin
    FetchL1Plugin_logic_waysWrite_tag_loaded = 1'bx;
    if(when_FetchL1Plugin_l220) begin
      FetchL1Plugin_logic_waysWrite_tag_loaded = 1'b0;
    end
    if(FetchL1Plugin_logic_invalidate_done) begin
      FetchL1Plugin_logic_waysWrite_tag_loaded = 1'b1;
    end
  end

  always @(*) begin
    FetchL1Plugin_logic_waysWrite_tag_error = 1'bx;
    if(FetchL1Plugin_logic_invalidate_done) begin
      FetchL1Plugin_logic_waysWrite_tag_error = (FetchL1Plugin_logic_bus_rsp_valid && FetchL1Plugin_logic_bus_rsp_payload_error);
    end
  end

  always @(*) begin
    FetchL1Plugin_logic_waysWrite_tag_address = 20'bxxxxxxxxxxxxxxxxxxxx;
    if(FetchL1Plugin_logic_invalidate_done) begin
      FetchL1Plugin_logic_waysWrite_tag_address = FetchL1Plugin_logic_refill_onRsp_address[31 : 12];
    end
  end

  assign _zz_FetchL1Plugin_logic_ways_0_read_rsp_loaded = FetchL1Plugin_logic_ways_0_mem_spinal_port1;
  assign FetchL1Plugin_logic_ways_0_read_rsp_loaded = _zz_FetchL1Plugin_logic_ways_0_read_rsp_loaded[0];
  assign FetchL1Plugin_logic_ways_0_read_rsp_error = _zz_FetchL1Plugin_logic_ways_0_read_rsp_loaded[1];
  assign FetchL1Plugin_logic_ways_0_read_rsp_address = _zz_FetchL1Plugin_logic_ways_0_read_rsp_loaded[21 : 2];
  assign fetch_logic_ctrls_1_down_FetchL1Plugin_logic_WAYS_TAGS_0_loaded = FetchL1Plugin_logic_ways_0_read_rsp_loaded;
  assign fetch_logic_ctrls_1_down_FetchL1Plugin_logic_WAYS_TAGS_0_error = FetchL1Plugin_logic_ways_0_read_rsp_error;
  assign fetch_logic_ctrls_1_down_FetchL1Plugin_logic_WAYS_TAGS_0_address = FetchL1Plugin_logic_ways_0_read_rsp_address;
  assign _zz_FetchL1Plugin_logic_ways_1_read_rsp_loaded = FetchL1Plugin_logic_ways_1_mem_spinal_port1;
  assign FetchL1Plugin_logic_ways_1_read_rsp_loaded = _zz_FetchL1Plugin_logic_ways_1_read_rsp_loaded[0];
  assign FetchL1Plugin_logic_ways_1_read_rsp_error = _zz_FetchL1Plugin_logic_ways_1_read_rsp_loaded[1];
  assign FetchL1Plugin_logic_ways_1_read_rsp_address = _zz_FetchL1Plugin_logic_ways_1_read_rsp_loaded[21 : 2];
  assign fetch_logic_ctrls_1_down_FetchL1Plugin_logic_WAYS_TAGS_1_loaded = FetchL1Plugin_logic_ways_1_read_rsp_loaded;
  assign fetch_logic_ctrls_1_down_FetchL1Plugin_logic_WAYS_TAGS_1_error = FetchL1Plugin_logic_ways_1_read_rsp_error;
  assign fetch_logic_ctrls_1_down_FetchL1Plugin_logic_WAYS_TAGS_1_address = FetchL1Plugin_logic_ways_1_read_rsp_address;
  assign FetchL1Plugin_logic_plru_read_rsp_0 = FetchL1Plugin_logic_plru_mem_spinal_port1[0 : 0];
  assign fetch_logic_ctrls_1_down_FetchL1Plugin_logic_PLRU_READ_0 = FetchL1Plugin_logic_plru_read_rsp_0;
  assign FetchL1Plugin_logic_invalidate_cmd_valid = (|TrapPlugin_logic_fetchL1Invalidate_0_cmd_valid);
  always @(*) begin
    FetchL1Plugin_logic_invalidate_canStart = 1'b1;
    if(when_FetchL1Plugin_l293) begin
      FetchL1Plugin_logic_invalidate_canStart = 1'b0;
    end
  end

  assign FetchL1Plugin_logic_invalidate_counterIncr = (FetchL1Plugin_logic_invalidate_counter + 7'h01);
  assign FetchL1Plugin_logic_invalidate_done = FetchL1Plugin_logic_invalidate_counter[6];
  assign FetchL1Plugin_logic_invalidate_last = FetchL1Plugin_logic_invalidate_counterIncr[6];
  assign when_FetchL1Plugin_l220 = (! FetchL1Plugin_logic_invalidate_done);
  assign when_FetchL1Plugin_l227 = ((FetchL1Plugin_logic_invalidate_done && FetchL1Plugin_logic_invalidate_cmd_valid) && FetchL1Plugin_logic_invalidate_canStart);
  always @(*) begin
    TrapPlugin_logic_fetchL1Invalidate_0_cmd_ready = 1'b0;
    if(when_FetchL1Plugin_l232) begin
      if(FetchL1Plugin_logic_invalidate_last) begin
        TrapPlugin_logic_fetchL1Invalidate_0_cmd_ready = 1'b1;
      end
    end
  end

  assign when_FetchL1Plugin_l232 = (! FetchL1Plugin_logic_invalidate_done);
  assign fetch_logic_ctrls_0_haltRequest_FetchL1Plugin_l233 = _zz_fetch_logic_ctrls_0_haltRequest_FetchL1Plugin_l233;
  assign FetchL1Plugin_logic_refill_slots_0_askCmd = (FetchL1Plugin_logic_refill_slots_0_valid && (! FetchL1Plugin_logic_refill_slots_0_cmdSent));
  assign FetchL1Plugin_logic_refill_hazard = (|(FetchL1Plugin_logic_refill_slots_0_valid && (FetchL1Plugin_logic_refill_slots_0_address[11 : 6] == FetchL1Plugin_logic_refill_start_address[11 : 6])));
  assign when_FetchL1Plugin_l271 = ((FetchL1Plugin_logic_refill_start_valid && FetchL1Plugin_logic_invalidate_done) && (! FetchL1Plugin_logic_refill_hazard));
  assign when_FetchL1Plugin_l293 = ((|FetchL1Plugin_logic_refill_slots_0_valid) || FetchL1Plugin_logic_refill_start_valid);
  assign FetchL1Plugin_logic_refill_onCmd_oh = (FetchL1Plugin_logic_refill_slots_0_askCmd && 1'b1);
  assign FetchL1Plugin_logic_bus_cmd_valid = (|FetchL1Plugin_logic_refill_onCmd_oh);
  assign FetchL1Plugin_logic_bus_cmd_payload_address = {FetchL1Plugin_logic_refill_slots_0_address[31 : 6],6'h0};
  assign FetchL1Plugin_logic_bus_cmd_payload_io = FetchL1Plugin_logic_refill_slots_0_isIo;
  assign FetchL1Plugin_logic_refill_onRsp_holdHarts = ((|FetchL1Plugin_logic_waysWrite_mask) || (|((FetchL1Plugin_logic_refill_slots_0_valid && (FetchL1Plugin_logic_refill_slots_0_address[11 : 6] == fetch_logic_ctrls_0_down_Fetch_WORD_PC[11 : 6])) && (! (1'b1 && (fetch_logic_ctrls_0_down_Fetch_WORD_PC[5 : 3] < FetchL1Plugin_logic_refill_onRsp_wordIndex))))));
  assign fetch_logic_ctrls_0_haltRequest_FetchL1Plugin_l317 = FetchL1Plugin_logic_refill_onRsp_holdHarts;
  assign FetchL1Plugin_logic_bus_rsp_fire = (FetchL1Plugin_logic_bus_rsp_valid && FetchL1Plugin_logic_bus_rsp_ready);
  assign FetchL1Plugin_logic_refill_onRsp_wayToAllocate = FetchL1Plugin_logic_refill_slots_0_wayToAllocate;
  assign FetchL1Plugin_logic_refill_onRsp_address = FetchL1Plugin_logic_refill_slots_0_address;
  assign when_FetchL1Plugin_l324 = (FetchL1Plugin_logic_bus_rsp_valid && (FetchL1Plugin_logic_refill_onRsp_firstCycle || FetchL1Plugin_logic_bus_rsp_payload_error));
  always @(*) begin
    FetchL1Plugin_logic_banks_0_write_valid = (FetchL1Plugin_logic_bus_rsp_valid && (FetchL1Plugin_logic_refill_onRsp_wayToAllocate == 1'b0));
    if(FetchL1Plugin_logic_initializer_busy) begin
      FetchL1Plugin_logic_banks_0_write_valid = 1'b1;
    end
  end

  always @(*) begin
    FetchL1Plugin_logic_banks_0_write_payload_address = {FetchL1Plugin_logic_refill_onRsp_address[11 : 6],FetchL1Plugin_logic_refill_onRsp_wordIndex};
    if(FetchL1Plugin_logic_initializer_busy) begin
      FetchL1Plugin_logic_banks_0_write_payload_address = FetchL1Plugin_logic_initializer_counter[8:0];
    end
  end

  always @(*) begin
    FetchL1Plugin_logic_banks_0_write_payload_data = FetchL1Plugin_logic_bus_rsp_payload_data;
    if(FetchL1Plugin_logic_initializer_busy) begin
      FetchL1Plugin_logic_banks_0_write_payload_data = 64'h0;
    end
  end

  always @(*) begin
    FetchL1Plugin_logic_banks_1_write_valid = (FetchL1Plugin_logic_bus_rsp_valid && (FetchL1Plugin_logic_refill_onRsp_wayToAllocate == 1'b1));
    if(FetchL1Plugin_logic_initializer_busy) begin
      FetchL1Plugin_logic_banks_1_write_valid = 1'b1;
    end
  end

  always @(*) begin
    FetchL1Plugin_logic_banks_1_write_payload_address = {FetchL1Plugin_logic_refill_onRsp_address[11 : 6],FetchL1Plugin_logic_refill_onRsp_wordIndex};
    if(FetchL1Plugin_logic_initializer_busy) begin
      FetchL1Plugin_logic_banks_1_write_payload_address = FetchL1Plugin_logic_initializer_counter[8:0];
    end
  end

  always @(*) begin
    FetchL1Plugin_logic_banks_1_write_payload_data = FetchL1Plugin_logic_bus_rsp_payload_data;
    if(FetchL1Plugin_logic_initializer_busy) begin
      FetchL1Plugin_logic_banks_1_write_payload_data = 64'h0;
    end
  end

  assign FetchL1Plugin_logic_bus_rsp_ready = 1'b1;
  assign when_FetchL1Plugin_l350 = (FetchL1Plugin_logic_refill_onRsp_wordIndex == 3'b111);
  assign FetchL1Plugin_logic_cmd_doIt = (fetch_logic_ctrls_1_up_ready || ((! fetch_logic_ctrls_1_up_valid) && 1'b1));
  assign FetchL1Plugin_logic_banks_0_read_cmd_valid = FetchL1Plugin_logic_cmd_doIt;
  assign FetchL1Plugin_logic_banks_0_read_cmd_payload = fetch_logic_ctrls_0_down_Fetch_WORD_PC[11 : 3];
  assign FetchL1Plugin_logic_banks_1_read_cmd_valid = FetchL1Plugin_logic_cmd_doIt;
  assign FetchL1Plugin_logic_banks_1_read_cmd_payload = fetch_logic_ctrls_0_down_Fetch_WORD_PC[11 : 3];
  assign FetchL1Plugin_logic_ways_0_read_cmd_valid = FetchL1Plugin_logic_cmd_doIt;
  assign FetchL1Plugin_logic_ways_0_read_cmd_payload = fetch_logic_ctrls_0_down_Fetch_WORD_PC[11 : 6];
  assign FetchL1Plugin_logic_ways_1_read_cmd_valid = FetchL1Plugin_logic_cmd_doIt;
  assign FetchL1Plugin_logic_ways_1_read_cmd_payload = fetch_logic_ctrls_0_down_Fetch_WORD_PC[11 : 6];
  assign FetchL1Plugin_logic_plru_read_cmd_valid = FetchL1Plugin_logic_cmd_doIt;
  assign FetchL1Plugin_logic_plru_read_cmd_payload = fetch_logic_ctrls_0_down_Fetch_WORD_PC[11 : 6];
  assign fetch_logic_ctrls_0_down_FetchL1Plugin_logic_cmd_PLRU_BYPASS_VALID = (FetchL1Plugin_logic_plru_write_valid && (FetchL1Plugin_logic_plru_write_payload_address == FetchL1Plugin_logic_plru_read_cmd_payload));
  assign fetch_logic_ctrls_0_down_FetchL1Plugin_logic_cmd_PLRU_BYPASS_DATA_0 = FetchL1Plugin_logic_plru_write_payload_data_0;
  assign fetch_logic_ctrls_0_down_FetchL1Plugin_logic_cmd_TAGS_UPDATE = (|FetchL1Plugin_logic_waysWrite_mask);
  assign fetch_logic_ctrls_0_down_FetchL1Plugin_logic_cmd_TAGS_UPDATE_ADDRESS = FetchL1Plugin_logic_waysWrite_address;
  always @(*) begin
    fetch_logic_ctrls_1_down_FetchL1Plugin_logic_PLRU_BYPASSED_0 = fetch_logic_ctrls_1_down_FetchL1Plugin_logic_PLRU_READ_0;
    if(fetch_logic_ctrls_1_down_FetchL1Plugin_logic_cmd_PLRU_BYPASS_VALID) begin
      fetch_logic_ctrls_1_down_FetchL1Plugin_logic_PLRU_BYPASSED_0 = fetch_logic_ctrls_1_down_FetchL1Plugin_logic_cmd_PLRU_BYPASS_DATA_0;
    end
  end

  assign fetch_logic_ctrls_1_down_FetchL1Plugin_logic_BANKS_MUXES_0 = fetch_logic_ctrls_1_down_FetchL1Plugin_logic_BANKS_WORDS_0[63 : 0];
  assign fetch_logic_ctrls_1_down_FetchL1Plugin_logic_BANKS_MUXES_1 = fetch_logic_ctrls_1_down_FetchL1Plugin_logic_BANKS_WORDS_1[63 : 0];
  assign fetch_logic_ctrls_2_down_Fetch_WORD = ((fetch_logic_ctrls_2_down_FetchL1Plugin_logic_WAYS_HITS_0 ? fetch_logic_ctrls_2_down_FetchL1Plugin_logic_BANKS_MUXES_0 : 64'h0) | (fetch_logic_ctrls_2_down_FetchL1Plugin_logic_WAYS_HITS_1 ? fetch_logic_ctrls_2_down_FetchL1Plugin_logic_BANKS_MUXES_1 : 64'h0));
  assign fetch_logic_ctrls_1_down_FetchL1Plugin_logic_HAZARD = (fetch_logic_ctrls_1_down_FetchL1Plugin_logic_cmd_TAGS_UPDATE && (fetch_logic_ctrls_1_down_FetchL1Plugin_logic_cmd_TAGS_UPDATE_ADDRESS == fetch_logic_ctrls_1_down_Fetch_WORD_PC[11 : 6]));
  assign FetchL1Plugin_logic_hits_w_0_indirect_wayTlbHits_0 = ((fetch_logic_ctrls_1_down_FetchL1Plugin_logic_WAYS_TAGS_0_address == fetch_logic_ctrls_1_down_MMU_WAYS_PHYSICAL_0[31 : 12]) && fetch_logic_ctrls_1_down_MMU_WAYS_OH[0]);
  assign FetchL1Plugin_logic_hits_w_0_indirect_wayTlbHits_1 = ((fetch_logic_ctrls_1_down_FetchL1Plugin_logic_WAYS_TAGS_0_address == fetch_logic_ctrls_1_down_MMU_WAYS_PHYSICAL_1[31 : 12]) && fetch_logic_ctrls_1_down_MMU_WAYS_OH[1]);
  assign FetchL1Plugin_logic_hits_w_0_indirect_wayTlbHits_2 = ((fetch_logic_ctrls_1_down_FetchL1Plugin_logic_WAYS_TAGS_0_address == fetch_logic_ctrls_1_down_MMU_WAYS_PHYSICAL_2[31 : 12]) && fetch_logic_ctrls_1_down_MMU_WAYS_OH[2]);
  assign FetchL1Plugin_logic_hits_w_0_indirect_translatedHits = (|{FetchL1Plugin_logic_hits_w_0_indirect_wayTlbHits_2,{FetchL1Plugin_logic_hits_w_0_indirect_wayTlbHits_1,FetchL1Plugin_logic_hits_w_0_indirect_wayTlbHits_0}});
  assign FetchL1Plugin_logic_hits_w_0_indirect_bypassHits = (fetch_logic_ctrls_1_down_FetchL1Plugin_logic_WAYS_TAGS_0_address == _zz_FetchL1Plugin_logic_hits_w_0_indirect_bypassHits);
  assign fetch_logic_ctrls_1_down_FetchL1Plugin_logic_WAYS_HITS_0 = ((fetch_logic_ctrls_1_down_MMU_BYPASS_TRANSLATION ? FetchL1Plugin_logic_hits_w_0_indirect_bypassHits : FetchL1Plugin_logic_hits_w_0_indirect_translatedHits) && fetch_logic_ctrls_1_down_FetchL1Plugin_logic_WAYS_TAGS_0_loaded);
  assign FetchL1Plugin_logic_hits_w_1_indirect_wayTlbHits_0 = ((fetch_logic_ctrls_1_down_FetchL1Plugin_logic_WAYS_TAGS_1_address == fetch_logic_ctrls_1_down_MMU_WAYS_PHYSICAL_0[31 : 12]) && fetch_logic_ctrls_1_down_MMU_WAYS_OH[0]);
  assign FetchL1Plugin_logic_hits_w_1_indirect_wayTlbHits_1 = ((fetch_logic_ctrls_1_down_FetchL1Plugin_logic_WAYS_TAGS_1_address == fetch_logic_ctrls_1_down_MMU_WAYS_PHYSICAL_1[31 : 12]) && fetch_logic_ctrls_1_down_MMU_WAYS_OH[1]);
  assign FetchL1Plugin_logic_hits_w_1_indirect_wayTlbHits_2 = ((fetch_logic_ctrls_1_down_FetchL1Plugin_logic_WAYS_TAGS_1_address == fetch_logic_ctrls_1_down_MMU_WAYS_PHYSICAL_2[31 : 12]) && fetch_logic_ctrls_1_down_MMU_WAYS_OH[2]);
  assign FetchL1Plugin_logic_hits_w_1_indirect_translatedHits = (|{FetchL1Plugin_logic_hits_w_1_indirect_wayTlbHits_2,{FetchL1Plugin_logic_hits_w_1_indirect_wayTlbHits_1,FetchL1Plugin_logic_hits_w_1_indirect_wayTlbHits_0}});
  assign FetchL1Plugin_logic_hits_w_1_indirect_bypassHits = (fetch_logic_ctrls_1_down_FetchL1Plugin_logic_WAYS_TAGS_1_address == _zz_FetchL1Plugin_logic_hits_w_1_indirect_bypassHits);
  assign fetch_logic_ctrls_1_down_FetchL1Plugin_logic_WAYS_HITS_1 = ((fetch_logic_ctrls_1_down_MMU_BYPASS_TRANSLATION ? FetchL1Plugin_logic_hits_w_1_indirect_bypassHits : FetchL1Plugin_logic_hits_w_1_indirect_translatedHits) && fetch_logic_ctrls_1_down_FetchL1Plugin_logic_WAYS_TAGS_1_loaded);
  assign fetch_logic_ctrls_1_down_FetchL1Plugin_logic_WAYS_HIT = (|{fetch_logic_ctrls_1_down_FetchL1Plugin_logic_WAYS_HITS_1,fetch_logic_ctrls_1_down_FetchL1Plugin_logic_WAYS_HITS_0});
  assign FetchL1Plugin_logic_ctrl_pmaPort_cmd_address = fetch_logic_ctrls_2_down_MMU_TRANSLATED;
  assign FetchL1Plugin_logic_ctrl_plruLogic_core_evict_logic_0_state = FetchL1Plugin_logic_ctrl_plruLogic_core_io_context_state_0[0];
  assign FetchL1Plugin_logic_ctrl_plruLogic_core_evict_sel_0 = (! FetchL1Plugin_logic_ctrl_plruLogic_core_evict_logic_0_state);
  assign FetchL1Plugin_logic_ctrl_plruLogic_core_io_evict_id = FetchL1Plugin_logic_ctrl_plruLogic_core_evict_sel_0;
  assign FetchL1Plugin_logic_ctrl_plruLogic_core_io_update_state_0[0] = FetchL1Plugin_logic_ctrl_plruLogic_core_io_update_id[0];
  assign FetchL1Plugin_logic_ctrl_plruLogic_core_io_context_state_0 = fetch_logic_ctrls_2_down_FetchL1Plugin_logic_PLRU_BYPASSED_0;
  assign FetchL1Plugin_logic_ctrl_plruLogic_core_io_update_id = fetch_logic_ctrls_2_down_FetchL1Plugin_logic_WAYS_HITS_1;
  always @(*) begin
    FetchL1Plugin_logic_plru_write_valid = FetchL1Plugin_logic_ctrl_plruLogic_buffer_regNext_valid;
    if(when_FetchL1Plugin_l567) begin
      FetchL1Plugin_logic_plru_write_valid = 1'b1;
    end
  end

  always @(*) begin
    FetchL1Plugin_logic_plru_write_payload_address = FetchL1Plugin_logic_ctrl_plruLogic_buffer_regNext_payload_address;
    if(when_FetchL1Plugin_l567) begin
      FetchL1Plugin_logic_plru_write_payload_address = FetchL1Plugin_logic_invalidate_counter[5:0];
    end
  end

  always @(*) begin
    FetchL1Plugin_logic_plru_write_payload_data_0 = FetchL1Plugin_logic_ctrl_plruLogic_buffer_regNext_payload_data_0;
    if(when_FetchL1Plugin_l567) begin
      FetchL1Plugin_logic_plru_write_payload_data_0 = _zz_FetchL1Plugin_logic_plru_write_payload_data_0[0 : 0];
    end
  end

  assign FetchL1Plugin_logic_ctrl_plruLogic_buffer_valid = (fetch_logic_ctrls_2_up_isValid && fetch_logic_ctrls_2_up_isReady);
  assign FetchL1Plugin_logic_ctrl_plruLogic_buffer_payload_address = fetch_logic_ctrls_2_down_Fetch_WORD_PC[11 : 6];
  assign FetchL1Plugin_logic_ctrl_plruLogic_buffer_payload_data_0 = FetchL1Plugin_logic_ctrl_plruLogic_core_io_update_state_0;
  assign FetchL1Plugin_logic_refill_start_wayToAllocate = FetchL1Plugin_logic_ctrl_plruLogic_core_io_evict_id;
  assign FetchL1Plugin_logic_ctrl_dataAccessFault = (_zz_FetchL1Plugin_logic_ctrl_dataAccessFault[0] && (! fetch_logic_ctrls_2_down_FetchL1Plugin_logic_HAZARD));
  always @(*) begin
    FetchL1Plugin_logic_trapPort_valid = 1'b0;
    if(when_FetchL1Plugin_l483) begin
      FetchL1Plugin_logic_trapPort_valid = 1'b1;
    end
    if(when_FetchL1Plugin_l489) begin
      FetchL1Plugin_logic_trapPort_valid = 1'b1;
    end
    if(when_FetchL1Plugin_l496) begin
      FetchL1Plugin_logic_trapPort_valid = 1'b1;
    end
    if(fetch_logic_ctrls_2_down_MMU_ACCESS_FAULT) begin
      FetchL1Plugin_logic_trapPort_valid = 1'b1;
    end
    if(fetch_logic_ctrls_2_down_MMU_REFILL) begin
      FetchL1Plugin_logic_trapPort_valid = 1'b1;
    end
    if(fetch_logic_ctrls_2_down_MMU_HAZARD) begin
      FetchL1Plugin_logic_trapPort_valid = 1'b1;
    end
    if(fetch_logic_ctrls_2_down_Fetch_PC_FAULT) begin
      FetchL1Plugin_logic_trapPort_valid = 1'b1;
    end
    if(when_FetchL1Plugin_l542) begin
      FetchL1Plugin_logic_trapPort_valid = 1'b0;
    end
  end

  assign FetchL1Plugin_logic_trapPort_payload_tval = fetch_logic_ctrls_2_down_Fetch_WORD_PC;
  always @(*) begin
    FetchL1Plugin_logic_trapPort_payload_exception = 1'bx;
    if(when_FetchL1Plugin_l483) begin
      FetchL1Plugin_logic_trapPort_payload_exception = 1'b0;
    end
    if(when_FetchL1Plugin_l489) begin
      FetchL1Plugin_logic_trapPort_payload_exception = 1'b1;
    end
    if(when_FetchL1Plugin_l496) begin
      FetchL1Plugin_logic_trapPort_payload_exception = 1'b1;
    end
    if(fetch_logic_ctrls_2_down_MMU_ACCESS_FAULT) begin
      FetchL1Plugin_logic_trapPort_payload_exception = 1'b1;
    end
    if(fetch_logic_ctrls_2_down_MMU_REFILL) begin
      FetchL1Plugin_logic_trapPort_payload_exception = 1'b0;
    end
    if(fetch_logic_ctrls_2_down_MMU_HAZARD) begin
      FetchL1Plugin_logic_trapPort_payload_exception = 1'b0;
    end
    if(fetch_logic_ctrls_2_down_Fetch_PC_FAULT) begin
      FetchL1Plugin_logic_trapPort_payload_exception = 1'b1;
    end
  end

  always @(*) begin
    FetchL1Plugin_logic_trapPort_payload_code = 4'bxxxx;
    if(when_FetchL1Plugin_l483) begin
      FetchL1Plugin_logic_trapPort_payload_code = 4'b0100;
    end
    if(when_FetchL1Plugin_l489) begin
      FetchL1Plugin_logic_trapPort_payload_code = 4'b0001;
    end
    if(when_FetchL1Plugin_l496) begin
      FetchL1Plugin_logic_trapPort_payload_code = 4'b1100;
    end
    if(fetch_logic_ctrls_2_down_MMU_ACCESS_FAULT) begin
      FetchL1Plugin_logic_trapPort_payload_code = 4'b0001;
    end
    if(fetch_logic_ctrls_2_down_MMU_REFILL) begin
      FetchL1Plugin_logic_trapPort_payload_code = 4'b0111;
    end
    if(fetch_logic_ctrls_2_down_MMU_HAZARD) begin
      FetchL1Plugin_logic_trapPort_payload_code = 4'b0100;
    end
    if(fetch_logic_ctrls_2_down_Fetch_PC_FAULT) begin
      FetchL1Plugin_logic_trapPort_payload_code = 4'b0001;
      if(when_FetchL1Plugin_l529) begin
        FetchL1Plugin_logic_trapPort_payload_code = 4'b1100;
      end
    end
  end

  assign _zz_59 = zz_FetchL1Plugin_logic_trapPort_payload_arg(1'b0);
  always @(*) FetchL1Plugin_logic_trapPort_payload_arg = _zz_59;
  always @(*) begin
    FetchL1Plugin_logic_ctrl_allowRefill = ((! fetch_logic_ctrls_2_down_FetchL1Plugin_logic_WAYS_HIT) && (! fetch_logic_ctrls_2_down_FetchL1Plugin_logic_HAZARD));
    if(when_FetchL1Plugin_l489) begin
      FetchL1Plugin_logic_ctrl_allowRefill = 1'b0;
    end
    if(when_FetchL1Plugin_l496) begin
      FetchL1Plugin_logic_ctrl_allowRefill = 1'b0;
    end
    if(fetch_logic_ctrls_2_down_MMU_ACCESS_FAULT) begin
      FetchL1Plugin_logic_ctrl_allowRefill = 1'b0;
    end
    if(fetch_logic_ctrls_2_down_MMU_REFILL) begin
      FetchL1Plugin_logic_ctrl_allowRefill = 1'b0;
    end
    if(fetch_logic_ctrls_2_down_MMU_HAZARD) begin
      FetchL1Plugin_logic_ctrl_allowRefill = 1'b0;
    end
    if(fetch_logic_ctrls_2_down_Fetch_PC_FAULT) begin
      FetchL1Plugin_logic_ctrl_allowRefill = 1'b0;
    end
  end

  assign when_FetchL1Plugin_l483 = ((! fetch_logic_ctrls_2_down_FetchL1Plugin_logic_WAYS_HIT) || fetch_logic_ctrls_2_down_FetchL1Plugin_logic_HAZARD);
  assign when_FetchL1Plugin_l489 = (FetchL1Plugin_logic_ctrl_dataAccessFault || FetchL1Plugin_logic_ctrl_pmaPort_rsp_fault);
  assign when_FetchL1Plugin_l496 = (fetch_logic_ctrls_2_down_MMU_PAGE_FAULT || (! fetch_logic_ctrls_2_down_MMU_ALLOW_EXECUTE));
  assign when_FetchL1Plugin_l529 = (! fetch_logic_ctrls_2_down_MMU_BYPASS_TRANSLATION);
  always @(*) begin
    FetchL1Plugin_logic_refill_start_valid = (FetchL1Plugin_logic_ctrl_allowRefill && (! FetchL1Plugin_logic_ctrl_trapSent));
    if(when_FetchL1Plugin_l546) begin
      FetchL1Plugin_logic_refill_start_valid = 1'b0;
    end
  end

  assign FetchL1Plugin_logic_refill_start_address = fetch_logic_ctrls_2_down_MMU_TRANSLATED;
  assign FetchL1Plugin_logic_refill_start_isIo = FetchL1Plugin_logic_ctrl_pmaPort_rsp_io;
  assign fetch_logic_ctrls_2_down_TRAP = (FetchL1Plugin_logic_trapPort_valid || FetchL1Plugin_logic_ctrl_trapSent);
  assign when_FetchL1Plugin_l542 = ((! fetch_logic_ctrls_2_up_isValid) || FetchL1Plugin_logic_ctrl_trapSent);
  assign when_FetchL1Plugin_l546 = ((! fetch_logic_ctrls_2_up_isValid) && 1'b1);
  assign when_FetchL1Plugin_l550 = (((! fetch_logic_ctrls_2_up_isValid) || fetch_logic_ctrls_2_down_isReady) || fetch_logic_ctrls_2_up_isCanceling);
  assign when_FetchL1Plugin_l567 = (! FetchL1Plugin_logic_invalidate_done);
  assign FetchL1Plugin_logic_initializer_busy = (! FetchL1Plugin_logic_initializer_counter[9]);
  assign toplevel_execute_ctrl0_down_AguPlugin_SIZE_lane0 = toplevel_execute_ctrl0_down_Decode_UOP_lane0[13 : 12];
  assign LsuPlugin_logic_flusher_wantExit = 1'b0;
  always @(*) begin
    LsuPlugin_logic_flusher_wantStart = 1'b0;
    case(LsuPlugin_logic_flusher_stateReg)
      LsuPlugin_logic_flusher_enumDef_CMD : begin
      end
      LsuPlugin_logic_flusher_enumDef_COMPLETION : begin
      end
      default : begin
        LsuPlugin_logic_flusher_wantStart = 1'b1;
      end
    endcase
  end

  assign LsuPlugin_logic_flusher_wantKill = 1'b0;
  assign TrapPlugin_logic_lsuL1Invalidate_0_cmd_ready = LsuPlugin_logic_flusher_arbiter_io_inputs_0_ready;
  assign LsuPlugin_logic_flusher_inflight = (|{(toplevel_execute_ctrl4_down_LsuL1_SEL_lane0 && toplevel_execute_ctrl4_down_LsuL1_FLUSH_lane0),(toplevel_execute_ctrl3_down_LsuL1_SEL_lane0 && toplevel_execute_ctrl3_down_LsuL1_FLUSH_lane0)});
  always @(*) begin
    PrivilegedPlugin_logic_harts_0_xretAwayFromMachine = 1'b0;
    case(TrapPlugin_logic_harts_0_trap_fsm_stateReg)
      TrapPlugin_logic_harts_0_trap_fsm_enumDef_RUNNING : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_enumDef_PROCESS_1 : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_enumDef_TRAP_EPC : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_enumDef_TRAP_TVAL : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_enumDef_TRAP_TVEC : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_enumDef_TRAP_APPLY : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_enumDef_XRET_EPC : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_enumDef_XRET_APPLY : begin
        if(when_TrapPlugin_l637) begin
          PrivilegedPlugin_logic_harts_0_xretAwayFromMachine = 1'b1;
        end
      end
      TrapPlugin_logic_harts_0_trap_fsm_enumDef_ATS_RSP : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_enumDef_JUMP : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_enumDef_LSU_FLUSH : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_enumDef_FETCH_FLUSH : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    PrivilegedPlugin_logic_harts_0_int_pending = 1'b0;
    if(TrapPlugin_logic_harts_0_interrupt_pendingInterrupt) begin
      PrivilegedPlugin_logic_harts_0_int_pending = 1'b1;
    end
  end

  assign PrivilegedPlugin_logic_harts_0_withMachinePrivilege = (2'b11 <= PrivilegedPlugin_logic_harts_0_privilege);
  assign PrivilegedPlugin_logic_harts_0_withSupervisorPrivilege = (2'b01 <= PrivilegedPlugin_logic_harts_0_privilege);
  assign PrivilegedPlugin_logic_harts_0_hartRunning = 1'b1;
  assign PrivilegedPlugin_logic_harts_0_debugMode = (! PrivilegedPlugin_logic_harts_0_hartRunning);
  always @(*) begin
    PrivilegedPlugin_logic_harts_0_m_status_sd = 1'b0;
    if(when_PrivilegedPlugin_l533) begin
      PrivilegedPlugin_logic_harts_0_m_status_sd = 1'b1;
    end
  end

  assign when_PrivilegedPlugin_l533 = (PrivilegedPlugin_logic_harts_0_m_status_fs == 2'b11);
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_1 = (when_CsrService_l188 && _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue);
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_2 = (when_CsrService_l188 && REG_CSR_834);
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_3 = (when_CsrService_l188 && REG_CSR_836);
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_4 = (when_CsrService_l188 && REG_CSR_772);
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_5 = (when_CsrService_l188 && REG_CSR_770);
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_6 = (when_CsrService_l188 && REG_CSR_771);
  assign _zz_when_TrapPlugin_l195 = (PrivilegedPlugin_logic_harts_0_m_ip_mtip && PrivilegedPlugin_logic_harts_0_m_ie_mtie);
  assign _zz_when_TrapPlugin_l195_1 = (PrivilegedPlugin_logic_harts_0_m_ip_msip && PrivilegedPlugin_logic_harts_0_m_ie_msie);
  assign _zz_when_TrapPlugin_l195_2 = (PrivilegedPlugin_logic_harts_0_m_ip_meip && PrivilegedPlugin_logic_harts_0_m_ie_meie);
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_7 = (when_CsrService_l188 && REG_CSR_322);
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_9 = (when_CsrService_l188 && _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_8);
  assign PrivilegedPlugin_logic_harts_0_s_ip_seipOr = (PrivilegedPlugin_logic_harts_0_s_ip_seipSoft || PrivilegedPlugin_logic_harts_0_s_ip_seipInput);
  assign PrivilegedPlugin_logic_harts_0_s_ip_seipMasked = (PrivilegedPlugin_logic_harts_0_s_ip_seipOr && PrivilegedPlugin_logic_harts_0_m_ideleg_se);
  assign PrivilegedPlugin_logic_harts_0_s_ip_stipMasked = (PrivilegedPlugin_logic_harts_0_s_ip_stip && PrivilegedPlugin_logic_harts_0_m_ideleg_st);
  assign PrivilegedPlugin_logic_harts_0_s_ip_ssipMasked = (PrivilegedPlugin_logic_harts_0_s_ip_ssip && PrivilegedPlugin_logic_harts_0_m_ideleg_ss);
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_10 = (when_CsrService_l188 && REG_CSR_260);
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_11 = (when_CsrService_l188 && REG_CSR_324);
  assign _zz_when_TrapPlugin_l195_3 = (PrivilegedPlugin_logic_harts_0_s_ip_ssip && PrivilegedPlugin_logic_harts_0_s_ie_ssie);
  assign _zz_when_TrapPlugin_l195_4 = (PrivilegedPlugin_logic_harts_0_s_ip_stip && PrivilegedPlugin_logic_harts_0_s_ie_stie);
  assign _zz_when_TrapPlugin_l195_5 = (PrivilegedPlugin_logic_harts_0_s_ip_seipOr && PrivilegedPlugin_logic_harts_0_s_ie_seie);
  assign PrivilegedPlugin_logic_defaultTrap_csrPrivilege = CsrAccessPlugin_bus_decode_address[9 : 8];
  assign PrivilegedPlugin_logic_defaultTrap_csrReadOnly = (CsrAccessPlugin_bus_decode_address[11 : 10] == 2'b11);
  assign when_PrivilegedPlugin_l679 = ((PrivilegedPlugin_logic_defaultTrap_csrReadOnly && CsrAccessPlugin_bus_decode_write) || (PrivilegedPlugin_logic_harts_0_privilege < PrivilegedPlugin_logic_defaultTrap_csrPrivilege));
  assign _zz_fetch_logic_ctrls_0_down_GSharePlugin_logic_HASH = fetch_logic_ctrls_0_down_Fetch_WORD_PC[14 : 3];
  assign fetch_logic_ctrls_0_down_GSharePlugin_logic_HASH = ({_zz_fetch_logic_ctrls_0_down_GSharePlugin_logic_HASH[0],{_zz_fetch_logic_ctrls_0_down_GSharePlugin_logic_HASH[1],{_zz_fetch_logic_ctrls_0_down_GSharePlugin_logic_HASH[2],{_zz_fetch_logic_ctrls_0_down_GSharePlugin_logic_HASH[3],{_zz_fetch_logic_ctrls_0_down_GSharePlugin_logic_HASH[4],{_zz_fetch_logic_ctrls_0_down_GSharePlugin_logic_HASH[5],{_zz_fetch_logic_ctrls_0_down_GSharePlugin_logic_HASH_1,{_zz_fetch_logic_ctrls_0_down_GSharePlugin_logic_HASH_2,_zz_fetch_logic_ctrls_0_down_GSharePlugin_logic_HASH_3}}}}}}}} ^ fetch_logic_ctrls_0_down_Prediction_BRANCH_HISTORY);
  assign fetch_logic_ctrls_0_down_GSharePlugin_logic_BYPASS_valid = GSharePlugin_logic_mem_write_valid;
  assign fetch_logic_ctrls_0_down_GSharePlugin_logic_BYPASS_payload_address = GSharePlugin_logic_mem_write_payload_address;
  assign fetch_logic_ctrls_0_down_GSharePlugin_logic_BYPASS_payload_data_0 = GSharePlugin_logic_mem_write_payload_data_0;
  assign fetch_logic_ctrls_0_down_GSharePlugin_logic_BYPASS_payload_data_1 = GSharePlugin_logic_mem_write_payload_data_1;
  assign fetch_logic_ctrls_0_down_GSharePlugin_logic_BYPASS_payload_data_2 = GSharePlugin_logic_mem_write_payload_data_2;
  assign fetch_logic_ctrls_0_down_GSharePlugin_logic_BYPASS_payload_data_3 = GSharePlugin_logic_mem_write_payload_data_3;
  assign _zz_fetch_logic_ctrls_1_down_GSharePlugin_GSHARE_COUNTER_0 = GSharePlugin_logic_mem_counter_spinal_port1;
  always @(*) begin
    fetch_logic_ctrls_1_down_GSharePlugin_GSHARE_COUNTER_0 = _zz_fetch_logic_ctrls_1_down_GSharePlugin_GSHARE_COUNTER_0[1 : 0];
    if(when_GSharePlugin_l82) begin
      fetch_logic_ctrls_1_down_GSharePlugin_GSHARE_COUNTER_0 = fetch_logic_ctrls_1_down_GSharePlugin_logic_BYPASS_payload_data_0;
    end
  end

  always @(*) begin
    fetch_logic_ctrls_1_down_GSharePlugin_GSHARE_COUNTER_1 = _zz_fetch_logic_ctrls_1_down_GSharePlugin_GSHARE_COUNTER_0[3 : 2];
    if(when_GSharePlugin_l82) begin
      fetch_logic_ctrls_1_down_GSharePlugin_GSHARE_COUNTER_1 = fetch_logic_ctrls_1_down_GSharePlugin_logic_BYPASS_payload_data_1;
    end
  end

  always @(*) begin
    fetch_logic_ctrls_1_down_GSharePlugin_GSHARE_COUNTER_2 = _zz_fetch_logic_ctrls_1_down_GSharePlugin_GSHARE_COUNTER_0[5 : 4];
    if(when_GSharePlugin_l82) begin
      fetch_logic_ctrls_1_down_GSharePlugin_GSHARE_COUNTER_2 = fetch_logic_ctrls_1_down_GSharePlugin_logic_BYPASS_payload_data_2;
    end
  end

  always @(*) begin
    fetch_logic_ctrls_1_down_GSharePlugin_GSHARE_COUNTER_3 = _zz_fetch_logic_ctrls_1_down_GSharePlugin_GSHARE_COUNTER_0[7 : 6];
    if(when_GSharePlugin_l82) begin
      fetch_logic_ctrls_1_down_GSharePlugin_GSHARE_COUNTER_3 = fetch_logic_ctrls_1_down_GSharePlugin_logic_BYPASS_payload_data_3;
    end
  end

  assign when_GSharePlugin_l82 = (fetch_logic_ctrls_1_down_GSharePlugin_logic_BYPASS_valid && (fetch_logic_ctrls_1_down_GSharePlugin_logic_BYPASS_payload_address == fetch_logic_ctrls_1_down_GSharePlugin_logic_HASH));
  always @(*) begin
    BtbPlugin_logic_ras_ptr_pushIt = 1'b0;
    if(BtbPlugin_logic_applyIt_rasLogic_pushValid) begin
      BtbPlugin_logic_ras_ptr_pushIt = 1'b1;
    end
  end

  always @(*) begin
    BtbPlugin_logic_ras_ptr_popIt = 1'b0;
    if(when_BtbPlugin_l218) begin
      BtbPlugin_logic_ras_ptr_popIt = 1'b1;
    end
  end

  always @(*) begin
    BtbPlugin_logic_ras_write_valid = BtbPlugin_logic_ras_ptr_pushIt;
    if(BtbPlugin_logic_initializer_busy) begin
      BtbPlugin_logic_ras_write_valid = 1'b1;
    end
  end

  always @(*) begin
    BtbPlugin_logic_ras_write_payload_address = BtbPlugin_logic_ras_ptr_push;
    if(BtbPlugin_logic_initializer_busy) begin
      BtbPlugin_logic_ras_write_payload_address = BtbPlugin_logic_initializer_counter[1:0];
    end
  end

  always @(*) begin
    BtbPlugin_logic_ras_write_payload_data = 31'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
    BtbPlugin_logic_ras_write_payload_data = (_zz_BtbPlugin_logic_ras_write_payload_data >>> 1'd1);
    if(BtbPlugin_logic_initializer_busy) begin
      BtbPlugin_logic_ras_write_payload_data = 31'h0;
    end
  end

  assign WhiteboxerPlugin_logic_fetch_fetchId = fetch_logic_ctrls_0_down_Fetch_ID;
  assign WhiteboxerPlugin_logic_decodes_0_fire = ((toplevel_decode_ctrls_0_up_LANE_SEL_0 && toplevel_decode_ctrls_0_up_isReady) && (! toplevel_decode_ctrls_0_lane0_upIsCancel));
  assign when_CtrlLaneApi_l46 = (toplevel_decode_ctrls_0_up_isReady || toplevel_decode_ctrls_0_lane0_upIsCancel);
  assign WhiteboxerPlugin_logic_decodes_0_spawn = (toplevel_decode_ctrls_0_up_LANE_SEL_0 && (! toplevel_decode_ctrls_0_up_LANE_SEL_0_regNext));
  assign WhiteboxerPlugin_logic_decodes_0_pc = _zz_WhiteboxerPlugin_logic_decodes_0_pc;
  assign WhiteboxerPlugin_logic_decodes_0_fetchId = toplevel_decode_ctrls_0_down_Fetch_ID_0;
  assign WhiteboxerPlugin_logic_decodes_0_decodeId = toplevel_decode_ctrls_0_down_Decode_DOP_ID_0;
  assign WhiteboxerPlugin_logic_decodes_1_fire = ((toplevel_decode_ctrls_0_up_LANE_SEL_1 && toplevel_decode_ctrls_0_up_isReady) && (! toplevel_decode_ctrls_0_lane1_upIsCancel));
  assign when_CtrlLaneApi_l46_1 = (toplevel_decode_ctrls_0_up_isReady || toplevel_decode_ctrls_0_lane1_upIsCancel);
  assign WhiteboxerPlugin_logic_decodes_1_spawn = (toplevel_decode_ctrls_0_up_LANE_SEL_1 && (! toplevel_decode_ctrls_0_up_LANE_SEL_1_regNext));
  assign WhiteboxerPlugin_logic_decodes_1_pc = _zz_WhiteboxerPlugin_logic_decodes_1_pc;
  assign WhiteboxerPlugin_logic_decodes_1_fetchId = toplevel_decode_ctrls_0_down_Fetch_ID_1;
  assign WhiteboxerPlugin_logic_decodes_1_decodeId = toplevel_decode_ctrls_0_down_Decode_DOP_ID_1;
  assign toplevel_execute_ctrl2_down_early0_BranchPlugin_logic_alu_EQ_lane0 = ($signed(toplevel_execute_ctrl2_down_early0_SrcPlugin_SRC1_lane0) == $signed(toplevel_execute_ctrl2_down_early0_SrcPlugin_SRC2_lane0));
  assign toplevel_execute_ctrl2_down_early0_BranchPlugin_logic_alu_btb_BAD_TARGET_lane0 = (toplevel_execute_ctrl2_down_Prediction_ALIGNED_JUMPED_PC_lane0 != toplevel_execute_ctrl2_down_early0_BranchPlugin_pcCalc_PC_TRUE_lane0);
  assign early0_BranchPlugin_logic_alu_expectedMsb = (MmuPlugin_api_fetchTranslationEnable ? _zz_early0_BranchPlugin_logic_alu_expectedMsb[31] : 1'b0);
  assign toplevel_execute_ctrl2_down_early0_BranchPlugin_logic_alu_MSB_FAILED_lane0 = ((toplevel_execute_ctrl2_down_BranchPlugin_BRANCH_CTRL_lane0 == BranchPlugin_BranchCtrlEnum_JALR) && 1'b0);
  assign switch_Misc_l241 = toplevel_execute_ctrl3_down_Decode_UOP_lane0[14 : 12];
  always @(*) begin
    casez(switch_Misc_l241)
      3'b000 : begin
        _zz_toplevel_execute_ctrl3_down_early0_BranchPlugin_logic_jumpLogic_COND_lane0 = toplevel_execute_ctrl3_down_early0_BranchPlugin_logic_alu_EQ_lane0;
      end
      3'b001 : begin
        _zz_toplevel_execute_ctrl3_down_early0_BranchPlugin_logic_jumpLogic_COND_lane0 = (! toplevel_execute_ctrl3_down_early0_BranchPlugin_logic_alu_EQ_lane0);
      end
      3'b1?1 : begin
        _zz_toplevel_execute_ctrl3_down_early0_BranchPlugin_logic_jumpLogic_COND_lane0 = (! toplevel_execute_ctrl3_down_early0_SrcPlugin_LESS_lane0);
      end
      default : begin
        _zz_toplevel_execute_ctrl3_down_early0_BranchPlugin_logic_jumpLogic_COND_lane0 = toplevel_execute_ctrl3_down_early0_SrcPlugin_LESS_lane0;
      end
    endcase
  end

  always @(*) begin
    case(toplevel_execute_ctrl3_down_BranchPlugin_BRANCH_CTRL_lane0)
      BranchPlugin_BranchCtrlEnum_JALR : begin
        _zz_toplevel_execute_ctrl3_down_early0_BranchPlugin_logic_jumpLogic_COND_lane0_1 = 1'b1;
      end
      BranchPlugin_BranchCtrlEnum_JAL : begin
        _zz_toplevel_execute_ctrl3_down_early0_BranchPlugin_logic_jumpLogic_COND_lane0_1 = 1'b1;
      end
      default : begin
        _zz_toplevel_execute_ctrl3_down_early0_BranchPlugin_logic_jumpLogic_COND_lane0_1 = _zz_toplevel_execute_ctrl3_down_early0_BranchPlugin_logic_jumpLogic_COND_lane0;
      end
    endcase
  end

  assign toplevel_execute_ctrl3_down_early0_BranchPlugin_logic_jumpLogic_COND_lane0 = _zz_toplevel_execute_ctrl3_down_early0_BranchPlugin_logic_jumpLogic_COND_lane0_1;
  assign toplevel_execute_ctrl3_down_early0_BranchPlugin_logic_jumpLogic_btb_REAL_TARGET_lane0 = (toplevel_execute_ctrl3_down_early0_BranchPlugin_logic_jumpLogic_COND_lane0 ? toplevel_execute_ctrl3_down_early0_BranchPlugin_pcCalc_PC_TRUE_lane0 : toplevel_execute_ctrl3_down_early0_BranchPlugin_pcCalc_PC_FALSE_lane0);
  assign early0_BranchPlugin_logic_jumpLogic_wrongCond = (toplevel_execute_ctrl3_down_Prediction_ALIGNED_JUMPED_lane0 != toplevel_execute_ctrl3_down_early0_BranchPlugin_logic_jumpLogic_COND_lane0);
  assign early0_BranchPlugin_logic_jumpLogic_needFix = ((early0_BranchPlugin_logic_jumpLogic_wrongCond || (toplevel_execute_ctrl3_down_early0_BranchPlugin_logic_jumpLogic_COND_lane0 && toplevel_execute_ctrl3_down_early0_BranchPlugin_logic_alu_btb_BAD_TARGET_lane0)) || toplevel_execute_ctrl3_down_early0_BranchPlugin_logic_alu_MSB_FAILED_lane0);
  assign early0_BranchPlugin_logic_jumpLogic_doIt = ((toplevel_execute_ctrl3_up_LANE_SEL_lane0 && toplevel_execute_ctrl3_down_early0_BranchPlugin_SEL_lane0) && early0_BranchPlugin_logic_jumpLogic_needFix);
  assign early0_BranchPlugin_logic_jumpLogic_history_fromFetch_slice = toplevel_execute_ctrl3_down_PC_lane0[2 : 1];
  assign early0_BranchPlugin_logic_jumpLogic_history_fromFetch_shifter = toplevel_execute_ctrl3_down_Prediction_BRANCH_HISTORY_lane0;
  assign when_BranchPlugin_l206 = ((early0_BranchPlugin_logic_jumpLogic_history_fromFetch_slice < 2'b00) && toplevel_execute_ctrl3_down_Prediction_ALIGNED_SLICES_BRANCH_lane0[0]);
  assign when_BranchPlugin_l206_1 = ((early0_BranchPlugin_logic_jumpLogic_history_fromFetch_slice < 2'b01) && toplevel_execute_ctrl3_down_Prediction_ALIGNED_SLICES_BRANCH_lane0[1]);
  assign when_BranchPlugin_l206_2 = ((early0_BranchPlugin_logic_jumpLogic_history_fromFetch_slice < 2'b10) && toplevel_execute_ctrl3_down_Prediction_ALIGNED_SLICES_BRANCH_lane0[2]);
  assign when_BranchPlugin_l210 = (toplevel_execute_ctrl3_down_BranchPlugin_BRANCH_CTRL_lane0 == BranchPlugin_BranchCtrlEnum_B);
  assign early0_BranchPlugin_logic_jumpLogic_history_next = early0_BranchPlugin_logic_jumpLogic_history_fromFetch_shifter_4;
  assign early0_BranchPlugin_logic_jumpLogic_history_fetched = toplevel_execute_ctrl3_down_Prediction_BRANCH_HISTORY_lane0;
  assign early0_BranchPlugin_logic_pcPort_valid = early0_BranchPlugin_logic_jumpLogic_doIt;
  assign early0_BranchPlugin_logic_pcPort_payload_fault = toplevel_execute_ctrl3_down_early0_BranchPlugin_logic_alu_MSB_FAILED_lane0;
  assign early0_BranchPlugin_logic_pcPort_payload_pc = toplevel_execute_ctrl3_down_early0_BranchPlugin_logic_jumpLogic_btb_REAL_TARGET_lane0;
  assign early0_BranchPlugin_logic_pcPort_payload_laneAge = toplevel_execute_ctrl3_down_LANE_AGE_lane0;
  assign early0_BranchPlugin_logic_historyPort_valid = early0_BranchPlugin_logic_jumpLogic_doIt;
  assign early0_BranchPlugin_logic_historyPort_payload_history = early0_BranchPlugin_logic_jumpLogic_history_next;
  assign early0_BranchPlugin_logic_historyPort_payload_age = toplevel_execute_ctrl3_down_LANE_AGE_lane0;
  assign early0_BranchPlugin_logic_flushPort_valid = early0_BranchPlugin_logic_jumpLogic_doIt;
  assign early0_BranchPlugin_logic_flushPort_payload_uopId = toplevel_execute_ctrl3_down_Decode_UOP_ID_lane0;
  assign early0_BranchPlugin_logic_flushPort_payload_laneAge = toplevel_execute_ctrl3_down_LANE_AGE_lane0;
  assign early0_BranchPlugin_logic_flushPort_payload_self = 1'b0;
  assign toplevel_execute_ctrl3_down_early0_BranchPlugin_logic_jumpLogic_MISSALIGNED_lane0 = ((toplevel_execute_ctrl3_down_early0_BranchPlugin_pcCalc_PC_TRUE_lane0[0 : 0] != 1'b0) && toplevel_execute_ctrl3_down_early0_BranchPlugin_logic_jumpLogic_COND_lane0);
  assign toplevel_execute_ctrl3_down_early0_BranchPlugin_logic_jumpLogic_IS_JAL_lane0 = (toplevel_execute_ctrl3_down_BranchPlugin_BRANCH_CTRL_lane0 == BranchPlugin_BranchCtrlEnum_JAL);
  assign toplevel_execute_ctrl3_down_early0_BranchPlugin_logic_jumpLogic_IS_JALR_lane0 = (toplevel_execute_ctrl3_down_BranchPlugin_BRANCH_CTRL_lane0 == BranchPlugin_BranchCtrlEnum_JALR);
  assign early0_BranchPlugin_logic_jumpLogic_rdLink = (|{(toplevel_execute_ctrl3_down_Decode_UOP_lane0[11 : 7] == 5'h05),(toplevel_execute_ctrl3_down_Decode_UOP_lane0[11 : 7] == 5'h01)});
  assign early0_BranchPlugin_logic_jumpLogic_rs1Link = (|{(toplevel_execute_ctrl3_down_Decode_UOP_lane0[19 : 15] == 5'h05),(toplevel_execute_ctrl3_down_Decode_UOP_lane0[19 : 15] == 5'h01)});
  assign early0_BranchPlugin_logic_jumpLogic_rdEquRs1 = (toplevel_execute_ctrl3_down_Decode_UOP_lane0[11 : 7] == toplevel_execute_ctrl3_down_Decode_UOP_lane0[19 : 15]);
  assign early0_BranchPlugin_logic_wb_valid = toplevel_execute_ctrl2_down_early0_BranchPlugin_SEL_lane0;
  assign early0_BranchPlugin_logic_wb_payload = toplevel_execute_ctrl2_down_early0_BranchPlugin_pcCalc_PC_FALSE_lane0;
  always @(*) begin
    early0_EnvPlugin_logic_flushPort_valid = 1'b0;
    if(when_EnvPlugin_l116) begin
      early0_EnvPlugin_logic_flushPort_valid = 1'b1;
    end
  end

  assign early0_EnvPlugin_logic_flushPort_payload_uopId = toplevel_execute_ctrl2_down_Decode_UOP_ID_lane0;
  assign early0_EnvPlugin_logic_flushPort_payload_laneAge = toplevel_execute_ctrl2_down_LANE_AGE_lane0;
  assign early0_EnvPlugin_logic_flushPort_payload_self = 1'b0;
  always @(*) begin
    early0_EnvPlugin_logic_trapPort_valid = 1'b0;
    if(when_EnvPlugin_l116) begin
      early0_EnvPlugin_logic_trapPort_valid = 1'b1;
    end
  end

  always @(*) begin
    early0_EnvPlugin_logic_trapPort_payload_exception = 1'b1;
    case(toplevel_execute_ctrl2_down_early0_EnvPlugin_OP_lane0)
      EnvPluginOp_EBREAK : begin
      end
      EnvPluginOp_ECALL : begin
      end
      EnvPluginOp_PRIV_RET : begin
        if(when_EnvPlugin_l83) begin
          early0_EnvPlugin_logic_trapPort_payload_exception = 1'b0;
        end
      end
      EnvPluginOp_WFI : begin
        if(when_EnvPlugin_l92) begin
          early0_EnvPlugin_logic_trapPort_payload_exception = 1'b0;
        end
      end
      EnvPluginOp_FENCE_I : begin
        early0_EnvPlugin_logic_trapPort_payload_exception = 1'b0;
      end
      default : begin
        if(when_EnvPlugin_l107) begin
          early0_EnvPlugin_logic_trapPort_payload_exception = 1'b0;
        end
      end
    endcase
  end

  assign early0_EnvPlugin_logic_trapPort_payload_tval = ((toplevel_execute_ctrl2_down_early0_EnvPlugin_OP_lane0 == EnvPluginOp_EBREAK) ? toplevel_execute_ctrl2_down_PC_lane0 : 32'h0);
  always @(*) begin
    early0_EnvPlugin_logic_trapPort_payload_code = 4'b0010;
    case(toplevel_execute_ctrl2_down_early0_EnvPlugin_OP_lane0)
      EnvPluginOp_EBREAK : begin
        early0_EnvPlugin_logic_trapPort_payload_code = 4'b0011;
      end
      EnvPluginOp_ECALL : begin
        early0_EnvPlugin_logic_trapPort_payload_code = (_zz_early0_EnvPlugin_logic_trapPort_payload_code | 4'b1000);
      end
      EnvPluginOp_PRIV_RET : begin
        if(when_EnvPlugin_l83) begin
          early0_EnvPlugin_logic_trapPort_payload_code = 4'b0001;
        end
      end
      EnvPluginOp_WFI : begin
        if(when_EnvPlugin_l92) begin
          early0_EnvPlugin_logic_trapPort_payload_code = 4'b1000;
        end
      end
      EnvPluginOp_FENCE_I : begin
        early0_EnvPlugin_logic_trapPort_payload_code = 4'b0010;
      end
      default : begin
        if(when_EnvPlugin_l107) begin
          early0_EnvPlugin_logic_trapPort_payload_code = 4'b0110;
        end
      end
    endcase
  end

  always @(*) begin
    early0_EnvPlugin_logic_trapPort_payload_arg = 3'bxxx;
    case(toplevel_execute_ctrl2_down_early0_EnvPlugin_OP_lane0)
      EnvPluginOp_EBREAK : begin
      end
      EnvPluginOp_ECALL : begin
      end
      EnvPluginOp_PRIV_RET : begin
        if(when_EnvPlugin_l83) begin
          early0_EnvPlugin_logic_trapPort_payload_arg[1 : 0] = early0_EnvPlugin_logic_exe_xretPriv;
        end
      end
      EnvPluginOp_WFI : begin
      end
      EnvPluginOp_FENCE_I : begin
      end
      default : begin
      end
    endcase
  end

  assign early0_EnvPlugin_logic_trapPort_payload_laneAge = toplevel_execute_ctrl2_down_LANE_AGE_lane0;
  assign early0_EnvPlugin_logic_exe_privilege = PrivilegedPlugin_logic_harts_0_privilege;
  assign early0_EnvPlugin_logic_exe_xretPriv = toplevel_execute_ctrl2_down_Decode_UOP_lane0[29 : 28];
  always @(*) begin
    early0_EnvPlugin_logic_exe_commit = 1'b0;
    case(toplevel_execute_ctrl2_down_early0_EnvPlugin_OP_lane0)
      EnvPluginOp_EBREAK : begin
      end
      EnvPluginOp_ECALL : begin
      end
      EnvPluginOp_PRIV_RET : begin
        if(when_EnvPlugin_l83) begin
          early0_EnvPlugin_logic_exe_commit = 1'b1;
        end
      end
      EnvPluginOp_WFI : begin
        if(when_EnvPlugin_l92) begin
          early0_EnvPlugin_logic_exe_commit = 1'b1;
        end
      end
      EnvPluginOp_FENCE_I : begin
        early0_EnvPlugin_logic_exe_commit = 1'b1;
      end
      default : begin
        if(when_EnvPlugin_l107) begin
          early0_EnvPlugin_logic_exe_commit = 1'b1;
        end
      end
    endcase
  end

  assign early0_EnvPlugin_logic_exe_retKo = ((PrivilegedPlugin_logic_harts_0_m_status_tsr && (early0_EnvPlugin_logic_exe_privilege == 2'b01)) && (early0_EnvPlugin_logic_exe_xretPriv == 2'b01));
  assign early0_EnvPlugin_logic_exe_vmaKo = (((early0_EnvPlugin_logic_exe_privilege == 2'b01) && PrivilegedPlugin_logic_harts_0_m_status_tvm) || (early0_EnvPlugin_logic_exe_privilege == 2'b00));
  assign when_EnvPlugin_l83 = ((early0_EnvPlugin_logic_exe_xretPriv <= PrivilegedPlugin_logic_harts_0_privilege) && (! early0_EnvPlugin_logic_exe_retKo));
  assign when_EnvPlugin_l92 = ((early0_EnvPlugin_logic_exe_privilege == 2'b11) || ((! PrivilegedPlugin_logic_harts_0_m_status_tw) && (1'b0 || (early0_EnvPlugin_logic_exe_privilege == 2'b01))));
  assign when_EnvPlugin_l107 = (! early0_EnvPlugin_logic_exe_vmaKo);
  assign when_EnvPlugin_l116 = (toplevel_execute_ctrl2_up_LANE_SEL_lane0 && toplevel_execute_ctrl2_down_early0_EnvPlugin_SEL_lane0);
  assign when_EnvPlugin_l120 = (! early0_EnvPlugin_logic_exe_commit);
  assign toplevel_execute_ctrl2_down_early1_BranchPlugin_logic_alu_EQ_lane1 = ($signed(toplevel_execute_ctrl2_down_early1_SrcPlugin_SRC1_lane1) == $signed(toplevel_execute_ctrl2_down_early1_SrcPlugin_SRC2_lane1));
  assign toplevel_execute_ctrl2_down_early1_BranchPlugin_logic_alu_btb_BAD_TARGET_lane1 = (toplevel_execute_ctrl2_down_Prediction_ALIGNED_JUMPED_PC_lane1 != toplevel_execute_ctrl2_down_early1_BranchPlugin_pcCalc_PC_TRUE_lane1);
  assign early1_BranchPlugin_logic_alu_expectedMsb = (MmuPlugin_api_fetchTranslationEnable ? _zz_early1_BranchPlugin_logic_alu_expectedMsb[31] : 1'b0);
  assign toplevel_execute_ctrl2_down_early1_BranchPlugin_logic_alu_MSB_FAILED_lane1 = ((toplevel_execute_ctrl2_down_BranchPlugin_BRANCH_CTRL_lane1 == BranchPlugin_BranchCtrlEnum_JALR) && 1'b0);
  assign switch_Misc_l241_1 = toplevel_execute_ctrl3_down_Decode_UOP_lane1[14 : 12];
  always @(*) begin
    casez(switch_Misc_l241_1)
      3'b000 : begin
        _zz_toplevel_execute_ctrl3_down_early1_BranchPlugin_logic_jumpLogic_COND_lane1 = toplevel_execute_ctrl3_down_early1_BranchPlugin_logic_alu_EQ_lane1;
      end
      3'b001 : begin
        _zz_toplevel_execute_ctrl3_down_early1_BranchPlugin_logic_jumpLogic_COND_lane1 = (! toplevel_execute_ctrl3_down_early1_BranchPlugin_logic_alu_EQ_lane1);
      end
      3'b1?1 : begin
        _zz_toplevel_execute_ctrl3_down_early1_BranchPlugin_logic_jumpLogic_COND_lane1 = (! toplevel_execute_ctrl3_down_early1_SrcPlugin_LESS_lane1);
      end
      default : begin
        _zz_toplevel_execute_ctrl3_down_early1_BranchPlugin_logic_jumpLogic_COND_lane1 = toplevel_execute_ctrl3_down_early1_SrcPlugin_LESS_lane1;
      end
    endcase
  end

  always @(*) begin
    case(toplevel_execute_ctrl3_down_BranchPlugin_BRANCH_CTRL_lane1)
      BranchPlugin_BranchCtrlEnum_JALR : begin
        _zz_toplevel_execute_ctrl3_down_early1_BranchPlugin_logic_jumpLogic_COND_lane1_1 = 1'b1;
      end
      BranchPlugin_BranchCtrlEnum_JAL : begin
        _zz_toplevel_execute_ctrl3_down_early1_BranchPlugin_logic_jumpLogic_COND_lane1_1 = 1'b1;
      end
      default : begin
        _zz_toplevel_execute_ctrl3_down_early1_BranchPlugin_logic_jumpLogic_COND_lane1_1 = _zz_toplevel_execute_ctrl3_down_early1_BranchPlugin_logic_jumpLogic_COND_lane1;
      end
    endcase
  end

  assign toplevel_execute_ctrl3_down_early1_BranchPlugin_logic_jumpLogic_COND_lane1 = _zz_toplevel_execute_ctrl3_down_early1_BranchPlugin_logic_jumpLogic_COND_lane1_1;
  assign toplevel_execute_ctrl3_down_early1_BranchPlugin_logic_jumpLogic_btb_REAL_TARGET_lane1 = (toplevel_execute_ctrl3_down_early1_BranchPlugin_logic_jumpLogic_COND_lane1 ? toplevel_execute_ctrl3_down_early1_BranchPlugin_pcCalc_PC_TRUE_lane1 : toplevel_execute_ctrl3_down_early1_BranchPlugin_pcCalc_PC_FALSE_lane1);
  assign early1_BranchPlugin_logic_jumpLogic_wrongCond = (toplevel_execute_ctrl3_down_Prediction_ALIGNED_JUMPED_lane1 != toplevel_execute_ctrl3_down_early1_BranchPlugin_logic_jumpLogic_COND_lane1);
  assign early1_BranchPlugin_logic_jumpLogic_needFix = ((early1_BranchPlugin_logic_jumpLogic_wrongCond || (toplevel_execute_ctrl3_down_early1_BranchPlugin_logic_jumpLogic_COND_lane1 && toplevel_execute_ctrl3_down_early1_BranchPlugin_logic_alu_btb_BAD_TARGET_lane1)) || toplevel_execute_ctrl3_down_early1_BranchPlugin_logic_alu_MSB_FAILED_lane1);
  assign early1_BranchPlugin_logic_jumpLogic_doIt = ((toplevel_execute_ctrl3_up_LANE_SEL_lane1 && toplevel_execute_ctrl3_down_early1_BranchPlugin_SEL_lane1) && early1_BranchPlugin_logic_jumpLogic_needFix);
  assign early1_BranchPlugin_logic_jumpLogic_history_fromFetch_slice = toplevel_execute_ctrl3_down_PC_lane1[2 : 1];
  assign early1_BranchPlugin_logic_jumpLogic_history_fromFetch_shifter = toplevel_execute_ctrl3_down_Prediction_BRANCH_HISTORY_lane1;
  assign when_BranchPlugin_l206_3 = ((early1_BranchPlugin_logic_jumpLogic_history_fromFetch_slice < 2'b00) && toplevel_execute_ctrl3_down_Prediction_ALIGNED_SLICES_BRANCH_lane1[0]);
  assign when_BranchPlugin_l206_4 = ((early1_BranchPlugin_logic_jumpLogic_history_fromFetch_slice < 2'b01) && toplevel_execute_ctrl3_down_Prediction_ALIGNED_SLICES_BRANCH_lane1[1]);
  assign when_BranchPlugin_l206_5 = ((early1_BranchPlugin_logic_jumpLogic_history_fromFetch_slice < 2'b10) && toplevel_execute_ctrl3_down_Prediction_ALIGNED_SLICES_BRANCH_lane1[2]);
  assign when_BranchPlugin_l210_1 = (toplevel_execute_ctrl3_down_BranchPlugin_BRANCH_CTRL_lane1 == BranchPlugin_BranchCtrlEnum_B);
  assign early1_BranchPlugin_logic_jumpLogic_history_next = early1_BranchPlugin_logic_jumpLogic_history_fromFetch_shifter_4;
  assign early1_BranchPlugin_logic_jumpLogic_history_fetched = toplevel_execute_ctrl3_down_Prediction_BRANCH_HISTORY_lane1;
  assign early1_BranchPlugin_logic_pcPort_valid = early1_BranchPlugin_logic_jumpLogic_doIt;
  assign early1_BranchPlugin_logic_pcPort_payload_fault = toplevel_execute_ctrl3_down_early1_BranchPlugin_logic_alu_MSB_FAILED_lane1;
  assign early1_BranchPlugin_logic_pcPort_payload_pc = toplevel_execute_ctrl3_down_early1_BranchPlugin_logic_jumpLogic_btb_REAL_TARGET_lane1;
  assign early1_BranchPlugin_logic_pcPort_payload_laneAge = toplevel_execute_ctrl3_down_LANE_AGE_lane1;
  assign early1_BranchPlugin_logic_historyPort_valid = early1_BranchPlugin_logic_jumpLogic_doIt;
  assign early1_BranchPlugin_logic_historyPort_payload_history = early1_BranchPlugin_logic_jumpLogic_history_next;
  assign early1_BranchPlugin_logic_historyPort_payload_age = toplevel_execute_ctrl3_down_LANE_AGE_lane1;
  assign early1_BranchPlugin_logic_flushPort_valid = early1_BranchPlugin_logic_jumpLogic_doIt;
  assign early1_BranchPlugin_logic_flushPort_payload_uopId = toplevel_execute_ctrl3_down_Decode_UOP_ID_lane1;
  assign early1_BranchPlugin_logic_flushPort_payload_laneAge = toplevel_execute_ctrl3_down_LANE_AGE_lane1;
  assign early1_BranchPlugin_logic_flushPort_payload_self = 1'b0;
  assign toplevel_execute_ctrl3_down_early1_BranchPlugin_logic_jumpLogic_MISSALIGNED_lane1 = ((toplevel_execute_ctrl3_down_early1_BranchPlugin_pcCalc_PC_TRUE_lane1[0 : 0] != 1'b0) && toplevel_execute_ctrl3_down_early1_BranchPlugin_logic_jumpLogic_COND_lane1);
  assign toplevel_execute_ctrl3_down_early1_BranchPlugin_logic_jumpLogic_IS_JAL_lane1 = (toplevel_execute_ctrl3_down_BranchPlugin_BRANCH_CTRL_lane1 == BranchPlugin_BranchCtrlEnum_JAL);
  assign toplevel_execute_ctrl3_down_early1_BranchPlugin_logic_jumpLogic_IS_JALR_lane1 = (toplevel_execute_ctrl3_down_BranchPlugin_BRANCH_CTRL_lane1 == BranchPlugin_BranchCtrlEnum_JALR);
  assign early1_BranchPlugin_logic_jumpLogic_rdLink = (|{(toplevel_execute_ctrl3_down_Decode_UOP_lane1[11 : 7] == 5'h05),(toplevel_execute_ctrl3_down_Decode_UOP_lane1[11 : 7] == 5'h01)});
  assign early1_BranchPlugin_logic_jumpLogic_rs1Link = (|{(toplevel_execute_ctrl3_down_Decode_UOP_lane1[19 : 15] == 5'h05),(toplevel_execute_ctrl3_down_Decode_UOP_lane1[19 : 15] == 5'h01)});
  assign early1_BranchPlugin_logic_jumpLogic_rdEquRs1 = (toplevel_execute_ctrl3_down_Decode_UOP_lane1[11 : 7] == toplevel_execute_ctrl3_down_Decode_UOP_lane1[19 : 15]);
  assign early1_BranchPlugin_logic_wb_valid = toplevel_execute_ctrl2_down_early1_BranchPlugin_SEL_lane1;
  assign early1_BranchPlugin_logic_wb_payload = toplevel_execute_ctrl2_down_early1_BranchPlugin_pcCalc_PC_FALSE_lane1;
  assign FetchL1TileLinkPlugin_logic_down_a_valid = FetchL1Plugin_logic_bus_cmd_valid;
  assign FetchL1TileLinkPlugin_logic_down_a_payload_opcode = A_GET;
  assign FetchL1TileLinkPlugin_logic_down_a_payload_param = 3'b000;
  assign FetchL1TileLinkPlugin_logic_down_a_payload_address = FetchL1Plugin_logic_bus_cmd_payload_address;
  assign FetchL1TileLinkPlugin_logic_down_a_payload_size = 3'b110;
  assign FetchL1Plugin_logic_bus_cmd_ready = FetchL1TileLinkPlugin_logic_down_a_ready;
  assign FetchL1Plugin_logic_bus_rsp_valid = FetchL1TileLinkPlugin_logic_down_d_valid;
  assign FetchL1Plugin_logic_bus_rsp_payload_data = FetchL1TileLinkPlugin_logic_down_d_payload_data;
  assign FetchL1Plugin_logic_bus_rsp_payload_error = (FetchL1TileLinkPlugin_logic_down_d_payload_denied || FetchL1TileLinkPlugin_logic_down_d_payload_corrupt);
  assign FetchL1TileLinkPlugin_logic_down_d_ready = 1'b1;
  assign MmuPlugin_logic_satpModeWrite = CsrAccessPlugin_bus_write_bits[31 : 31];
  always @(*) begin
    _zz_toplevel_execute_ctrl1_down_early0_SrcPlugin_SRC1_lane0 = 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
    case(toplevel_execute_ctrl1_down_early0_SrcPlugin_logic_SRC1_CTRL_lane0)
      1'b0 : begin
        _zz_toplevel_execute_ctrl1_down_early0_SrcPlugin_SRC1_lane0 = toplevel_execute_ctrl1_down_integer_RS1_lane0;
      end
      default : begin
        _zz_toplevel_execute_ctrl1_down_early0_SrcPlugin_SRC1_lane0 = {toplevel_execute_ctrl1_down_Decode_UOP_lane0[31 : 12],12'h0};
      end
    endcase
  end

  assign toplevel_execute_ctrl1_down_early0_SrcPlugin_SRC1_lane0 = _zz_toplevel_execute_ctrl1_down_early0_SrcPlugin_SRC1_lane0;
  always @(*) begin
    _zz_toplevel_execute_ctrl1_down_early0_SrcPlugin_SRC2_lane0 = 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
    case(toplevel_execute_ctrl1_down_early0_SrcPlugin_logic_SRC2_CTRL_lane0)
      2'b00 : begin
        _zz_toplevel_execute_ctrl1_down_early0_SrcPlugin_SRC2_lane0 = toplevel_execute_ctrl1_down_integer_RS2_lane0;
      end
      2'b01 : begin
        _zz_toplevel_execute_ctrl1_down_early0_SrcPlugin_SRC2_lane0 = {{20{_zz__zz_toplevel_execute_ctrl1_down_early0_SrcPlugin_SRC2_lane0[11]}}, _zz__zz_toplevel_execute_ctrl1_down_early0_SrcPlugin_SRC2_lane0};
      end
      2'b10 : begin
        _zz_toplevel_execute_ctrl1_down_early0_SrcPlugin_SRC2_lane0 = toplevel_execute_ctrl1_down_PC_lane0;
      end
      default : begin
        _zz_toplevel_execute_ctrl1_down_early0_SrcPlugin_SRC2_lane0 = {{20{_zz__zz_toplevel_execute_ctrl1_down_early0_SrcPlugin_SRC2_lane0_1[11]}}, _zz__zz_toplevel_execute_ctrl1_down_early0_SrcPlugin_SRC2_lane0_1};
      end
    endcase
  end

  assign toplevel_execute_ctrl1_down_early0_SrcPlugin_SRC2_lane0 = _zz_toplevel_execute_ctrl1_down_early0_SrcPlugin_SRC2_lane0;
  always @(*) begin
    early0_SrcPlugin_logic_addsub_combined_rs2Patched = toplevel_execute_ctrl2_down_early0_SrcPlugin_SRC2_lane0;
    if(toplevel_execute_ctrl2_down_SrcStageables_REVERT_lane0) begin
      early0_SrcPlugin_logic_addsub_combined_rs2Patched = (~ toplevel_execute_ctrl2_down_early0_SrcPlugin_SRC2_lane0);
    end
    if(toplevel_execute_ctrl2_down_SrcStageables_ZERO_lane0) begin
      early0_SrcPlugin_logic_addsub_combined_rs2Patched = 32'h0;
    end
  end

  assign toplevel_execute_ctrl2_down_early0_SrcPlugin_ADD_SUB_lane0 = ($signed(_zz_toplevel_execute_ctrl2_down_early0_SrcPlugin_ADD_SUB_lane0) + $signed(_zz_toplevel_execute_ctrl2_down_early0_SrcPlugin_ADD_SUB_lane0_1));
  assign toplevel_execute_ctrl2_down_early0_SrcPlugin_LESS_lane0 = ((toplevel_execute_ctrl2_down_early0_SrcPlugin_SRC1_lane0[31] == toplevel_execute_ctrl2_down_early0_SrcPlugin_SRC2_lane0[31]) ? toplevel_execute_ctrl2_down_early0_SrcPlugin_ADD_SUB_lane0[31] : (toplevel_execute_ctrl2_down_SrcStageables_UNSIGNED_lane0 ? toplevel_execute_ctrl2_down_early0_SrcPlugin_SRC2_lane0[31] : toplevel_execute_ctrl2_down_early0_SrcPlugin_SRC1_lane0[31]));
  assign lane0_IntFormatPlugin_logic_stages_0_hits = early0_IntAluPlugin_logic_wb_valid;
  assign lane0_IntFormatPlugin_logic_stages_0_wb_valid = (toplevel_execute_ctrl2_up_LANE_SEL_lane0 && (|lane0_IntFormatPlugin_logic_stages_0_hits));
  assign lane0_IntFormatPlugin_logic_stages_0_raw = early0_IntAluPlugin_logic_wb_payload;
  assign lane0_IntFormatPlugin_logic_stages_0_wb_payload = lane0_IntFormatPlugin_logic_stages_0_raw;
  assign lane0_IntFormatPlugin_logic_stages_1_hits = {CsrAccessPlugin_logic_wbWi_valid,{early0_DivPlugin_logic_formatBus_valid,early0_BarrelShifterPlugin_logic_wb_valid}};
  assign lane0_IntFormatPlugin_logic_stages_1_wb_valid = (toplevel_execute_ctrl3_up_LANE_SEL_lane0 && (|lane0_IntFormatPlugin_logic_stages_1_hits));
  assign lane0_IntFormatPlugin_logic_stages_1_raw = (((lane0_IntFormatPlugin_logic_stages_1_hits[0] ? early0_BarrelShifterPlugin_logic_wb_payload : 32'h0) | (lane0_IntFormatPlugin_logic_stages_1_hits[1] ? early0_DivPlugin_logic_formatBus_payload : 32'h0)) | (lane0_IntFormatPlugin_logic_stages_1_hits[2] ? CsrAccessPlugin_logic_wbWi_payload : 32'h0));
  assign lane0_IntFormatPlugin_logic_stages_1_wb_payload = lane0_IntFormatPlugin_logic_stages_1_raw;
  assign lane0_IntFormatPlugin_logic_stages_2_hits = {LsuPlugin_logic_iwb_valid,{late0_BarrelShifterPlugin_logic_wb_valid,{late0_IntAluPlugin_logic_wb_valid,early0_MulPlugin_logic_formatBus_valid}}};
  assign lane0_IntFormatPlugin_logic_stages_2_wb_valid = (toplevel_execute_ctrl4_up_LANE_SEL_lane0 && (|lane0_IntFormatPlugin_logic_stages_2_hits));
  assign lane0_IntFormatPlugin_logic_stages_2_raw = (((lane0_IntFormatPlugin_logic_stages_2_hits[0] ? early0_MulPlugin_logic_formatBus_payload : 32'h0) | (lane0_IntFormatPlugin_logic_stages_2_hits[1] ? late0_IntAluPlugin_logic_wb_payload : 32'h0)) | ((lane0_IntFormatPlugin_logic_stages_2_hits[2] ? late0_BarrelShifterPlugin_logic_wb_payload : 32'h0) | (lane0_IntFormatPlugin_logic_stages_2_hits[3] ? LsuPlugin_logic_iwb_payload : 32'h0)));
  always @(*) begin
    lane0_IntFormatPlugin_logic_stages_2_wb_payload = lane0_IntFormatPlugin_logic_stages_2_raw;
    if(lane0_IntFormatPlugin_logic_stages_2_segments_0_doIt) begin
      lane0_IntFormatPlugin_logic_stages_2_wb_payload[15 : 8] = {8{lane0_IntFormatPlugin_logic_stages_2_segments_0_sign_value}};
    end
    if(lane0_IntFormatPlugin_logic_stages_2_segments_1_doIt) begin
      lane0_IntFormatPlugin_logic_stages_2_wb_payload[31 : 16] = {16{lane0_IntFormatPlugin_logic_stages_2_segments_1_sign_value}};
    end
  end

  assign lane0_IntFormatPlugin_logic_stages_2_segments_0_sign_sels_0 = lane0_IntFormatPlugin_logic_stages_2_raw[7];
  always @(*) begin
    _zz_lane0_IntFormatPlugin_logic_stages_2_segments_0_sign_value = 1'bx;
    case(toplevel_execute_ctrl4_down_lane0_IntFormatPlugin_logic_WIDTH_ID_lane0)
      2'b00 : begin
        _zz_lane0_IntFormatPlugin_logic_stages_2_segments_0_sign_value = lane0_IntFormatPlugin_logic_stages_2_segments_0_sign_sels_0;
      end
      default : begin
      end
    endcase
  end

  assign lane0_IntFormatPlugin_logic_stages_2_segments_0_sign_value = (toplevel_execute_ctrl4_down_lane0_IntFormatPlugin_logic_SIGNED_lane0 && _zz_lane0_IntFormatPlugin_logic_stages_2_segments_0_sign_value);
  assign lane0_IntFormatPlugin_logic_stages_2_segments_0_doIt = (toplevel_execute_ctrl4_down_lane0_IntFormatPlugin_logic_WIDTH_ID_lane0 < 2'b01);
  assign lane0_IntFormatPlugin_logic_stages_2_segments_1_sign_sels_0 = lane0_IntFormatPlugin_logic_stages_2_raw[7];
  assign lane0_IntFormatPlugin_logic_stages_2_segments_1_sign_sels_1 = lane0_IntFormatPlugin_logic_stages_2_raw[15];
  always @(*) begin
    _zz_lane0_IntFormatPlugin_logic_stages_2_segments_1_sign_value = 1'bx;
    case(toplevel_execute_ctrl4_down_lane0_IntFormatPlugin_logic_WIDTH_ID_lane0)
      2'b00 : begin
        _zz_lane0_IntFormatPlugin_logic_stages_2_segments_1_sign_value = lane0_IntFormatPlugin_logic_stages_2_segments_1_sign_sels_0;
      end
      2'b01 : begin
        _zz_lane0_IntFormatPlugin_logic_stages_2_segments_1_sign_value = lane0_IntFormatPlugin_logic_stages_2_segments_1_sign_sels_1;
      end
      default : begin
      end
    endcase
  end

  assign lane0_IntFormatPlugin_logic_stages_2_segments_1_sign_value = (toplevel_execute_ctrl4_down_lane0_IntFormatPlugin_logic_SIGNED_lane0 && _zz_lane0_IntFormatPlugin_logic_stages_2_segments_1_sign_value);
  assign lane0_IntFormatPlugin_logic_stages_2_segments_1_doIt = (toplevel_execute_ctrl4_down_lane0_IntFormatPlugin_logic_WIDTH_ID_lane0 < 2'b10);
  always @(*) begin
    _zz_toplevel_execute_ctrl3_down_late0_SrcPlugin_SRC1_lane0 = 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
    case(toplevel_execute_ctrl3_down_late0_SrcPlugin_logic_SRC1_CTRL_lane0)
      1'b0 : begin
        _zz_toplevel_execute_ctrl3_down_late0_SrcPlugin_SRC1_lane0 = toplevel_execute_ctrl3_down_integer_RS1_lane0;
      end
      default : begin
        _zz_toplevel_execute_ctrl3_down_late0_SrcPlugin_SRC1_lane0 = {toplevel_execute_ctrl3_down_Decode_UOP_lane0[31 : 12],12'h0};
      end
    endcase
  end

  assign toplevel_execute_ctrl3_down_late0_SrcPlugin_SRC1_lane0 = _zz_toplevel_execute_ctrl3_down_late0_SrcPlugin_SRC1_lane0;
  always @(*) begin
    _zz_toplevel_execute_ctrl3_down_late0_SrcPlugin_SRC2_lane0 = 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
    case(toplevel_execute_ctrl3_down_late0_SrcPlugin_logic_SRC2_CTRL_lane0)
      2'b00 : begin
        _zz_toplevel_execute_ctrl3_down_late0_SrcPlugin_SRC2_lane0 = toplevel_execute_ctrl3_down_integer_RS2_lane0;
      end
      2'b01 : begin
        _zz_toplevel_execute_ctrl3_down_late0_SrcPlugin_SRC2_lane0 = {{20{_zz__zz_toplevel_execute_ctrl3_down_late0_SrcPlugin_SRC2_lane0[11]}}, _zz__zz_toplevel_execute_ctrl3_down_late0_SrcPlugin_SRC2_lane0};
      end
      2'b10 : begin
        _zz_toplevel_execute_ctrl3_down_late0_SrcPlugin_SRC2_lane0 = toplevel_execute_ctrl3_down_PC_lane0;
      end
      default : begin
      end
    endcase
  end

  assign toplevel_execute_ctrl3_down_late0_SrcPlugin_SRC2_lane0 = _zz_toplevel_execute_ctrl3_down_late0_SrcPlugin_SRC2_lane0;
  always @(*) begin
    late0_SrcPlugin_logic_addsub_combined_rs2Patched = toplevel_execute_ctrl4_down_late0_SrcPlugin_SRC2_lane0;
    if(toplevel_execute_ctrl4_down_SrcStageables_REVERT_lane0) begin
      late0_SrcPlugin_logic_addsub_combined_rs2Patched = (~ toplevel_execute_ctrl4_down_late0_SrcPlugin_SRC2_lane0);
    end
    if(toplevel_execute_ctrl4_down_SrcStageables_ZERO_lane0) begin
      late0_SrcPlugin_logic_addsub_combined_rs2Patched = 32'h0;
    end
  end

  assign toplevel_execute_ctrl4_down_late0_SrcPlugin_ADD_SUB_lane0 = ($signed(_zz_toplevel_execute_ctrl4_down_late0_SrcPlugin_ADD_SUB_lane0) + $signed(_zz_toplevel_execute_ctrl4_down_late0_SrcPlugin_ADD_SUB_lane0_1));
  assign toplevel_execute_ctrl4_down_late0_SrcPlugin_LESS_lane0 = ((toplevel_execute_ctrl4_down_late0_SrcPlugin_SRC1_lane0[31] == toplevel_execute_ctrl4_down_late0_SrcPlugin_SRC2_lane0[31]) ? toplevel_execute_ctrl4_down_late0_SrcPlugin_ADD_SUB_lane0[31] : (toplevel_execute_ctrl4_down_SrcStageables_UNSIGNED_lane0 ? toplevel_execute_ctrl4_down_late0_SrcPlugin_SRC2_lane0[31] : toplevel_execute_ctrl4_down_late0_SrcPlugin_SRC1_lane0[31]));
  always @(*) begin
    _zz_toplevel_execute_ctrl1_down_early1_SrcPlugin_SRC1_lane1 = 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
    case(toplevel_execute_ctrl1_down_early1_SrcPlugin_logic_SRC1_CTRL_lane1)
      1'b0 : begin
        _zz_toplevel_execute_ctrl1_down_early1_SrcPlugin_SRC1_lane1 = toplevel_execute_ctrl1_down_integer_RS1_lane1;
      end
      default : begin
        _zz_toplevel_execute_ctrl1_down_early1_SrcPlugin_SRC1_lane1 = {toplevel_execute_ctrl1_down_Decode_UOP_lane1[31 : 12],12'h0};
      end
    endcase
  end

  assign toplevel_execute_ctrl1_down_early1_SrcPlugin_SRC1_lane1 = _zz_toplevel_execute_ctrl1_down_early1_SrcPlugin_SRC1_lane1;
  always @(*) begin
    _zz_toplevel_execute_ctrl1_down_early1_SrcPlugin_SRC2_lane1 = 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
    case(toplevel_execute_ctrl1_down_early1_SrcPlugin_logic_SRC2_CTRL_lane1)
      2'b00 : begin
        _zz_toplevel_execute_ctrl1_down_early1_SrcPlugin_SRC2_lane1 = toplevel_execute_ctrl1_down_integer_RS2_lane1;
      end
      2'b01 : begin
        _zz_toplevel_execute_ctrl1_down_early1_SrcPlugin_SRC2_lane1 = {{20{_zz__zz_toplevel_execute_ctrl1_down_early1_SrcPlugin_SRC2_lane1[11]}}, _zz__zz_toplevel_execute_ctrl1_down_early1_SrcPlugin_SRC2_lane1};
      end
      2'b10 : begin
        _zz_toplevel_execute_ctrl1_down_early1_SrcPlugin_SRC2_lane1 = toplevel_execute_ctrl1_down_PC_lane1;
      end
      default : begin
      end
    endcase
  end

  assign toplevel_execute_ctrl1_down_early1_SrcPlugin_SRC2_lane1 = _zz_toplevel_execute_ctrl1_down_early1_SrcPlugin_SRC2_lane1;
  always @(*) begin
    early1_SrcPlugin_logic_addsub_combined_rs2Patched = toplevel_execute_ctrl2_down_early1_SrcPlugin_SRC2_lane1;
    if(toplevel_execute_ctrl2_down_SrcStageables_REVERT_lane1) begin
      early1_SrcPlugin_logic_addsub_combined_rs2Patched = (~ toplevel_execute_ctrl2_down_early1_SrcPlugin_SRC2_lane1);
    end
    if(toplevel_execute_ctrl2_down_SrcStageables_ZERO_lane1) begin
      early1_SrcPlugin_logic_addsub_combined_rs2Patched = 32'h0;
    end
  end

  assign toplevel_execute_ctrl2_down_early1_SrcPlugin_ADD_SUB_lane1 = ($signed(_zz_toplevel_execute_ctrl2_down_early1_SrcPlugin_ADD_SUB_lane1) + $signed(_zz_toplevel_execute_ctrl2_down_early1_SrcPlugin_ADD_SUB_lane1_1));
  assign toplevel_execute_ctrl2_down_early1_SrcPlugin_LESS_lane1 = ((toplevel_execute_ctrl2_down_early1_SrcPlugin_SRC1_lane1[31] == toplevel_execute_ctrl2_down_early1_SrcPlugin_SRC2_lane1[31]) ? toplevel_execute_ctrl2_down_early1_SrcPlugin_ADD_SUB_lane1[31] : (toplevel_execute_ctrl2_down_SrcStageables_UNSIGNED_lane1 ? toplevel_execute_ctrl2_down_early1_SrcPlugin_SRC2_lane1[31] : toplevel_execute_ctrl2_down_early1_SrcPlugin_SRC1_lane1[31]));
  assign lane1_IntFormatPlugin_logic_stages_0_hits = early1_IntAluPlugin_logic_wb_valid;
  assign lane1_IntFormatPlugin_logic_stages_0_wb_valid = (toplevel_execute_ctrl2_up_LANE_SEL_lane1 && (|lane1_IntFormatPlugin_logic_stages_0_hits));
  assign lane1_IntFormatPlugin_logic_stages_0_raw = early1_IntAluPlugin_logic_wb_payload;
  assign lane1_IntFormatPlugin_logic_stages_0_wb_payload = lane1_IntFormatPlugin_logic_stages_0_raw;
  assign lane1_IntFormatPlugin_logic_stages_1_hits = early1_BarrelShifterPlugin_logic_wb_valid;
  assign lane1_IntFormatPlugin_logic_stages_1_wb_valid = (toplevel_execute_ctrl3_up_LANE_SEL_lane1 && (|lane1_IntFormatPlugin_logic_stages_1_hits));
  assign lane1_IntFormatPlugin_logic_stages_1_raw = early1_BarrelShifterPlugin_logic_wb_payload;
  assign lane1_IntFormatPlugin_logic_stages_1_wb_payload = lane1_IntFormatPlugin_logic_stages_1_raw;
  assign lane1_IntFormatPlugin_logic_stages_2_hits = {late1_BarrelShifterPlugin_logic_wb_valid,late1_IntAluPlugin_logic_wb_valid};
  assign lane1_IntFormatPlugin_logic_stages_2_wb_valid = (toplevel_execute_ctrl4_up_LANE_SEL_lane1 && (|lane1_IntFormatPlugin_logic_stages_2_hits));
  assign lane1_IntFormatPlugin_logic_stages_2_raw = ((lane1_IntFormatPlugin_logic_stages_2_hits[0] ? late1_IntAluPlugin_logic_wb_payload : 32'h0) | (lane1_IntFormatPlugin_logic_stages_2_hits[1] ? late1_BarrelShifterPlugin_logic_wb_payload : 32'h0));
  assign lane1_IntFormatPlugin_logic_stages_2_wb_payload = lane1_IntFormatPlugin_logic_stages_2_raw;
  always @(*) begin
    _zz_toplevel_execute_ctrl3_down_late1_SrcPlugin_SRC1_lane1 = 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
    case(toplevel_execute_ctrl3_down_late1_SrcPlugin_logic_SRC1_CTRL_lane1)
      1'b0 : begin
        _zz_toplevel_execute_ctrl3_down_late1_SrcPlugin_SRC1_lane1 = toplevel_execute_ctrl3_down_integer_RS1_lane1;
      end
      default : begin
        _zz_toplevel_execute_ctrl3_down_late1_SrcPlugin_SRC1_lane1 = {toplevel_execute_ctrl3_down_Decode_UOP_lane1[31 : 12],12'h0};
      end
    endcase
  end

  assign toplevel_execute_ctrl3_down_late1_SrcPlugin_SRC1_lane1 = _zz_toplevel_execute_ctrl3_down_late1_SrcPlugin_SRC1_lane1;
  always @(*) begin
    _zz_toplevel_execute_ctrl3_down_late1_SrcPlugin_SRC2_lane1 = 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
    case(toplevel_execute_ctrl3_down_late1_SrcPlugin_logic_SRC2_CTRL_lane1)
      2'b00 : begin
        _zz_toplevel_execute_ctrl3_down_late1_SrcPlugin_SRC2_lane1 = toplevel_execute_ctrl3_down_integer_RS2_lane1;
      end
      2'b01 : begin
        _zz_toplevel_execute_ctrl3_down_late1_SrcPlugin_SRC2_lane1 = {{20{_zz__zz_toplevel_execute_ctrl3_down_late1_SrcPlugin_SRC2_lane1[11]}}, _zz__zz_toplevel_execute_ctrl3_down_late1_SrcPlugin_SRC2_lane1};
      end
      2'b10 : begin
        _zz_toplevel_execute_ctrl3_down_late1_SrcPlugin_SRC2_lane1 = toplevel_execute_ctrl3_down_PC_lane1;
      end
      default : begin
      end
    endcase
  end

  assign toplevel_execute_ctrl3_down_late1_SrcPlugin_SRC2_lane1 = _zz_toplevel_execute_ctrl3_down_late1_SrcPlugin_SRC2_lane1;
  always @(*) begin
    late1_SrcPlugin_logic_addsub_combined_rs2Patched = toplevel_execute_ctrl4_down_late1_SrcPlugin_SRC2_lane1;
    if(toplevel_execute_ctrl4_down_SrcStageables_REVERT_lane1) begin
      late1_SrcPlugin_logic_addsub_combined_rs2Patched = (~ toplevel_execute_ctrl4_down_late1_SrcPlugin_SRC2_lane1);
    end
    if(toplevel_execute_ctrl4_down_SrcStageables_ZERO_lane1) begin
      late1_SrcPlugin_logic_addsub_combined_rs2Patched = 32'h0;
    end
  end

  assign toplevel_execute_ctrl4_down_late1_SrcPlugin_ADD_SUB_lane1 = ($signed(_zz_toplevel_execute_ctrl4_down_late1_SrcPlugin_ADD_SUB_lane1) + $signed(_zz_toplevel_execute_ctrl4_down_late1_SrcPlugin_ADD_SUB_lane1_1));
  assign toplevel_execute_ctrl4_down_late1_SrcPlugin_LESS_lane1 = ((toplevel_execute_ctrl4_down_late1_SrcPlugin_SRC1_lane1[31] == toplevel_execute_ctrl4_down_late1_SrcPlugin_SRC2_lane1[31]) ? toplevel_execute_ctrl4_down_late1_SrcPlugin_ADD_SUB_lane1[31] : (toplevel_execute_ctrl4_down_SrcStageables_UNSIGNED_lane1 ? toplevel_execute_ctrl4_down_late1_SrcPlugin_SRC2_lane1[31] : toplevel_execute_ctrl4_down_late1_SrcPlugin_SRC1_lane1[31]));
  assign toplevel_execute_ctrl4_down_late0_BranchPlugin_logic_alu_EQ_lane0 = ($signed(toplevel_execute_ctrl4_down_late0_SrcPlugin_SRC1_lane0) == $signed(toplevel_execute_ctrl4_down_late0_SrcPlugin_SRC2_lane0));
  assign toplevel_execute_ctrl4_down_late0_BranchPlugin_logic_alu_btb_BAD_TARGET_lane0 = (toplevel_execute_ctrl4_down_Prediction_ALIGNED_JUMPED_PC_lane0 != toplevel_execute_ctrl4_down_early0_BranchPlugin_pcCalc_PC_TRUE_lane0);
  assign late0_BranchPlugin_logic_alu_expectedMsb = (MmuPlugin_api_fetchTranslationEnable ? _zz_late0_BranchPlugin_logic_alu_expectedMsb[31] : 1'b0);
  assign toplevel_execute_ctrl4_down_late0_BranchPlugin_logic_alu_MSB_FAILED_lane0 = ((toplevel_execute_ctrl4_down_BranchPlugin_BRANCH_CTRL_lane0 == BranchPlugin_BranchCtrlEnum_JALR) && 1'b0);
  assign switch_Misc_l241_2 = toplevel_execute_ctrl4_down_Decode_UOP_lane0[14 : 12];
  always @(*) begin
    casez(switch_Misc_l241_2)
      3'b000 : begin
        _zz_toplevel_execute_ctrl4_down_late0_BranchPlugin_logic_jumpLogic_COND_lane0 = toplevel_execute_ctrl4_down_late0_BranchPlugin_logic_alu_EQ_lane0;
      end
      3'b001 : begin
        _zz_toplevel_execute_ctrl4_down_late0_BranchPlugin_logic_jumpLogic_COND_lane0 = (! toplevel_execute_ctrl4_down_late0_BranchPlugin_logic_alu_EQ_lane0);
      end
      3'b1?1 : begin
        _zz_toplevel_execute_ctrl4_down_late0_BranchPlugin_logic_jumpLogic_COND_lane0 = (! toplevel_execute_ctrl4_down_late0_SrcPlugin_LESS_lane0);
      end
      default : begin
        _zz_toplevel_execute_ctrl4_down_late0_BranchPlugin_logic_jumpLogic_COND_lane0 = toplevel_execute_ctrl4_down_late0_SrcPlugin_LESS_lane0;
      end
    endcase
  end

  always @(*) begin
    case(toplevel_execute_ctrl4_down_BranchPlugin_BRANCH_CTRL_lane0)
      BranchPlugin_BranchCtrlEnum_JALR : begin
        _zz_toplevel_execute_ctrl4_down_late0_BranchPlugin_logic_jumpLogic_COND_lane0_1 = 1'b1;
      end
      BranchPlugin_BranchCtrlEnum_JAL : begin
        _zz_toplevel_execute_ctrl4_down_late0_BranchPlugin_logic_jumpLogic_COND_lane0_1 = 1'b1;
      end
      default : begin
        _zz_toplevel_execute_ctrl4_down_late0_BranchPlugin_logic_jumpLogic_COND_lane0_1 = _zz_toplevel_execute_ctrl4_down_late0_BranchPlugin_logic_jumpLogic_COND_lane0;
      end
    endcase
  end

  assign toplevel_execute_ctrl4_down_late0_BranchPlugin_logic_jumpLogic_COND_lane0 = _zz_toplevel_execute_ctrl4_down_late0_BranchPlugin_logic_jumpLogic_COND_lane0_1;
  assign toplevel_execute_ctrl4_down_late0_BranchPlugin_logic_jumpLogic_btb_REAL_TARGET_lane0 = (toplevel_execute_ctrl4_down_late0_BranchPlugin_logic_jumpLogic_COND_lane0 ? toplevel_execute_ctrl4_down_early0_BranchPlugin_pcCalc_PC_TRUE_lane0 : toplevel_execute_ctrl4_down_early0_BranchPlugin_pcCalc_PC_FALSE_lane0);
  assign late0_BranchPlugin_logic_jumpLogic_wrongCond = (toplevel_execute_ctrl4_down_Prediction_ALIGNED_JUMPED_lane0 != toplevel_execute_ctrl4_down_late0_BranchPlugin_logic_jumpLogic_COND_lane0);
  assign late0_BranchPlugin_logic_jumpLogic_needFix = ((late0_BranchPlugin_logic_jumpLogic_wrongCond || (toplevel_execute_ctrl4_down_late0_BranchPlugin_logic_jumpLogic_COND_lane0 && toplevel_execute_ctrl4_down_late0_BranchPlugin_logic_alu_btb_BAD_TARGET_lane0)) || toplevel_execute_ctrl4_down_late0_BranchPlugin_logic_alu_MSB_FAILED_lane0);
  assign late0_BranchPlugin_logic_jumpLogic_doIt = ((toplevel_execute_ctrl4_up_LANE_SEL_lane0 && toplevel_execute_ctrl4_down_late0_BranchPlugin_SEL_lane0) && late0_BranchPlugin_logic_jumpLogic_needFix);
  assign late0_BranchPlugin_logic_jumpLogic_history_fromFetch_slice = toplevel_execute_ctrl4_down_PC_lane0[2 : 1];
  assign late0_BranchPlugin_logic_jumpLogic_history_fromFetch_shifter = toplevel_execute_ctrl4_down_Prediction_BRANCH_HISTORY_lane0;
  assign when_BranchPlugin_l206_6 = ((late0_BranchPlugin_logic_jumpLogic_history_fromFetch_slice < 2'b00) && toplevel_execute_ctrl4_down_Prediction_ALIGNED_SLICES_BRANCH_lane0[0]);
  assign when_BranchPlugin_l206_7 = ((late0_BranchPlugin_logic_jumpLogic_history_fromFetch_slice < 2'b01) && toplevel_execute_ctrl4_down_Prediction_ALIGNED_SLICES_BRANCH_lane0[1]);
  assign when_BranchPlugin_l206_8 = ((late0_BranchPlugin_logic_jumpLogic_history_fromFetch_slice < 2'b10) && toplevel_execute_ctrl4_down_Prediction_ALIGNED_SLICES_BRANCH_lane0[2]);
  assign when_BranchPlugin_l210_2 = (toplevel_execute_ctrl4_down_BranchPlugin_BRANCH_CTRL_lane0 == BranchPlugin_BranchCtrlEnum_B);
  assign late0_BranchPlugin_logic_jumpLogic_history_next = late0_BranchPlugin_logic_jumpLogic_history_fromFetch_shifter_4;
  assign late0_BranchPlugin_logic_jumpLogic_history_fetched = toplevel_execute_ctrl4_down_Prediction_BRANCH_HISTORY_lane0;
  assign late0_BranchPlugin_logic_pcPort_valid = late0_BranchPlugin_logic_jumpLogic_doIt;
  assign late0_BranchPlugin_logic_pcPort_payload_fault = toplevel_execute_ctrl4_down_late0_BranchPlugin_logic_alu_MSB_FAILED_lane0;
  assign late0_BranchPlugin_logic_pcPort_payload_pc = toplevel_execute_ctrl4_down_late0_BranchPlugin_logic_jumpLogic_btb_REAL_TARGET_lane0;
  assign late0_BranchPlugin_logic_pcPort_payload_laneAge = toplevel_execute_ctrl4_down_LANE_AGE_lane0;
  assign late0_BranchPlugin_logic_historyPort_valid = late0_BranchPlugin_logic_jumpLogic_doIt;
  assign late0_BranchPlugin_logic_historyPort_payload_history = late0_BranchPlugin_logic_jumpLogic_history_next;
  assign late0_BranchPlugin_logic_historyPort_payload_age = toplevel_execute_ctrl4_down_LANE_AGE_lane0;
  assign late0_BranchPlugin_logic_flushPort_valid = late0_BranchPlugin_logic_jumpLogic_doIt;
  assign late0_BranchPlugin_logic_flushPort_payload_uopId = toplevel_execute_ctrl4_down_Decode_UOP_ID_lane0;
  assign late0_BranchPlugin_logic_flushPort_payload_laneAge = toplevel_execute_ctrl4_down_LANE_AGE_lane0;
  assign late0_BranchPlugin_logic_flushPort_payload_self = 1'b0;
  assign toplevel_execute_ctrl4_down_late0_BranchPlugin_logic_jumpLogic_MISSALIGNED_lane0 = ((toplevel_execute_ctrl4_down_early0_BranchPlugin_pcCalc_PC_TRUE_lane0[0 : 0] != 1'b0) && toplevel_execute_ctrl4_down_late0_BranchPlugin_logic_jumpLogic_COND_lane0);
  assign toplevel_execute_ctrl4_down_late0_BranchPlugin_logic_jumpLogic_IS_JAL_lane0 = (toplevel_execute_ctrl4_down_BranchPlugin_BRANCH_CTRL_lane0 == BranchPlugin_BranchCtrlEnum_JAL);
  assign toplevel_execute_ctrl4_down_late0_BranchPlugin_logic_jumpLogic_IS_JALR_lane0 = (toplevel_execute_ctrl4_down_BranchPlugin_BRANCH_CTRL_lane0 == BranchPlugin_BranchCtrlEnum_JALR);
  assign late0_BranchPlugin_logic_jumpLogic_rdLink = (|{(toplevel_execute_ctrl4_down_Decode_UOP_lane0[11 : 7] == 5'h05),(toplevel_execute_ctrl4_down_Decode_UOP_lane0[11 : 7] == 5'h01)});
  assign late0_BranchPlugin_logic_jumpLogic_rs1Link = (|{(toplevel_execute_ctrl4_down_Decode_UOP_lane0[19 : 15] == 5'h05),(toplevel_execute_ctrl4_down_Decode_UOP_lane0[19 : 15] == 5'h01)});
  assign late0_BranchPlugin_logic_jumpLogic_rdEquRs1 = (toplevel_execute_ctrl4_down_Decode_UOP_lane0[11 : 7] == toplevel_execute_ctrl4_down_Decode_UOP_lane0[19 : 15]);
  assign late0_BranchPlugin_logic_jumpLogic_learn_valid = (((toplevel_execute_ctrl4_up_LANE_SEL_lane0 && toplevel_execute_ctrl4_down_isReady) && (! toplevel_execute_lane0_ctrls_4_upIsCancel)) && (|{toplevel_execute_ctrl4_down_late0_BranchPlugin_SEL_lane0,toplevel_execute_ctrl4_down_early0_BranchPlugin_SEL_lane0}));
  assign late0_BranchPlugin_logic_jumpLogic_learn_payload_taken = toplevel_execute_ctrl4_down_late0_BranchPlugin_logic_jumpLogic_COND_lane0;
  assign late0_BranchPlugin_logic_jumpLogic_learn_payload_pcTarget = toplevel_execute_ctrl4_down_early0_BranchPlugin_pcCalc_PC_TRUE_lane0;
  assign late0_BranchPlugin_logic_jumpLogic_learn_payload_pcOnLastSlice = toplevel_execute_ctrl4_down_early0_BranchPlugin_pcCalc_PC_LAST_SLICE_lane0;
  assign late0_BranchPlugin_logic_jumpLogic_learn_payload_isBranch = (toplevel_execute_ctrl4_down_BranchPlugin_BRANCH_CTRL_lane0 == BranchPlugin_BranchCtrlEnum_B);
  assign late0_BranchPlugin_logic_jumpLogic_learn_payload_isPush = ((toplevel_execute_ctrl4_down_late0_BranchPlugin_logic_jumpLogic_IS_JAL_lane0 || toplevel_execute_ctrl4_down_late0_BranchPlugin_logic_jumpLogic_IS_JALR_lane0) && late0_BranchPlugin_logic_jumpLogic_rdLink);
  assign late0_BranchPlugin_logic_jumpLogic_learn_payload_isPop = (toplevel_execute_ctrl4_down_late0_BranchPlugin_logic_jumpLogic_IS_JALR_lane0 && (((! late0_BranchPlugin_logic_jumpLogic_rdLink) && late0_BranchPlugin_logic_jumpLogic_rs1Link) || ((late0_BranchPlugin_logic_jumpLogic_rdLink && late0_BranchPlugin_logic_jumpLogic_rs1Link) && (! late0_BranchPlugin_logic_jumpLogic_rdEquRs1))));
  assign late0_BranchPlugin_logic_jumpLogic_learn_payload_wasWrong = late0_BranchPlugin_logic_jumpLogic_needFix;
  assign late0_BranchPlugin_logic_jumpLogic_learn_payload_badPredictedTarget = toplevel_execute_ctrl4_down_late0_BranchPlugin_logic_alu_btb_BAD_TARGET_lane0;
  assign late0_BranchPlugin_logic_jumpLogic_learn_payload_history = late0_BranchPlugin_logic_jumpLogic_history_fetched;
  assign late0_BranchPlugin_logic_jumpLogic_learn_payload_uopId = toplevel_execute_ctrl4_down_Decode_UOP_ID_lane0;
  assign late0_BranchPlugin_logic_jumpLogic_learn_payload_ctx_GSharePlugin_GSHARE_COUNTER_0 = toplevel_execute_ctrl4_down_GSharePlugin_GSHARE_COUNTER_lane0_0;
  assign late0_BranchPlugin_logic_jumpLogic_learn_payload_ctx_GSharePlugin_GSHARE_COUNTER_1 = toplevel_execute_ctrl4_down_GSharePlugin_GSHARE_COUNTER_lane0_1;
  assign late0_BranchPlugin_logic_jumpLogic_learn_payload_ctx_GSharePlugin_GSHARE_COUNTER_2 = toplevel_execute_ctrl4_down_GSharePlugin_GSHARE_COUNTER_lane0_2;
  assign late0_BranchPlugin_logic_jumpLogic_learn_payload_ctx_GSharePlugin_GSHARE_COUNTER_3 = toplevel_execute_ctrl4_down_GSharePlugin_GSHARE_COUNTER_lane0_3;
  assign late0_BranchPlugin_logic_wb_valid = toplevel_execute_ctrl4_down_late0_BranchPlugin_SEL_lane0;
  assign late0_BranchPlugin_logic_wb_payload = toplevel_execute_ctrl4_down_early0_BranchPlugin_pcCalc_PC_FALSE_lane0;
  assign toplevel_execute_ctrl4_down_late1_BranchPlugin_logic_alu_EQ_lane1 = ($signed(toplevel_execute_ctrl4_down_late1_SrcPlugin_SRC1_lane1) == $signed(toplevel_execute_ctrl4_down_late1_SrcPlugin_SRC2_lane1));
  assign toplevel_execute_ctrl4_down_late1_BranchPlugin_logic_alu_btb_BAD_TARGET_lane1 = (toplevel_execute_ctrl4_down_Prediction_ALIGNED_JUMPED_PC_lane1 != toplevel_execute_ctrl4_down_early1_BranchPlugin_pcCalc_PC_TRUE_lane1);
  assign late1_BranchPlugin_logic_alu_expectedMsb = (MmuPlugin_api_fetchTranslationEnable ? _zz_late1_BranchPlugin_logic_alu_expectedMsb[31] : 1'b0);
  assign toplevel_execute_ctrl4_down_late1_BranchPlugin_logic_alu_MSB_FAILED_lane1 = ((toplevel_execute_ctrl4_down_BranchPlugin_BRANCH_CTRL_lane1 == BranchPlugin_BranchCtrlEnum_JALR) && 1'b0);
  assign switch_Misc_l241_3 = toplevel_execute_ctrl4_down_Decode_UOP_lane1[14 : 12];
  always @(*) begin
    casez(switch_Misc_l241_3)
      3'b000 : begin
        _zz_toplevel_execute_ctrl4_down_late1_BranchPlugin_logic_jumpLogic_COND_lane1 = toplevel_execute_ctrl4_down_late1_BranchPlugin_logic_alu_EQ_lane1;
      end
      3'b001 : begin
        _zz_toplevel_execute_ctrl4_down_late1_BranchPlugin_logic_jumpLogic_COND_lane1 = (! toplevel_execute_ctrl4_down_late1_BranchPlugin_logic_alu_EQ_lane1);
      end
      3'b1?1 : begin
        _zz_toplevel_execute_ctrl4_down_late1_BranchPlugin_logic_jumpLogic_COND_lane1 = (! toplevel_execute_ctrl4_down_late1_SrcPlugin_LESS_lane1);
      end
      default : begin
        _zz_toplevel_execute_ctrl4_down_late1_BranchPlugin_logic_jumpLogic_COND_lane1 = toplevel_execute_ctrl4_down_late1_SrcPlugin_LESS_lane1;
      end
    endcase
  end

  always @(*) begin
    case(toplevel_execute_ctrl4_down_BranchPlugin_BRANCH_CTRL_lane1)
      BranchPlugin_BranchCtrlEnum_JALR : begin
        _zz_toplevel_execute_ctrl4_down_late1_BranchPlugin_logic_jumpLogic_COND_lane1_1 = 1'b1;
      end
      BranchPlugin_BranchCtrlEnum_JAL : begin
        _zz_toplevel_execute_ctrl4_down_late1_BranchPlugin_logic_jumpLogic_COND_lane1_1 = 1'b1;
      end
      default : begin
        _zz_toplevel_execute_ctrl4_down_late1_BranchPlugin_logic_jumpLogic_COND_lane1_1 = _zz_toplevel_execute_ctrl4_down_late1_BranchPlugin_logic_jumpLogic_COND_lane1;
      end
    endcase
  end

  assign toplevel_execute_ctrl4_down_late1_BranchPlugin_logic_jumpLogic_COND_lane1 = _zz_toplevel_execute_ctrl4_down_late1_BranchPlugin_logic_jumpLogic_COND_lane1_1;
  assign toplevel_execute_ctrl4_down_late1_BranchPlugin_logic_jumpLogic_btb_REAL_TARGET_lane1 = (toplevel_execute_ctrl4_down_late1_BranchPlugin_logic_jumpLogic_COND_lane1 ? toplevel_execute_ctrl4_down_early1_BranchPlugin_pcCalc_PC_TRUE_lane1 : toplevel_execute_ctrl4_down_early1_BranchPlugin_pcCalc_PC_FALSE_lane1);
  assign late1_BranchPlugin_logic_jumpLogic_wrongCond = (toplevel_execute_ctrl4_down_Prediction_ALIGNED_JUMPED_lane1 != toplevel_execute_ctrl4_down_late1_BranchPlugin_logic_jumpLogic_COND_lane1);
  assign late1_BranchPlugin_logic_jumpLogic_needFix = ((late1_BranchPlugin_logic_jumpLogic_wrongCond || (toplevel_execute_ctrl4_down_late1_BranchPlugin_logic_jumpLogic_COND_lane1 && toplevel_execute_ctrl4_down_late1_BranchPlugin_logic_alu_btb_BAD_TARGET_lane1)) || toplevel_execute_ctrl4_down_late1_BranchPlugin_logic_alu_MSB_FAILED_lane1);
  assign late1_BranchPlugin_logic_jumpLogic_doIt = ((toplevel_execute_ctrl4_up_LANE_SEL_lane1 && toplevel_execute_ctrl4_down_late1_BranchPlugin_SEL_lane1) && late1_BranchPlugin_logic_jumpLogic_needFix);
  assign late1_BranchPlugin_logic_jumpLogic_history_fromFetch_slice = toplevel_execute_ctrl4_down_PC_lane1[2 : 1];
  assign late1_BranchPlugin_logic_jumpLogic_history_fromFetch_shifter = toplevel_execute_ctrl4_down_Prediction_BRANCH_HISTORY_lane1;
  assign when_BranchPlugin_l206_9 = ((late1_BranchPlugin_logic_jumpLogic_history_fromFetch_slice < 2'b00) && toplevel_execute_ctrl4_down_Prediction_ALIGNED_SLICES_BRANCH_lane1[0]);
  assign when_BranchPlugin_l206_10 = ((late1_BranchPlugin_logic_jumpLogic_history_fromFetch_slice < 2'b01) && toplevel_execute_ctrl4_down_Prediction_ALIGNED_SLICES_BRANCH_lane1[1]);
  assign when_BranchPlugin_l206_11 = ((late1_BranchPlugin_logic_jumpLogic_history_fromFetch_slice < 2'b10) && toplevel_execute_ctrl4_down_Prediction_ALIGNED_SLICES_BRANCH_lane1[2]);
  assign when_BranchPlugin_l210_3 = (toplevel_execute_ctrl4_down_BranchPlugin_BRANCH_CTRL_lane1 == BranchPlugin_BranchCtrlEnum_B);
  assign late1_BranchPlugin_logic_jumpLogic_history_next = late1_BranchPlugin_logic_jumpLogic_history_fromFetch_shifter_4;
  assign late1_BranchPlugin_logic_jumpLogic_history_fetched = toplevel_execute_ctrl4_down_Prediction_BRANCH_HISTORY_lane1;
  assign late1_BranchPlugin_logic_pcPort_valid = late1_BranchPlugin_logic_jumpLogic_doIt;
  assign late1_BranchPlugin_logic_pcPort_payload_fault = toplevel_execute_ctrl4_down_late1_BranchPlugin_logic_alu_MSB_FAILED_lane1;
  assign late1_BranchPlugin_logic_pcPort_payload_pc = toplevel_execute_ctrl4_down_late1_BranchPlugin_logic_jumpLogic_btb_REAL_TARGET_lane1;
  assign late1_BranchPlugin_logic_pcPort_payload_laneAge = toplevel_execute_ctrl4_down_LANE_AGE_lane1;
  assign late1_BranchPlugin_logic_historyPort_valid = late1_BranchPlugin_logic_jumpLogic_doIt;
  assign late1_BranchPlugin_logic_historyPort_payload_history = late1_BranchPlugin_logic_jumpLogic_history_next;
  assign late1_BranchPlugin_logic_historyPort_payload_age = toplevel_execute_ctrl4_down_LANE_AGE_lane1;
  assign late1_BranchPlugin_logic_flushPort_valid = late1_BranchPlugin_logic_jumpLogic_doIt;
  assign late1_BranchPlugin_logic_flushPort_payload_uopId = toplevel_execute_ctrl4_down_Decode_UOP_ID_lane1;
  assign late1_BranchPlugin_logic_flushPort_payload_laneAge = toplevel_execute_ctrl4_down_LANE_AGE_lane1;
  assign late1_BranchPlugin_logic_flushPort_payload_self = 1'b0;
  assign toplevel_execute_ctrl4_down_late1_BranchPlugin_logic_jumpLogic_MISSALIGNED_lane1 = ((toplevel_execute_ctrl4_down_early1_BranchPlugin_pcCalc_PC_TRUE_lane1[0 : 0] != 1'b0) && toplevel_execute_ctrl4_down_late1_BranchPlugin_logic_jumpLogic_COND_lane1);
  assign toplevel_execute_ctrl4_down_late1_BranchPlugin_logic_jumpLogic_IS_JAL_lane1 = (toplevel_execute_ctrl4_down_BranchPlugin_BRANCH_CTRL_lane1 == BranchPlugin_BranchCtrlEnum_JAL);
  assign toplevel_execute_ctrl4_down_late1_BranchPlugin_logic_jumpLogic_IS_JALR_lane1 = (toplevel_execute_ctrl4_down_BranchPlugin_BRANCH_CTRL_lane1 == BranchPlugin_BranchCtrlEnum_JALR);
  assign late1_BranchPlugin_logic_jumpLogic_rdLink = (|{(toplevel_execute_ctrl4_down_Decode_UOP_lane1[11 : 7] == 5'h05),(toplevel_execute_ctrl4_down_Decode_UOP_lane1[11 : 7] == 5'h01)});
  assign late1_BranchPlugin_logic_jumpLogic_rs1Link = (|{(toplevel_execute_ctrl4_down_Decode_UOP_lane1[19 : 15] == 5'h05),(toplevel_execute_ctrl4_down_Decode_UOP_lane1[19 : 15] == 5'h01)});
  assign late1_BranchPlugin_logic_jumpLogic_rdEquRs1 = (toplevel_execute_ctrl4_down_Decode_UOP_lane1[11 : 7] == toplevel_execute_ctrl4_down_Decode_UOP_lane1[19 : 15]);
  assign late1_BranchPlugin_logic_jumpLogic_learn_valid = (((toplevel_execute_ctrl4_up_LANE_SEL_lane1 && toplevel_execute_ctrl4_down_isReady) && (! toplevel_execute_lane1_ctrls_4_upIsCancel)) && (|{toplevel_execute_ctrl4_down_late1_BranchPlugin_SEL_lane1,toplevel_execute_ctrl4_down_early1_BranchPlugin_SEL_lane1}));
  assign late1_BranchPlugin_logic_jumpLogic_learn_payload_taken = toplevel_execute_ctrl4_down_late1_BranchPlugin_logic_jumpLogic_COND_lane1;
  assign late1_BranchPlugin_logic_jumpLogic_learn_payload_pcTarget = toplevel_execute_ctrl4_down_early1_BranchPlugin_pcCalc_PC_TRUE_lane1;
  assign late1_BranchPlugin_logic_jumpLogic_learn_payload_pcOnLastSlice = toplevel_execute_ctrl4_down_early1_BranchPlugin_pcCalc_PC_LAST_SLICE_lane1;
  assign late1_BranchPlugin_logic_jumpLogic_learn_payload_isBranch = (toplevel_execute_ctrl4_down_BranchPlugin_BRANCH_CTRL_lane1 == BranchPlugin_BranchCtrlEnum_B);
  assign late1_BranchPlugin_logic_jumpLogic_learn_payload_isPush = ((toplevel_execute_ctrl4_down_late1_BranchPlugin_logic_jumpLogic_IS_JAL_lane1 || toplevel_execute_ctrl4_down_late1_BranchPlugin_logic_jumpLogic_IS_JALR_lane1) && late1_BranchPlugin_logic_jumpLogic_rdLink);
  assign late1_BranchPlugin_logic_jumpLogic_learn_payload_isPop = (toplevel_execute_ctrl4_down_late1_BranchPlugin_logic_jumpLogic_IS_JALR_lane1 && (((! late1_BranchPlugin_logic_jumpLogic_rdLink) && late1_BranchPlugin_logic_jumpLogic_rs1Link) || ((late1_BranchPlugin_logic_jumpLogic_rdLink && late1_BranchPlugin_logic_jumpLogic_rs1Link) && (! late1_BranchPlugin_logic_jumpLogic_rdEquRs1))));
  assign late1_BranchPlugin_logic_jumpLogic_learn_payload_wasWrong = late1_BranchPlugin_logic_jumpLogic_needFix;
  assign late1_BranchPlugin_logic_jumpLogic_learn_payload_badPredictedTarget = toplevel_execute_ctrl4_down_late1_BranchPlugin_logic_alu_btb_BAD_TARGET_lane1;
  assign late1_BranchPlugin_logic_jumpLogic_learn_payload_history = late1_BranchPlugin_logic_jumpLogic_history_fetched;
  assign late1_BranchPlugin_logic_jumpLogic_learn_payload_uopId = toplevel_execute_ctrl4_down_Decode_UOP_ID_lane1;
  assign late1_BranchPlugin_logic_jumpLogic_learn_payload_ctx_GSharePlugin_GSHARE_COUNTER_0 = toplevel_execute_ctrl4_down_GSharePlugin_GSHARE_COUNTER_lane1_0;
  assign late1_BranchPlugin_logic_jumpLogic_learn_payload_ctx_GSharePlugin_GSHARE_COUNTER_1 = toplevel_execute_ctrl4_down_GSharePlugin_GSHARE_COUNTER_lane1_1;
  assign late1_BranchPlugin_logic_jumpLogic_learn_payload_ctx_GSharePlugin_GSHARE_COUNTER_2 = toplevel_execute_ctrl4_down_GSharePlugin_GSHARE_COUNTER_lane1_2;
  assign late1_BranchPlugin_logic_jumpLogic_learn_payload_ctx_GSharePlugin_GSHARE_COUNTER_3 = toplevel_execute_ctrl4_down_GSharePlugin_GSHARE_COUNTER_lane1_3;
  assign late1_BranchPlugin_logic_wb_valid = toplevel_execute_ctrl4_down_late1_BranchPlugin_SEL_lane1;
  assign late1_BranchPlugin_logic_wb_payload = toplevel_execute_ctrl4_down_early1_BranchPlugin_pcCalc_PC_FALSE_lane1;
  always @(*) begin
    late0_BranchPlugin_logic_jumpLogic_learn_ready = late0_BranchPlugin_logic_jumpLogic_learn_m2sPipe_ready;
    if(when_Stream_l393) begin
      late0_BranchPlugin_logic_jumpLogic_learn_ready = 1'b1;
    end
  end

  assign when_Stream_l393 = (! late0_BranchPlugin_logic_jumpLogic_learn_m2sPipe_valid);
  assign late0_BranchPlugin_logic_jumpLogic_learn_m2sPipe_valid = late0_BranchPlugin_logic_jumpLogic_learn_rValid;
  assign late0_BranchPlugin_logic_jumpLogic_learn_m2sPipe_payload_pcOnLastSlice = late0_BranchPlugin_logic_jumpLogic_learn_rData_pcOnLastSlice;
  assign late0_BranchPlugin_logic_jumpLogic_learn_m2sPipe_payload_pcTarget = late0_BranchPlugin_logic_jumpLogic_learn_rData_pcTarget;
  assign late0_BranchPlugin_logic_jumpLogic_learn_m2sPipe_payload_taken = late0_BranchPlugin_logic_jumpLogic_learn_rData_taken;
  assign late0_BranchPlugin_logic_jumpLogic_learn_m2sPipe_payload_isBranch = late0_BranchPlugin_logic_jumpLogic_learn_rData_isBranch;
  assign late0_BranchPlugin_logic_jumpLogic_learn_m2sPipe_payload_isPush = late0_BranchPlugin_logic_jumpLogic_learn_rData_isPush;
  assign late0_BranchPlugin_logic_jumpLogic_learn_m2sPipe_payload_isPop = late0_BranchPlugin_logic_jumpLogic_learn_rData_isPop;
  assign late0_BranchPlugin_logic_jumpLogic_learn_m2sPipe_payload_wasWrong = late0_BranchPlugin_logic_jumpLogic_learn_rData_wasWrong;
  assign late0_BranchPlugin_logic_jumpLogic_learn_m2sPipe_payload_badPredictedTarget = late0_BranchPlugin_logic_jumpLogic_learn_rData_badPredictedTarget;
  assign late0_BranchPlugin_logic_jumpLogic_learn_m2sPipe_payload_history = late0_BranchPlugin_logic_jumpLogic_learn_rData_history;
  assign late0_BranchPlugin_logic_jumpLogic_learn_m2sPipe_payload_uopId = late0_BranchPlugin_logic_jumpLogic_learn_rData_uopId;
  assign late0_BranchPlugin_logic_jumpLogic_learn_m2sPipe_payload_ctx_GSharePlugin_GSHARE_COUNTER_0 = late0_BranchPlugin_logic_jumpLogic_learn_rData_ctx_GSharePlugin_GSHARE_COUNTER_0;
  assign late0_BranchPlugin_logic_jumpLogic_learn_m2sPipe_payload_ctx_GSharePlugin_GSHARE_COUNTER_1 = late0_BranchPlugin_logic_jumpLogic_learn_rData_ctx_GSharePlugin_GSHARE_COUNTER_1;
  assign late0_BranchPlugin_logic_jumpLogic_learn_m2sPipe_payload_ctx_GSharePlugin_GSHARE_COUNTER_2 = late0_BranchPlugin_logic_jumpLogic_learn_rData_ctx_GSharePlugin_GSHARE_COUNTER_2;
  assign late0_BranchPlugin_logic_jumpLogic_learn_m2sPipe_payload_ctx_GSharePlugin_GSHARE_COUNTER_3 = late0_BranchPlugin_logic_jumpLogic_learn_rData_ctx_GSharePlugin_GSHARE_COUNTER_3;
  always @(*) begin
    late1_BranchPlugin_logic_jumpLogic_learn_ready = late1_BranchPlugin_logic_jumpLogic_learn_m2sPipe_ready;
    if(when_Stream_l393_1) begin
      late1_BranchPlugin_logic_jumpLogic_learn_ready = 1'b1;
    end
  end

  assign when_Stream_l393_1 = (! late1_BranchPlugin_logic_jumpLogic_learn_m2sPipe_valid);
  assign late1_BranchPlugin_logic_jumpLogic_learn_m2sPipe_valid = late1_BranchPlugin_logic_jumpLogic_learn_rValid;
  assign late1_BranchPlugin_logic_jumpLogic_learn_m2sPipe_payload_pcOnLastSlice = late1_BranchPlugin_logic_jumpLogic_learn_rData_pcOnLastSlice;
  assign late1_BranchPlugin_logic_jumpLogic_learn_m2sPipe_payload_pcTarget = late1_BranchPlugin_logic_jumpLogic_learn_rData_pcTarget;
  assign late1_BranchPlugin_logic_jumpLogic_learn_m2sPipe_payload_taken = late1_BranchPlugin_logic_jumpLogic_learn_rData_taken;
  assign late1_BranchPlugin_logic_jumpLogic_learn_m2sPipe_payload_isBranch = late1_BranchPlugin_logic_jumpLogic_learn_rData_isBranch;
  assign late1_BranchPlugin_logic_jumpLogic_learn_m2sPipe_payload_isPush = late1_BranchPlugin_logic_jumpLogic_learn_rData_isPush;
  assign late1_BranchPlugin_logic_jumpLogic_learn_m2sPipe_payload_isPop = late1_BranchPlugin_logic_jumpLogic_learn_rData_isPop;
  assign late1_BranchPlugin_logic_jumpLogic_learn_m2sPipe_payload_wasWrong = late1_BranchPlugin_logic_jumpLogic_learn_rData_wasWrong;
  assign late1_BranchPlugin_logic_jumpLogic_learn_m2sPipe_payload_badPredictedTarget = late1_BranchPlugin_logic_jumpLogic_learn_rData_badPredictedTarget;
  assign late1_BranchPlugin_logic_jumpLogic_learn_m2sPipe_payload_history = late1_BranchPlugin_logic_jumpLogic_learn_rData_history;
  assign late1_BranchPlugin_logic_jumpLogic_learn_m2sPipe_payload_uopId = late1_BranchPlugin_logic_jumpLogic_learn_rData_uopId;
  assign late1_BranchPlugin_logic_jumpLogic_learn_m2sPipe_payload_ctx_GSharePlugin_GSHARE_COUNTER_0 = late1_BranchPlugin_logic_jumpLogic_learn_rData_ctx_GSharePlugin_GSHARE_COUNTER_0;
  assign late1_BranchPlugin_logic_jumpLogic_learn_m2sPipe_payload_ctx_GSharePlugin_GSHARE_COUNTER_1 = late1_BranchPlugin_logic_jumpLogic_learn_rData_ctx_GSharePlugin_GSHARE_COUNTER_1;
  assign late1_BranchPlugin_logic_jumpLogic_learn_m2sPipe_payload_ctx_GSharePlugin_GSHARE_COUNTER_2 = late1_BranchPlugin_logic_jumpLogic_learn_rData_ctx_GSharePlugin_GSHARE_COUNTER_2;
  assign late1_BranchPlugin_logic_jumpLogic_learn_m2sPipe_payload_ctx_GSharePlugin_GSHARE_COUNTER_3 = late1_BranchPlugin_logic_jumpLogic_learn_rData_ctx_GSharePlugin_GSHARE_COUNTER_3;
  assign late0_BranchPlugin_logic_jumpLogic_learn_m2sPipe_ready = streamArbiter_10_io_inputs_0_ready;
  assign late1_BranchPlugin_logic_jumpLogic_learn_m2sPipe_ready = streamArbiter_10_io_inputs_1_ready;
  assign streamArbiter_10_io_output_combStage_valid = streamArbiter_10_io_output_valid;
  assign streamArbiter_10_io_output_combStage_payload_pcOnLastSlice = streamArbiter_10_io_output_payload_pcOnLastSlice;
  assign streamArbiter_10_io_output_combStage_payload_pcTarget = streamArbiter_10_io_output_payload_pcTarget;
  assign streamArbiter_10_io_output_combStage_payload_taken = streamArbiter_10_io_output_payload_taken;
  assign streamArbiter_10_io_output_combStage_payload_isBranch = streamArbiter_10_io_output_payload_isBranch;
  assign streamArbiter_10_io_output_combStage_payload_isPush = streamArbiter_10_io_output_payload_isPush;
  assign streamArbiter_10_io_output_combStage_payload_isPop = streamArbiter_10_io_output_payload_isPop;
  assign streamArbiter_10_io_output_combStage_payload_wasWrong = streamArbiter_10_io_output_payload_wasWrong;
  assign streamArbiter_10_io_output_combStage_payload_badPredictedTarget = streamArbiter_10_io_output_payload_badPredictedTarget;
  assign streamArbiter_10_io_output_combStage_payload_history = streamArbiter_10_io_output_payload_history;
  assign streamArbiter_10_io_output_combStage_payload_uopId = streamArbiter_10_io_output_payload_uopId;
  assign streamArbiter_10_io_output_combStage_payload_ctx_GSharePlugin_GSHARE_COUNTER_0 = streamArbiter_10_io_output_payload_ctx_GSharePlugin_GSHARE_COUNTER_0;
  assign streamArbiter_10_io_output_combStage_payload_ctx_GSharePlugin_GSHARE_COUNTER_1 = streamArbiter_10_io_output_payload_ctx_GSharePlugin_GSHARE_COUNTER_1;
  assign streamArbiter_10_io_output_combStage_payload_ctx_GSharePlugin_GSHARE_COUNTER_2 = streamArbiter_10_io_output_payload_ctx_GSharePlugin_GSHARE_COUNTER_2;
  assign streamArbiter_10_io_output_combStage_payload_ctx_GSharePlugin_GSHARE_COUNTER_3 = streamArbiter_10_io_output_payload_ctx_GSharePlugin_GSHARE_COUNTER_3;
  assign streamArbiter_10_io_output_combStage_ready = 1'b1;
  assign LearnPlugin_logic_learn_valid = streamArbiter_10_io_output_combStage_valid;
  assign LearnPlugin_logic_learn_payload_pcOnLastSlice = streamArbiter_10_io_output_combStage_payload_pcOnLastSlice;
  assign LearnPlugin_logic_learn_payload_pcTarget = streamArbiter_10_io_output_combStage_payload_pcTarget;
  assign LearnPlugin_logic_learn_payload_taken = streamArbiter_10_io_output_combStage_payload_taken;
  assign LearnPlugin_logic_learn_payload_isBranch = streamArbiter_10_io_output_combStage_payload_isBranch;
  assign LearnPlugin_logic_learn_payload_isPush = streamArbiter_10_io_output_combStage_payload_isPush;
  assign LearnPlugin_logic_learn_payload_isPop = streamArbiter_10_io_output_combStage_payload_isPop;
  assign LearnPlugin_logic_learn_payload_wasWrong = streamArbiter_10_io_output_combStage_payload_wasWrong;
  assign LearnPlugin_logic_learn_payload_badPredictedTarget = streamArbiter_10_io_output_combStage_payload_badPredictedTarget;
  assign LearnPlugin_logic_learn_payload_history = streamArbiter_10_io_output_combStage_payload_history;
  assign LearnPlugin_logic_learn_payload_uopId = streamArbiter_10_io_output_combStage_payload_uopId;
  assign LearnPlugin_logic_learn_payload_ctx_GSharePlugin_GSHARE_COUNTER_0 = streamArbiter_10_io_output_combStage_payload_ctx_GSharePlugin_GSHARE_COUNTER_0;
  assign LearnPlugin_logic_learn_payload_ctx_GSharePlugin_GSHARE_COUNTER_1 = streamArbiter_10_io_output_combStage_payload_ctx_GSharePlugin_GSHARE_COUNTER_1;
  assign LearnPlugin_logic_learn_payload_ctx_GSharePlugin_GSHARE_COUNTER_2 = streamArbiter_10_io_output_combStage_payload_ctx_GSharePlugin_GSHARE_COUNTER_2;
  assign LearnPlugin_logic_learn_payload_ctx_GSharePlugin_GSHARE_COUNTER_3 = streamArbiter_10_io_output_combStage_payload_ctx_GSharePlugin_GSHARE_COUNTER_3;
  assign toplevel_execute_ctrl2_COMPLETED_lane1_bypass = (toplevel_execute_ctrl2_up_COMPLETED_lane1 || toplevel_execute_ctrl2_down_COMPLETION_AT_2_lane1);
  assign toplevel_execute_ctrl3_COMPLETED_lane1_bypass = (toplevel_execute_ctrl3_up_COMPLETED_lane1 || toplevel_execute_ctrl3_down_COMPLETION_AT_3_lane1);
  assign toplevel_execute_ctrl4_COMPLETED_lane1_bypass = (toplevel_execute_ctrl4_up_COMPLETED_lane1 || toplevel_execute_ctrl4_down_COMPLETION_AT_4_lane1);
  assign execute_lane1_api_hartsInflight[0] = (|{(toplevel_execute_ctrl4_up_LANE_SEL_lane1 && 1'b1),{(toplevel_execute_ctrl3_up_LANE_SEL_lane1 && 1'b1),{(toplevel_execute_ctrl2_up_LANE_SEL_lane1 && 1'b1),(toplevel_execute_ctrl1_up_LANE_SEL_lane1 && 1'b1)}}});
  assign _zz_GSharePlugin_logic_onLearn_hash = LearnPlugin_logic_learn_payload_pcOnLastSlice[14 : 3];
  assign GSharePlugin_logic_onLearn_hash = ({_zz_GSharePlugin_logic_onLearn_hash[0],{_zz_GSharePlugin_logic_onLearn_hash[1],{_zz_GSharePlugin_logic_onLearn_hash[2],{_zz_GSharePlugin_logic_onLearn_hash[3],{_zz_GSharePlugin_logic_onLearn_hash[4],{_zz_GSharePlugin_logic_onLearn_hash[5],{_zz_GSharePlugin_logic_onLearn_hash_1,{_zz_GSharePlugin_logic_onLearn_hash_2,_zz_GSharePlugin_logic_onLearn_hash_3}}}}}}}} ^ LearnPlugin_logic_learn_payload_history);
  assign GSharePlugin_logic_onLearn_incrValue = (LearnPlugin_logic_learn_payload_taken ? 2'b01 : 2'b11);
  always @(*) begin
    GSharePlugin_logic_onLearn_overflow = 1'b0;
    if(when_GSharePlugin_l104) begin
      GSharePlugin_logic_onLearn_overflow = 1'b1;
    end
    if(when_GSharePlugin_l104_1) begin
      GSharePlugin_logic_onLearn_overflow = 1'b1;
    end
    if(when_GSharePlugin_l104_2) begin
      GSharePlugin_logic_onLearn_overflow = 1'b1;
    end
    if(when_GSharePlugin_l104_3) begin
      GSharePlugin_logic_onLearn_overflow = 1'b1;
    end
  end

  assign GSharePlugin_logic_onLearn_updated_0 = (LearnPlugin_logic_learn_payload_ctx_GSharePlugin_GSHARE_COUNTER_0 + ((LearnPlugin_logic_learn_payload_pcOnLastSlice[2 : 1] == 2'b00) ? GSharePlugin_logic_onLearn_incrValue : 2'b00));
  assign when_GSharePlugin_l104 = (((LearnPlugin_logic_learn_payload_taken && LearnPlugin_logic_learn_payload_ctx_GSharePlugin_GSHARE_COUNTER_0[1]) && (! GSharePlugin_logic_onLearn_updated_0[1])) || (((! LearnPlugin_logic_learn_payload_taken) && (! LearnPlugin_logic_learn_payload_ctx_GSharePlugin_GSHARE_COUNTER_0[1])) && GSharePlugin_logic_onLearn_updated_0[1]));
  assign GSharePlugin_logic_onLearn_updated_1 = (LearnPlugin_logic_learn_payload_ctx_GSharePlugin_GSHARE_COUNTER_1 + ((LearnPlugin_logic_learn_payload_pcOnLastSlice[2 : 1] == 2'b01) ? GSharePlugin_logic_onLearn_incrValue : 2'b00));
  assign when_GSharePlugin_l104_1 = (((LearnPlugin_logic_learn_payload_taken && LearnPlugin_logic_learn_payload_ctx_GSharePlugin_GSHARE_COUNTER_1[1]) && (! GSharePlugin_logic_onLearn_updated_1[1])) || (((! LearnPlugin_logic_learn_payload_taken) && (! LearnPlugin_logic_learn_payload_ctx_GSharePlugin_GSHARE_COUNTER_1[1])) && GSharePlugin_logic_onLearn_updated_1[1]));
  assign GSharePlugin_logic_onLearn_updated_2 = (LearnPlugin_logic_learn_payload_ctx_GSharePlugin_GSHARE_COUNTER_2 + ((LearnPlugin_logic_learn_payload_pcOnLastSlice[2 : 1] == 2'b10) ? GSharePlugin_logic_onLearn_incrValue : 2'b00));
  assign when_GSharePlugin_l104_2 = (((LearnPlugin_logic_learn_payload_taken && LearnPlugin_logic_learn_payload_ctx_GSharePlugin_GSHARE_COUNTER_2[1]) && (! GSharePlugin_logic_onLearn_updated_2[1])) || (((! LearnPlugin_logic_learn_payload_taken) && (! LearnPlugin_logic_learn_payload_ctx_GSharePlugin_GSHARE_COUNTER_2[1])) && GSharePlugin_logic_onLearn_updated_2[1]));
  assign GSharePlugin_logic_onLearn_updated_3 = (LearnPlugin_logic_learn_payload_ctx_GSharePlugin_GSHARE_COUNTER_3 + ((LearnPlugin_logic_learn_payload_pcOnLastSlice[2 : 1] == 2'b11) ? GSharePlugin_logic_onLearn_incrValue : 2'b00));
  assign when_GSharePlugin_l104_3 = (((LearnPlugin_logic_learn_payload_taken && LearnPlugin_logic_learn_payload_ctx_GSharePlugin_GSHARE_COUNTER_3[1]) && (! GSharePlugin_logic_onLearn_updated_3[1])) || (((! LearnPlugin_logic_learn_payload_taken) && (! LearnPlugin_logic_learn_payload_ctx_GSharePlugin_GSHARE_COUNTER_3[1])) && GSharePlugin_logic_onLearn_updated_3[1]));
  always @(*) begin
    GSharePlugin_logic_mem_write_valid = ((LearnPlugin_logic_learn_valid && LearnPlugin_logic_learn_payload_isBranch) && (! GSharePlugin_logic_onLearn_overflow));
    if(GSharePlugin_logic_initializer_busy) begin
      GSharePlugin_logic_mem_write_valid = 1'b1;
    end
  end

  always @(*) begin
    GSharePlugin_logic_mem_write_payload_address = GSharePlugin_logic_onLearn_hash;
    if(GSharePlugin_logic_initializer_busy) begin
      GSharePlugin_logic_mem_write_payload_address = GSharePlugin_logic_initializer_counter[11:0];
    end
  end

  always @(*) begin
    GSharePlugin_logic_mem_write_payload_data_0 = GSharePlugin_logic_onLearn_updated_0;
    if(GSharePlugin_logic_initializer_busy) begin
      GSharePlugin_logic_mem_write_payload_data_0 = _zz_GSharePlugin_logic_mem_write_payload_data_0[1 : 0];
    end
  end

  always @(*) begin
    GSharePlugin_logic_mem_write_payload_data_1 = GSharePlugin_logic_onLearn_updated_1;
    if(GSharePlugin_logic_initializer_busy) begin
      GSharePlugin_logic_mem_write_payload_data_1 = _zz_GSharePlugin_logic_mem_write_payload_data_0[3 : 2];
    end
  end

  always @(*) begin
    GSharePlugin_logic_mem_write_payload_data_2 = GSharePlugin_logic_onLearn_updated_2;
    if(GSharePlugin_logic_initializer_busy) begin
      GSharePlugin_logic_mem_write_payload_data_2 = _zz_GSharePlugin_logic_mem_write_payload_data_0[5 : 4];
    end
  end

  always @(*) begin
    GSharePlugin_logic_mem_write_payload_data_3 = GSharePlugin_logic_onLearn_updated_3;
    if(GSharePlugin_logic_initializer_busy) begin
      GSharePlugin_logic_mem_write_payload_data_3 = _zz_GSharePlugin_logic_mem_write_payload_data_0[7 : 6];
    end
  end

  assign GSharePlugin_logic_initializer_busy = (! GSharePlugin_logic_initializer_counter[12]);
  assign _zz_GSharePlugin_logic_mem_write_payload_data_0 = 8'h0;
  assign BtbPlugin_logic_onLearn_hash = LearnPlugin_logic_learn_payload_pcOnLastSlice[26 : 11];
  always @(*) begin
    BtbPlugin_logic_onLearn_port_valid = (LearnPlugin_logic_learn_valid && (LearnPlugin_logic_learn_payload_badPredictedTarget && LearnPlugin_logic_learn_payload_taken));
    if(DecoderPlugin_logic_forgetPort_valid) begin
      BtbPlugin_logic_onLearn_port_valid = DecoderPlugin_logic_forgetPort_valid;
    end
    if(BtbPlugin_logic_initializer_busy) begin
      BtbPlugin_logic_onLearn_port_valid = 1'b1;
    end
  end

  always @(*) begin
    BtbPlugin_logic_onLearn_port_payload_address = _zz_BtbPlugin_logic_onLearn_port_payload_address[7:0];
    if(DecoderPlugin_logic_forgetPort_valid) begin
      BtbPlugin_logic_onLearn_port_payload_address = _zz_BtbPlugin_logic_onLearn_port_payload_address_1[7:0];
    end
    if(BtbPlugin_logic_initializer_busy) begin
      BtbPlugin_logic_onLearn_port_payload_address = BtbPlugin_logic_initializer_counter[7:0];
    end
  end

  always @(*) begin
    BtbPlugin_logic_onLearn_port_payload_mask = (2'b01 <<< LearnPlugin_logic_learn_payload_pcOnLastSlice[2 : 2]);
    if(DecoderPlugin_logic_forgetPort_valid) begin
      BtbPlugin_logic_onLearn_port_payload_mask = (2'b01 <<< DecoderPlugin_logic_forgetPort_payload_pcOnLastSlice[2 : 2]);
    end
    if(BtbPlugin_logic_initializer_busy) begin
      BtbPlugin_logic_onLearn_port_payload_mask = 2'b11;
    end
  end

  always @(*) begin
    BtbPlugin_logic_onLearn_port_payload_data_0_hash = BtbPlugin_logic_onLearn_hash;
    if(DecoderPlugin_logic_forgetPort_valid) begin
      BtbPlugin_logic_onLearn_port_payload_data_0_hash = (~ BtbPlugin_logic_onForget_hash);
    end
    if(BtbPlugin_logic_initializer_busy) begin
      BtbPlugin_logic_onLearn_port_payload_data_0_hash = 16'hffff;
    end
  end

  always @(*) begin
    BtbPlugin_logic_onLearn_port_payload_data_0_sliceLow = LearnPlugin_logic_learn_payload_pcOnLastSlice[1 : 1];
    if(DecoderPlugin_logic_forgetPort_valid) begin
      BtbPlugin_logic_onLearn_port_payload_data_0_sliceLow = DecoderPlugin_logic_forgetPort_payload_pcOnLastSlice[1 : 1];
    end
    if(BtbPlugin_logic_initializer_busy) begin
      BtbPlugin_logic_onLearn_port_payload_data_0_sliceLow = 1'b0;
    end
  end

  assign BtbPlugin_logic_onLearn_port_payload_data_0_pcTarget = (LearnPlugin_logic_learn_payload_pcTarget >>> 1'd1);
  always @(*) begin
    BtbPlugin_logic_onLearn_port_payload_data_0_isBranch = LearnPlugin_logic_learn_payload_isBranch;
    if(DecoderPlugin_logic_forgetPort_valid) begin
      BtbPlugin_logic_onLearn_port_payload_data_0_isBranch = 1'b0;
    end
    if(BtbPlugin_logic_initializer_busy) begin
      BtbPlugin_logic_onLearn_port_payload_data_0_isBranch = 1'b0;
    end
  end

  always @(*) begin
    BtbPlugin_logic_onLearn_port_payload_data_0_isPush = LearnPlugin_logic_learn_payload_isPush;
    if(DecoderPlugin_logic_forgetPort_valid) begin
      BtbPlugin_logic_onLearn_port_payload_data_0_isPush = 1'b0;
    end
    if(BtbPlugin_logic_initializer_busy) begin
      BtbPlugin_logic_onLearn_port_payload_data_0_isPush = 1'b0;
    end
  end

  always @(*) begin
    BtbPlugin_logic_onLearn_port_payload_data_0_isPop = LearnPlugin_logic_learn_payload_isPop;
    if(DecoderPlugin_logic_forgetPort_valid) begin
      BtbPlugin_logic_onLearn_port_payload_data_0_isPop = 1'b0;
    end
    if(BtbPlugin_logic_initializer_busy) begin
      BtbPlugin_logic_onLearn_port_payload_data_0_isPop = 1'b0;
    end
  end

  always @(*) begin
    BtbPlugin_logic_onLearn_port_payload_data_1_hash = BtbPlugin_logic_onLearn_hash;
    if(DecoderPlugin_logic_forgetPort_valid) begin
      BtbPlugin_logic_onLearn_port_payload_data_1_hash = (~ BtbPlugin_logic_onForget_hash);
    end
    if(BtbPlugin_logic_initializer_busy) begin
      BtbPlugin_logic_onLearn_port_payload_data_1_hash = 16'hffff;
    end
  end

  always @(*) begin
    BtbPlugin_logic_onLearn_port_payload_data_1_sliceLow = LearnPlugin_logic_learn_payload_pcOnLastSlice[1 : 1];
    if(DecoderPlugin_logic_forgetPort_valid) begin
      BtbPlugin_logic_onLearn_port_payload_data_1_sliceLow = DecoderPlugin_logic_forgetPort_payload_pcOnLastSlice[1 : 1];
    end
    if(BtbPlugin_logic_initializer_busy) begin
      BtbPlugin_logic_onLearn_port_payload_data_1_sliceLow = 1'b0;
    end
  end

  assign BtbPlugin_logic_onLearn_port_payload_data_1_pcTarget = (LearnPlugin_logic_learn_payload_pcTarget >>> 1'd1);
  always @(*) begin
    BtbPlugin_logic_onLearn_port_payload_data_1_isBranch = LearnPlugin_logic_learn_payload_isBranch;
    if(DecoderPlugin_logic_forgetPort_valid) begin
      BtbPlugin_logic_onLearn_port_payload_data_1_isBranch = 1'b0;
    end
    if(BtbPlugin_logic_initializer_busy) begin
      BtbPlugin_logic_onLearn_port_payload_data_1_isBranch = 1'b0;
    end
  end

  always @(*) begin
    BtbPlugin_logic_onLearn_port_payload_data_1_isPush = LearnPlugin_logic_learn_payload_isPush;
    if(DecoderPlugin_logic_forgetPort_valid) begin
      BtbPlugin_logic_onLearn_port_payload_data_1_isPush = 1'b0;
    end
    if(BtbPlugin_logic_initializer_busy) begin
      BtbPlugin_logic_onLearn_port_payload_data_1_isPush = 1'b0;
    end
  end

  always @(*) begin
    BtbPlugin_logic_onLearn_port_payload_data_1_isPop = LearnPlugin_logic_learn_payload_isPop;
    if(DecoderPlugin_logic_forgetPort_valid) begin
      BtbPlugin_logic_onLearn_port_payload_data_1_isPop = 1'b0;
    end
    if(BtbPlugin_logic_initializer_busy) begin
      BtbPlugin_logic_onLearn_port_payload_data_1_isPop = 1'b0;
    end
  end

  assign toplevel_execute_ctrl2_COMPLETED_lane0_bypass = (toplevel_execute_ctrl2_up_COMPLETED_lane0 || toplevel_execute_ctrl2_down_COMPLETION_AT_2_lane0);
  assign toplevel_execute_ctrl3_COMPLETED_lane0_bypass = (toplevel_execute_ctrl3_up_COMPLETED_lane0 || toplevel_execute_ctrl3_down_COMPLETION_AT_3_lane0);
  assign toplevel_execute_ctrl4_COMPLETED_lane0_bypass = (toplevel_execute_ctrl4_up_COMPLETED_lane0 || toplevel_execute_ctrl4_down_COMPLETION_AT_4_lane0);
  assign execute_lane0_api_hartsInflight[0] = (|{(toplevel_execute_ctrl4_up_LANE_SEL_lane0 && 1'b1),{(toplevel_execute_ctrl3_up_LANE_SEL_lane0 && 1'b1),{(toplevel_execute_ctrl2_up_LANE_SEL_lane0 && 1'b1),(toplevel_execute_ctrl1_up_LANE_SEL_lane0 && 1'b1)}}});
  assign when_DecoderPlugin_l135 = (toplevel_decode_ctrls_1_up_isMoving && 1'b1);
  assign DecoderPlugin_logic_interrupt_async = PrivilegedPlugin_logic_harts_0_int_pending;
  assign when_DecoderPlugin_l143 = (((! toplevel_decode_ctrls_1_up_valid) || toplevel_decode_ctrls_1_up_ready) || toplevel_decode_ctrls_1_up_isCanceling);
  assign _zz_toplevel_decode_ctrls_1_down_DispatchPlugin_MAY_FLUSH_0 = ((toplevel_decode_ctrls_1_down_Decode_INSTRUCTION_0 & 32'h00000018) == 32'h0);
  assign toplevel_decode_ctrls_1_down_RS1_ENABLE_0 = _zz_toplevel_decode_ctrls_1_down_RS1_ENABLE_0[0];
  assign toplevel_decode_ctrls_1_down_RS1_PHYS_0 = toplevel_decode_ctrls_1_down_Decode_INSTRUCTION_0[19 : 15];
  assign toplevel_decode_ctrls_1_down_RS2_ENABLE_0 = _zz_toplevel_decode_ctrls_1_down_RS2_ENABLE_0[0];
  assign toplevel_decode_ctrls_1_down_RS2_PHYS_0 = toplevel_decode_ctrls_1_down_Decode_INSTRUCTION_0[24 : 20];
  assign _zz_toplevel_decode_ctrls_1_down_DispatchPlugin_logic_LANES_LAYER_HIT_0_0 = ((toplevel_decode_ctrls_1_down_Decode_INSTRUCTION_0 & 32'h0000000c) == 32'h00000004);
  assign _zz_toplevel_decode_ctrls_1_down_DispatchPlugin_logic_LANES_LAYER_HIT_3_0 = ((toplevel_decode_ctrls_1_down_Decode_INSTRUCTION_0 & 32'h00000048) == 32'h00000048);
  always @(*) begin
    toplevel_decode_ctrls_1_down_RD_ENABLE_0 = _zz_toplevel_decode_ctrls_1_down_RD_ENABLE_0[0];
    if(when_DecoderPlugin_l234) begin
      toplevel_decode_ctrls_1_down_RD_ENABLE_0 = 1'b0;
    end
  end

  assign toplevel_decode_ctrls_1_down_RD_PHYS_0 = toplevel_decode_ctrls_1_down_Decode_INSTRUCTION_0[11 : 7];
  assign toplevel_decode_ctrls_1_down_Decode_LEGAL_0 = ((|{((toplevel_decode_ctrls_1_down_Decode_INSTRUCTION_0 & 32'h0000005f) == 32'h00000017),{((toplevel_decode_ctrls_1_down_Decode_INSTRUCTION_0 & 32'h0000007f) == 32'h0000006f),{((toplevel_decode_ctrls_1_down_Decode_INSTRUCTION_0 & _zz_toplevel_decode_ctrls_1_down_Decode_LEGAL_0) == 32'h00001073),{(_zz_toplevel_decode_ctrls_1_down_Decode_LEGAL_0_1 == _zz_toplevel_decode_ctrls_1_down_Decode_LEGAL_0_2),{_zz_toplevel_decode_ctrls_1_down_Decode_LEGAL_0_3,{_zz_toplevel_decode_ctrls_1_down_Decode_LEGAL_0_4,_zz_toplevel_decode_ctrls_1_down_Decode_LEGAL_0_5}}}}}}) && (! toplevel_decode_ctrls_1_down_Decode_DECOMPRESSION_FAULT_0));
  assign DecoderPlugin_logic_laneLogic_0_interruptPending = DecoderPlugin_logic_interrupt_buffered[0];
  always @(*) begin
    DecoderPlugin_logic_laneLogic_0_trapPort_valid = 1'b0;
    if(when_DecoderPlugin_l216) begin
      DecoderPlugin_logic_laneLogic_0_trapPort_valid = ((! toplevel_decode_ctrls_1_up_TRAP_0) || DecoderPlugin_logic_laneLogic_0_interruptPending);
      if(DecoderPlugin_logic_laneLogic_0_fixer_doIt) begin
        DecoderPlugin_logic_laneLogic_0_trapPort_valid = 1'b1;
      end
    end
  end

  always @(*) begin
    DecoderPlugin_logic_laneLogic_0_trapPort_payload_exception = 1'b1;
    if(DecoderPlugin_logic_laneLogic_0_fixer_doIt) begin
      DecoderPlugin_logic_laneLogic_0_trapPort_payload_exception = 1'b0;
    end
    if(DecoderPlugin_logic_laneLogic_0_interruptPending) begin
      DecoderPlugin_logic_laneLogic_0_trapPort_payload_exception = 1'b0;
    end
  end

  assign DecoderPlugin_logic_laneLogic_0_trapPort_payload_tval = toplevel_decode_ctrls_1_down_Decode_INSTRUCTION_RAW_0;
  always @(*) begin
    DecoderPlugin_logic_laneLogic_0_trapPort_payload_code = 4'b0010;
    if(DecoderPlugin_logic_laneLogic_0_fixer_doIt) begin
      DecoderPlugin_logic_laneLogic_0_trapPort_payload_code = 4'b0100;
    end
    if(DecoderPlugin_logic_laneLogic_0_interruptPending) begin
      DecoderPlugin_logic_laneLogic_0_trapPort_payload_code = 4'b0000;
    end
  end

  assign DecoderPlugin_logic_laneLogic_0_trapPort_payload_laneAge = 2'b00;
  assign DecoderPlugin_logic_laneLogic_0_trapPort_payload_arg = 3'b000;
  assign _zz_toplevel_decode_ctrls_1_down_DispatchPlugin_logic_LANES_LAYER_HIT_0_0_1 = ((toplevel_decode_ctrls_1_down_Decode_INSTRUCTION_0 & 32'h00000050) == 32'h00000040);
  assign DecoderPlugin_logic_laneLogic_0_fixer_isJb = _zz_DecoderPlugin_logic_laneLogic_0_fixer_isJb[0];
  assign DecoderPlugin_logic_laneLogic_0_fixer_doIt = (toplevel_decode_ctrls_1_up_LANE_SEL_0 && ((toplevel_decode_ctrls_1_down_Prediction_ALIGNED_JUMPED_0 && (! DecoderPlugin_logic_laneLogic_0_fixer_isJb)) || toplevel_decode_ctrls_1_down_Prediction_ALIGN_REDO_0));
  assign when_CtrlLaneApi_l46_2 = (toplevel_decode_ctrls_1_up_isReady || toplevel_decode_ctrls_1_lane0_upIsCancel);
  assign DecoderPlugin_logic_laneLogic_0_completionPort_valid = ((toplevel_decode_ctrls_1_up_LANE_SEL_0 && toplevel_decode_ctrls_1_down_TRAP_0) && (toplevel_decode_ctrls_1_up_LANE_SEL_0 && (! toplevel_decode_ctrls_1_up_LANE_SEL_0_regNext)));
  assign DecoderPlugin_logic_laneLogic_0_completionPort_payload_uopId = toplevel_decode_ctrls_1_down_Decode_UOP_ID_0;
  assign DecoderPlugin_logic_laneLogic_0_completionPort_payload_trap = 1'b1;
  assign DecoderPlugin_logic_laneLogic_0_completionPort_payload_commit = 1'b0;
  assign when_DecoderPlugin_l216 = (toplevel_decode_ctrls_1_up_LANE_SEL_0 && (((! toplevel_decode_ctrls_1_down_Decode_LEGAL_0) || DecoderPlugin_logic_laneLogic_0_interruptPending) || DecoderPlugin_logic_laneLogic_0_fixer_doIt));
  assign DecoderPlugin_logic_laneLogic_0_flushPort_valid = (toplevel_decode_ctrls_1_up_LANE_SEL_0 && toplevel_decode_ctrls_1_down_TRAP_0);
  assign DecoderPlugin_logic_laneLogic_0_flushPort_payload_uopId = toplevel_decode_ctrls_1_down_Decode_UOP_ID_0;
  assign DecoderPlugin_logic_laneLogic_0_flushPort_payload_laneAge = 1'b0;
  assign DecoderPlugin_logic_laneLogic_0_flushPort_payload_self = 1'b0;
  assign when_DecoderPlugin_l234 = ((toplevel_decode_ctrls_1_down_Decode_INSTRUCTION_0[11 : 7] == 5'h0) && (|1'b1));
  assign toplevel_decode_ctrls_1_down_Decode_UOP_0 = toplevel_decode_ctrls_1_down_Decode_INSTRUCTION_0;
  assign DecoderPlugin_logic_laneLogic_0_uopIdBase = DecoderPlugin_logic_harts_0_uopId;
  assign toplevel_decode_ctrls_1_down_Decode_UOP_ID_0 = (DecoderPlugin_logic_laneLogic_0_uopIdBase + 16'h0);
  assign _zz_toplevel_decode_ctrls_1_down_DispatchPlugin_MAY_FLUSH_1 = ((toplevel_decode_ctrls_1_down_Decode_INSTRUCTION_1 & 32'h00000018) == 32'h0);
  assign toplevel_decode_ctrls_1_down_RS1_ENABLE_1 = _zz_toplevel_decode_ctrls_1_down_RS1_ENABLE_1[0];
  assign toplevel_decode_ctrls_1_down_RS1_PHYS_1 = toplevel_decode_ctrls_1_down_Decode_INSTRUCTION_1[19 : 15];
  assign toplevel_decode_ctrls_1_down_RS2_ENABLE_1 = _zz_toplevel_decode_ctrls_1_down_RS2_ENABLE_1[0];
  assign toplevel_decode_ctrls_1_down_RS2_PHYS_1 = toplevel_decode_ctrls_1_down_Decode_INSTRUCTION_1[24 : 20];
  assign _zz_toplevel_decode_ctrls_1_down_DispatchPlugin_logic_LANES_LAYER_HIT_0_1 = ((toplevel_decode_ctrls_1_down_Decode_INSTRUCTION_1 & 32'h0000000c) == 32'h00000004);
  assign _zz_toplevel_decode_ctrls_1_down_DispatchPlugin_logic_LANES_LAYER_HIT_3_1 = ((toplevel_decode_ctrls_1_down_Decode_INSTRUCTION_1 & 32'h00000048) == 32'h00000048);
  always @(*) begin
    toplevel_decode_ctrls_1_down_RD_ENABLE_1 = _zz_toplevel_decode_ctrls_1_down_RD_ENABLE_1[0];
    if(when_DecoderPlugin_l234_1) begin
      toplevel_decode_ctrls_1_down_RD_ENABLE_1 = 1'b0;
    end
  end

  assign toplevel_decode_ctrls_1_down_RD_PHYS_1 = toplevel_decode_ctrls_1_down_Decode_INSTRUCTION_1[11 : 7];
  assign toplevel_decode_ctrls_1_down_Decode_LEGAL_1 = ((|{((toplevel_decode_ctrls_1_down_Decode_INSTRUCTION_1 & 32'h0000005f) == 32'h00000017),{((toplevel_decode_ctrls_1_down_Decode_INSTRUCTION_1 & 32'h0000007f) == 32'h0000006f),{((toplevel_decode_ctrls_1_down_Decode_INSTRUCTION_1 & _zz_toplevel_decode_ctrls_1_down_Decode_LEGAL_1) == 32'h00001073),{(_zz_toplevel_decode_ctrls_1_down_Decode_LEGAL_1_1 == _zz_toplevel_decode_ctrls_1_down_Decode_LEGAL_1_2),{_zz_toplevel_decode_ctrls_1_down_Decode_LEGAL_1_3,{_zz_toplevel_decode_ctrls_1_down_Decode_LEGAL_1_4,_zz_toplevel_decode_ctrls_1_down_Decode_LEGAL_1_5}}}}}}) && (! toplevel_decode_ctrls_1_down_Decode_DECOMPRESSION_FAULT_1));
  assign DecoderPlugin_logic_laneLogic_1_interruptPending = DecoderPlugin_logic_interrupt_buffered[0];
  always @(*) begin
    DecoderPlugin_logic_laneLogic_1_trapPort_valid = 1'b0;
    if(when_DecoderPlugin_l216_1) begin
      DecoderPlugin_logic_laneLogic_1_trapPort_valid = ((! toplevel_decode_ctrls_1_up_TRAP_1) || DecoderPlugin_logic_laneLogic_1_interruptPending);
      if(DecoderPlugin_logic_laneLogic_1_fixer_doIt) begin
        DecoderPlugin_logic_laneLogic_1_trapPort_valid = 1'b1;
      end
    end
  end

  always @(*) begin
    DecoderPlugin_logic_laneLogic_1_trapPort_payload_exception = 1'b1;
    if(DecoderPlugin_logic_laneLogic_1_fixer_doIt) begin
      DecoderPlugin_logic_laneLogic_1_trapPort_payload_exception = 1'b0;
    end
    if(DecoderPlugin_logic_laneLogic_1_interruptPending) begin
      DecoderPlugin_logic_laneLogic_1_trapPort_payload_exception = 1'b0;
    end
  end

  assign DecoderPlugin_logic_laneLogic_1_trapPort_payload_tval = toplevel_decode_ctrls_1_down_Decode_INSTRUCTION_RAW_1;
  always @(*) begin
    DecoderPlugin_logic_laneLogic_1_trapPort_payload_code = 4'b0010;
    if(DecoderPlugin_logic_laneLogic_1_fixer_doIt) begin
      DecoderPlugin_logic_laneLogic_1_trapPort_payload_code = 4'b0100;
    end
    if(DecoderPlugin_logic_laneLogic_1_interruptPending) begin
      DecoderPlugin_logic_laneLogic_1_trapPort_payload_code = 4'b0000;
    end
  end

  assign DecoderPlugin_logic_laneLogic_1_trapPort_payload_laneAge = 2'b01;
  assign DecoderPlugin_logic_laneLogic_1_trapPort_payload_arg = 3'b000;
  assign _zz_toplevel_decode_ctrls_1_down_DispatchPlugin_logic_LANES_LAYER_HIT_0_1_1 = ((toplevel_decode_ctrls_1_down_Decode_INSTRUCTION_1 & 32'h00000050) == 32'h00000040);
  assign DecoderPlugin_logic_laneLogic_1_fixer_isJb = _zz_DecoderPlugin_logic_laneLogic_1_fixer_isJb[0];
  assign DecoderPlugin_logic_laneLogic_1_fixer_doIt = (toplevel_decode_ctrls_1_up_LANE_SEL_1 && ((toplevel_decode_ctrls_1_down_Prediction_ALIGNED_JUMPED_1 && (! DecoderPlugin_logic_laneLogic_1_fixer_isJb)) || toplevel_decode_ctrls_1_down_Prediction_ALIGN_REDO_1));
  assign when_CtrlLaneApi_l46_3 = (toplevel_decode_ctrls_1_up_isReady || toplevel_decode_ctrls_1_lane1_upIsCancel);
  assign DecoderPlugin_logic_laneLogic_1_completionPort_valid = ((toplevel_decode_ctrls_1_up_LANE_SEL_1 && toplevel_decode_ctrls_1_down_TRAP_1) && (toplevel_decode_ctrls_1_up_LANE_SEL_1 && (! toplevel_decode_ctrls_1_up_LANE_SEL_1_regNext)));
  assign DecoderPlugin_logic_laneLogic_1_completionPort_payload_uopId = toplevel_decode_ctrls_1_down_Decode_UOP_ID_1;
  assign DecoderPlugin_logic_laneLogic_1_completionPort_payload_trap = 1'b1;
  assign DecoderPlugin_logic_laneLogic_1_completionPort_payload_commit = 1'b0;
  assign when_DecoderPlugin_l216_1 = (toplevel_decode_ctrls_1_up_LANE_SEL_1 && (((! toplevel_decode_ctrls_1_down_Decode_LEGAL_1) || DecoderPlugin_logic_laneLogic_1_interruptPending) || DecoderPlugin_logic_laneLogic_1_fixer_doIt));
  assign DecoderPlugin_logic_laneLogic_1_flushPort_valid = (toplevel_decode_ctrls_1_up_LANE_SEL_1 && toplevel_decode_ctrls_1_down_TRAP_1);
  assign DecoderPlugin_logic_laneLogic_1_flushPort_payload_uopId = toplevel_decode_ctrls_1_down_Decode_UOP_ID_1;
  assign DecoderPlugin_logic_laneLogic_1_flushPort_payload_laneAge = 1'b1;
  assign DecoderPlugin_logic_laneLogic_1_flushPort_payload_self = 1'b0;
  assign when_DecoderPlugin_l234_1 = ((toplevel_decode_ctrls_1_down_Decode_INSTRUCTION_1[11 : 7] == 5'h0) && (|1'b1));
  assign toplevel_decode_ctrls_1_down_Decode_UOP_1 = toplevel_decode_ctrls_1_down_Decode_INSTRUCTION_1;
  assign DecoderPlugin_logic_laneLogic_1_uopIdBase = DecoderPlugin_logic_harts_0_uopId;
  assign toplevel_decode_ctrls_1_down_Decode_UOP_ID_1 = (DecoderPlugin_logic_laneLogic_1_uopIdBase + 16'h0001);
  assign _zz_CsrRamPlugin_csrMapper_ramAddress = CsrAccessPlugin_bus_decode_address;
  assign CsrRamPlugin_csrMapper_ramAddress = {(|((_zz_CsrRamPlugin_csrMapper_ramAddress & 12'h200) == 12'h200)),{(|{((_zz_CsrRamPlugin_csrMapper_ramAddress & _zz_CsrRamPlugin_csrMapper_ramAddress_1) == 12'h002),((_zz_CsrRamPlugin_csrMapper_ramAddress & _zz_CsrRamPlugin_csrMapper_ramAddress_2) == 12'h0)}),(|((_zz_CsrRamPlugin_csrMapper_ramAddress & 12'h003) == 12'h001))}};
  always @(*) begin
    CsrRamPlugin_csrMapper_withRead = 1'b0;
    if(when_CsrAccessPlugin_l264) begin
      CsrRamPlugin_csrMapper_withRead = 1'b1;
    end
  end

  assign CsrRamPlugin_csrMapper_read_valid = (CsrRamPlugin_csrMapper_withRead && (! CsrRamPlugin_api_holdRead));
  assign CsrRamPlugin_csrMapper_read_address = CsrRamPlugin_csrMapper_ramAddress;
  assign when_CsrRamPlugin_l77 = (CsrRamPlugin_csrMapper_withRead && (! CsrRamPlugin_csrMapper_read_ready));
  always @(*) begin
    CsrRamPlugin_csrMapper_doWrite = 1'b0;
    if(when_CsrAccessPlugin_l356_2) begin
      CsrRamPlugin_csrMapper_doWrite = 1'b1;
    end
  end

  assign when_CsrRamPlugin_l84 = (CsrRamPlugin_csrMapper_write_valid && CsrRamPlugin_csrMapper_write_ready);
  assign CsrRamPlugin_csrMapper_write_valid = ((CsrRamPlugin_csrMapper_doWrite && (! CsrRamPlugin_csrMapper_fired)) && (! CsrRamPlugin_api_holdWrite));
  assign CsrRamPlugin_csrMapper_write_address = CsrRamPlugin_csrMapper_ramAddress;
  assign CsrRamPlugin_csrMapper_write_data = CsrAccessPlugin_bus_write_bits;
  assign when_CsrRamPlugin_l88 = ((CsrRamPlugin_csrMapper_doWrite && (! CsrRamPlugin_csrMapper_fired)) && (! CsrRamPlugin_csrMapper_write_ready));
  assign lane0_integer_WriteBackPlugin_logic_stages_0_hits = {lane0_IntFormatPlugin_logic_stages_0_wb_valid,early0_BranchPlugin_logic_wb_valid};
  assign lane0_integer_WriteBackPlugin_logic_stages_0_muxed = ((lane0_integer_WriteBackPlugin_logic_stages_0_hits[0] ? early0_BranchPlugin_logic_wb_payload : 32'h0) | (lane0_integer_WriteBackPlugin_logic_stages_0_hits[1] ? lane0_IntFormatPlugin_logic_stages_0_wb_payload : 32'h0));
  assign toplevel_execute_ctrl2_lane0_integer_WriteBackPlugin_logic_DATA_lane0_bypass = lane0_integer_WriteBackPlugin_logic_stages_0_muxed;
  assign lane0_integer_WriteBackPlugin_logic_stages_0_write_valid = (((((toplevel_execute_ctrl2_down_LANE_SEL_lane0 && toplevel_execute_ctrl2_down_isReady) && (! toplevel_execute_lane0_ctrls_2_downIsCancel)) && (|lane0_integer_WriteBackPlugin_logic_stages_0_hits)) && toplevel_execute_ctrl2_up_RD_ENABLE_lane0) && toplevel_execute_ctrl2_down_COMMIT_lane0);
  assign lane0_integer_WriteBackPlugin_logic_stages_0_write_payload_uopId = toplevel_execute_ctrl2_down_Decode_UOP_ID_lane0;
  assign lane0_integer_WriteBackPlugin_logic_stages_0_write_payload_data = lane0_integer_WriteBackPlugin_logic_stages_0_muxed;
  assign lane0_integer_WriteBackPlugin_logic_stages_1_hits = lane0_IntFormatPlugin_logic_stages_1_wb_valid;
  assign lane0_integer_WriteBackPlugin_logic_stages_1_muxed = (lane0_integer_WriteBackPlugin_logic_stages_1_hits[0] ? lane0_IntFormatPlugin_logic_stages_1_wb_payload : 32'h0);
  assign lane0_integer_WriteBackPlugin_logic_stages_1_merged = (toplevel_execute_ctrl3_up_lane0_integer_WriteBackPlugin_logic_DATA_lane0 | lane0_integer_WriteBackPlugin_logic_stages_1_muxed);
  assign toplevel_execute_ctrl3_lane0_integer_WriteBackPlugin_logic_DATA_lane0_bypass = lane0_integer_WriteBackPlugin_logic_stages_1_merged;
  assign lane0_integer_WriteBackPlugin_logic_stages_1_write_valid = (((((toplevel_execute_ctrl3_down_LANE_SEL_lane0 && toplevel_execute_ctrl3_down_isReady) && (! toplevel_execute_lane0_ctrls_3_downIsCancel)) && (|lane0_integer_WriteBackPlugin_logic_stages_1_hits)) && toplevel_execute_ctrl3_up_RD_ENABLE_lane0) && toplevel_execute_ctrl3_down_COMMIT_lane0);
  assign lane0_integer_WriteBackPlugin_logic_stages_1_write_payload_uopId = toplevel_execute_ctrl3_down_Decode_UOP_ID_lane0;
  assign lane0_integer_WriteBackPlugin_logic_stages_1_write_payload_data = lane0_integer_WriteBackPlugin_logic_stages_1_muxed;
  assign lane0_integer_WriteBackPlugin_logic_stages_2_hits = {lane0_IntFormatPlugin_logic_stages_2_wb_valid,late0_BranchPlugin_logic_wb_valid};
  assign lane0_integer_WriteBackPlugin_logic_stages_2_muxed = ((lane0_integer_WriteBackPlugin_logic_stages_2_hits[0] ? late0_BranchPlugin_logic_wb_payload : 32'h0) | (lane0_integer_WriteBackPlugin_logic_stages_2_hits[1] ? lane0_IntFormatPlugin_logic_stages_2_wb_payload : 32'h0));
  assign lane0_integer_WriteBackPlugin_logic_stages_2_merged = (toplevel_execute_ctrl4_up_lane0_integer_WriteBackPlugin_logic_DATA_lane0 | lane0_integer_WriteBackPlugin_logic_stages_2_muxed);
  assign toplevel_execute_ctrl4_lane0_integer_WriteBackPlugin_logic_DATA_lane0_bypass = lane0_integer_WriteBackPlugin_logic_stages_2_merged;
  assign lane0_integer_WriteBackPlugin_logic_stages_2_write_valid = (((((toplevel_execute_ctrl4_down_LANE_SEL_lane0 && toplevel_execute_ctrl4_down_isReady) && (! toplevel_execute_lane0_ctrls_4_downIsCancel)) && (|lane0_integer_WriteBackPlugin_logic_stages_2_hits)) && toplevel_execute_ctrl4_up_RD_ENABLE_lane0) && toplevel_execute_ctrl4_down_COMMIT_lane0);
  assign lane0_integer_WriteBackPlugin_logic_stages_2_write_payload_uopId = toplevel_execute_ctrl4_down_Decode_UOP_ID_lane0;
  assign lane0_integer_WriteBackPlugin_logic_stages_2_write_payload_data = lane0_integer_WriteBackPlugin_logic_stages_2_muxed;
  assign lane0_integer_WriteBackPlugin_logic_write_port_valid = (((((toplevel_execute_ctrl4_up_LANE_SEL_lane0 && toplevel_execute_ctrl4_down_isReady) && (! toplevel_execute_lane0_ctrls_4_upIsCancel)) && toplevel_execute_ctrl4_up_RD_ENABLE_lane0) && toplevel_execute_ctrl4_down_lane0_integer_WriteBackPlugin_SEL_lane0) && toplevel_execute_ctrl4_down_COMMIT_lane0);
  assign lane0_integer_WriteBackPlugin_logic_write_port_address = toplevel_execute_ctrl4_down_RD_PHYS_lane0;
  assign lane0_integer_WriteBackPlugin_logic_write_port_data = toplevel_execute_ctrl4_down_lane0_integer_WriteBackPlugin_logic_DATA_lane0;
  assign lane0_integer_WriteBackPlugin_logic_write_port_uopId = toplevel_execute_ctrl4_down_Decode_UOP_ID_lane0;
  assign lane1_integer_WriteBackPlugin_logic_stages_0_hits = {lane1_IntFormatPlugin_logic_stages_0_wb_valid,early1_BranchPlugin_logic_wb_valid};
  assign lane1_integer_WriteBackPlugin_logic_stages_0_muxed = ((lane1_integer_WriteBackPlugin_logic_stages_0_hits[0] ? early1_BranchPlugin_logic_wb_payload : 32'h0) | (lane1_integer_WriteBackPlugin_logic_stages_0_hits[1] ? lane1_IntFormatPlugin_logic_stages_0_wb_payload : 32'h0));
  assign toplevel_execute_ctrl2_lane1_integer_WriteBackPlugin_logic_DATA_lane1_bypass = lane1_integer_WriteBackPlugin_logic_stages_0_muxed;
  assign lane1_integer_WriteBackPlugin_logic_stages_0_write_valid = (((((toplevel_execute_ctrl2_down_LANE_SEL_lane1 && toplevel_execute_ctrl2_down_isReady) && (! toplevel_execute_lane1_ctrls_2_downIsCancel)) && (|lane1_integer_WriteBackPlugin_logic_stages_0_hits)) && toplevel_execute_ctrl2_up_RD_ENABLE_lane1) && toplevel_execute_ctrl2_down_COMMIT_lane1);
  assign lane1_integer_WriteBackPlugin_logic_stages_0_write_payload_uopId = toplevel_execute_ctrl2_down_Decode_UOP_ID_lane1;
  assign lane1_integer_WriteBackPlugin_logic_stages_0_write_payload_data = lane1_integer_WriteBackPlugin_logic_stages_0_muxed;
  assign lane1_integer_WriteBackPlugin_logic_stages_1_hits = lane1_IntFormatPlugin_logic_stages_1_wb_valid;
  assign lane1_integer_WriteBackPlugin_logic_stages_1_muxed = (lane1_integer_WriteBackPlugin_logic_stages_1_hits[0] ? lane1_IntFormatPlugin_logic_stages_1_wb_payload : 32'h0);
  assign lane1_integer_WriteBackPlugin_logic_stages_1_merged = (toplevel_execute_ctrl3_up_lane1_integer_WriteBackPlugin_logic_DATA_lane1 | lane1_integer_WriteBackPlugin_logic_stages_1_muxed);
  assign toplevel_execute_ctrl3_lane1_integer_WriteBackPlugin_logic_DATA_lane1_bypass = lane1_integer_WriteBackPlugin_logic_stages_1_merged;
  assign lane1_integer_WriteBackPlugin_logic_stages_1_write_valid = (((((toplevel_execute_ctrl3_down_LANE_SEL_lane1 && toplevel_execute_ctrl3_down_isReady) && (! toplevel_execute_lane1_ctrls_3_downIsCancel)) && (|lane1_integer_WriteBackPlugin_logic_stages_1_hits)) && toplevel_execute_ctrl3_up_RD_ENABLE_lane1) && toplevel_execute_ctrl3_down_COMMIT_lane1);
  assign lane1_integer_WriteBackPlugin_logic_stages_1_write_payload_uopId = toplevel_execute_ctrl3_down_Decode_UOP_ID_lane1;
  assign lane1_integer_WriteBackPlugin_logic_stages_1_write_payload_data = lane1_integer_WriteBackPlugin_logic_stages_1_muxed;
  assign lane1_integer_WriteBackPlugin_logic_stages_2_hits = {lane1_IntFormatPlugin_logic_stages_2_wb_valid,late1_BranchPlugin_logic_wb_valid};
  assign lane1_integer_WriteBackPlugin_logic_stages_2_muxed = ((lane1_integer_WriteBackPlugin_logic_stages_2_hits[0] ? late1_BranchPlugin_logic_wb_payload : 32'h0) | (lane1_integer_WriteBackPlugin_logic_stages_2_hits[1] ? lane1_IntFormatPlugin_logic_stages_2_wb_payload : 32'h0));
  assign lane1_integer_WriteBackPlugin_logic_stages_2_merged = (toplevel_execute_ctrl4_up_lane1_integer_WriteBackPlugin_logic_DATA_lane1 | lane1_integer_WriteBackPlugin_logic_stages_2_muxed);
  assign toplevel_execute_ctrl4_lane1_integer_WriteBackPlugin_logic_DATA_lane1_bypass = lane1_integer_WriteBackPlugin_logic_stages_2_merged;
  assign lane1_integer_WriteBackPlugin_logic_stages_2_write_valid = (((((toplevel_execute_ctrl4_down_LANE_SEL_lane1 && toplevel_execute_ctrl4_down_isReady) && (! toplevel_execute_lane1_ctrls_4_downIsCancel)) && (|lane1_integer_WriteBackPlugin_logic_stages_2_hits)) && toplevel_execute_ctrl4_up_RD_ENABLE_lane1) && toplevel_execute_ctrl4_down_COMMIT_lane1);
  assign lane1_integer_WriteBackPlugin_logic_stages_2_write_payload_uopId = toplevel_execute_ctrl4_down_Decode_UOP_ID_lane1;
  assign lane1_integer_WriteBackPlugin_logic_stages_2_write_payload_data = lane1_integer_WriteBackPlugin_logic_stages_2_muxed;
  assign lane1_integer_WriteBackPlugin_logic_write_port_valid = (((((toplevel_execute_ctrl4_up_LANE_SEL_lane1 && toplevel_execute_ctrl4_down_isReady) && (! toplevel_execute_lane1_ctrls_4_upIsCancel)) && toplevel_execute_ctrl4_up_RD_ENABLE_lane1) && toplevel_execute_ctrl4_down_lane1_integer_WriteBackPlugin_SEL_lane1) && toplevel_execute_ctrl4_down_COMMIT_lane1);
  assign lane1_integer_WriteBackPlugin_logic_write_port_address = toplevel_execute_ctrl4_down_RD_PHYS_lane1;
  assign lane1_integer_WriteBackPlugin_logic_write_port_data = toplevel_execute_ctrl4_down_lane1_integer_WriteBackPlugin_logic_DATA_lane1;
  assign lane1_integer_WriteBackPlugin_logic_write_port_uopId = toplevel_execute_ctrl4_down_Decode_UOP_ID_lane1;
  assign DispatchPlugin_logic_trapPendings[0] = (|(DispatchPlugin_logic_slots_0_ctx_valid && DispatchPlugin_logic_slots_0_ctx_hm_TRAP));
  assign DispatchPlugin_logic_candidates_0_moving = (((! DispatchPlugin_logic_candidates_0_ctx_valid) || DispatchPlugin_logic_candidates_0_fire) || DispatchPlugin_logic_candidates_0_cancel);
  assign DispatchPlugin_logic_candidates_1_moving = (((! DispatchPlugin_logic_candidates_1_ctx_valid) || DispatchPlugin_logic_candidates_1_fire) || DispatchPlugin_logic_candidates_1_cancel);
  assign DispatchPlugin_logic_candidates_2_moving = (((! DispatchPlugin_logic_candidates_2_ctx_valid) || DispatchPlugin_logic_candidates_2_fire) || DispatchPlugin_logic_candidates_2_cancel);
  assign DispatchPlugin_logic_candidates_0_age = 1'b0;
  assign DispatchPlugin_logic_candidates_1_age = _zz_DispatchPlugin_logic_candidates_1_age;
  assign DispatchPlugin_logic_candidates_2_age = _zz_DispatchPlugin_logic_candidates_2_age[0:0];
  assign DispatchPlugin_logic_rsHazardChecker_0_onLl_0_onRs_0_hazard = (DispatchPlugin_logic_candidates_0_ctx_hm_RS1_ENABLE && (|{((((DispatchPlugin_logic_candidates_0_ctx_hm_DispatchPlugin_logic_hcs_0_onRs_0_ENABLES_0 && toplevel_execute_ctrl2_up_RD_ENABLE_lane1) && (toplevel_execute_ctrl2_up_RD_PHYS_lane1 == DispatchPlugin_logic_candidates_0_ctx_hm_RS1_PHYS)) && 1'b1) && (! toplevel_execute_ctrl2_down_BYPASSED_AT_3_lane1)),{(((_zz_DispatchPlugin_logic_rsHazardChecker_0_onLl_0_onRs_0_hazard && _zz_DispatchPlugin_logic_rsHazardChecker_0_onLl_0_onRs_0_hazard_1) && 1'b1) && (! toplevel_execute_ctrl1_down_BYPASSED_AT_2_lane1)),{((_zz_DispatchPlugin_logic_rsHazardChecker_0_onLl_0_onRs_0_hazard_2 && _zz_DispatchPlugin_logic_rsHazardChecker_0_onLl_0_onRs_0_hazard_3) && (! toplevel_execute_ctrl2_down_BYPASSED_AT_3_lane0)),((_zz_DispatchPlugin_logic_rsHazardChecker_0_onLl_0_onRs_0_hazard_4 && _zz_DispatchPlugin_logic_rsHazardChecker_0_onLl_0_onRs_0_hazard_5) && (! toplevel_execute_ctrl1_down_BYPASSED_AT_2_lane0))}}}));
  assign DispatchPlugin_logic_rsHazardChecker_0_onLl_0_onRs_1_hazard = (DispatchPlugin_logic_candidates_0_ctx_hm_RS2_ENABLE && (|{((((DispatchPlugin_logic_candidates_0_ctx_hm_DispatchPlugin_logic_hcs_0_onRs_1_ENABLES_0 && toplevel_execute_ctrl2_up_RD_ENABLE_lane1) && (toplevel_execute_ctrl2_up_RD_PHYS_lane1 == DispatchPlugin_logic_candidates_0_ctx_hm_RS2_PHYS)) && 1'b1) && (! toplevel_execute_ctrl2_down_BYPASSED_AT_3_lane1)),{(((_zz_DispatchPlugin_logic_rsHazardChecker_0_onLl_0_onRs_1_hazard && _zz_DispatchPlugin_logic_rsHazardChecker_0_onLl_0_onRs_1_hazard_1) && 1'b1) && (! toplevel_execute_ctrl1_down_BYPASSED_AT_2_lane1)),{((_zz_DispatchPlugin_logic_rsHazardChecker_0_onLl_0_onRs_1_hazard_2 && _zz_DispatchPlugin_logic_rsHazardChecker_0_onLl_0_onRs_1_hazard_3) && (! toplevel_execute_ctrl2_down_BYPASSED_AT_3_lane0)),((_zz_DispatchPlugin_logic_rsHazardChecker_0_onLl_0_onRs_1_hazard_4 && _zz_DispatchPlugin_logic_rsHazardChecker_0_onLl_0_onRs_1_hazard_5) && (! toplevel_execute_ctrl1_down_BYPASSED_AT_2_lane0))}}}));
  always @(*) begin
    DispatchPlugin_logic_candidates_0_rsHazards[0] = (|{DispatchPlugin_logic_rsHazardChecker_0_onLl_0_onRs_1_hazard,DispatchPlugin_logic_rsHazardChecker_0_onLl_0_onRs_0_hazard});
    DispatchPlugin_logic_candidates_0_rsHazards[1] = (|{DispatchPlugin_logic_rsHazardChecker_0_onLl_1_onRs_1_hazard,DispatchPlugin_logic_rsHazardChecker_0_onLl_1_onRs_0_hazard});
    DispatchPlugin_logic_candidates_0_rsHazards[2] = (|{DispatchPlugin_logic_rsHazardChecker_0_onLl_2_onRs_1_hazard,DispatchPlugin_logic_rsHazardChecker_0_onLl_2_onRs_0_hazard});
    DispatchPlugin_logic_candidates_0_rsHazards[3] = (|{DispatchPlugin_logic_rsHazardChecker_0_onLl_3_onRs_1_hazard,DispatchPlugin_logic_rsHazardChecker_0_onLl_3_onRs_0_hazard});
  end

  assign DispatchPlugin_logic_rsHazardChecker_0_onLl_1_onRs_0_hazard = (DispatchPlugin_logic_candidates_0_ctx_hm_RS1_ENABLE && (|{((((DispatchPlugin_logic_candidates_0_ctx_hm_DispatchPlugin_logic_hcs_1_onRs_0_ENABLES_0 && toplevel_execute_ctrl2_up_RD_ENABLE_lane1) && (toplevel_execute_ctrl2_up_RD_PHYS_lane1 == DispatchPlugin_logic_candidates_0_ctx_hm_RS1_PHYS)) && 1'b1) && (! toplevel_execute_ctrl2_down_BYPASSED_AT_3_lane1)),{(((_zz_DispatchPlugin_logic_rsHazardChecker_0_onLl_1_onRs_0_hazard && _zz_DispatchPlugin_logic_rsHazardChecker_0_onLl_1_onRs_0_hazard_1) && 1'b1) && (! toplevel_execute_ctrl1_down_BYPASSED_AT_2_lane1)),{((_zz_DispatchPlugin_logic_rsHazardChecker_0_onLl_1_onRs_0_hazard_2 && _zz_DispatchPlugin_logic_rsHazardChecker_0_onLl_1_onRs_0_hazard_3) && (! toplevel_execute_ctrl2_down_BYPASSED_AT_3_lane0)),((_zz_DispatchPlugin_logic_rsHazardChecker_0_onLl_1_onRs_0_hazard_4 && _zz_DispatchPlugin_logic_rsHazardChecker_0_onLl_1_onRs_0_hazard_5) && (! toplevel_execute_ctrl1_down_BYPASSED_AT_2_lane0))}}}));
  assign DispatchPlugin_logic_rsHazardChecker_0_onLl_1_onRs_1_hazard = (DispatchPlugin_logic_candidates_0_ctx_hm_RS2_ENABLE && (|{((((DispatchPlugin_logic_candidates_0_ctx_hm_DispatchPlugin_logic_hcs_1_onRs_1_ENABLES_0 && toplevel_execute_ctrl2_up_RD_ENABLE_lane1) && (toplevel_execute_ctrl2_up_RD_PHYS_lane1 == DispatchPlugin_logic_candidates_0_ctx_hm_RS2_PHYS)) && 1'b1) && (! toplevel_execute_ctrl2_down_BYPASSED_AT_3_lane1)),{(((_zz_DispatchPlugin_logic_rsHazardChecker_0_onLl_1_onRs_1_hazard && _zz_DispatchPlugin_logic_rsHazardChecker_0_onLl_1_onRs_1_hazard_1) && 1'b1) && (! toplevel_execute_ctrl1_down_BYPASSED_AT_2_lane1)),{((_zz_DispatchPlugin_logic_rsHazardChecker_0_onLl_1_onRs_1_hazard_2 && _zz_DispatchPlugin_logic_rsHazardChecker_0_onLl_1_onRs_1_hazard_3) && (! toplevel_execute_ctrl2_down_BYPASSED_AT_3_lane0)),((_zz_DispatchPlugin_logic_rsHazardChecker_0_onLl_1_onRs_1_hazard_4 && _zz_DispatchPlugin_logic_rsHazardChecker_0_onLl_1_onRs_1_hazard_5) && (! toplevel_execute_ctrl1_down_BYPASSED_AT_2_lane0))}}}));
  assign DispatchPlugin_logic_rsHazardChecker_0_onLl_2_onRs_0_hazard = (DispatchPlugin_logic_candidates_0_ctx_hm_RS1_ENABLE && 1'b0);
  assign DispatchPlugin_logic_rsHazardChecker_0_onLl_2_onRs_1_hazard = (DispatchPlugin_logic_candidates_0_ctx_hm_RS2_ENABLE && 1'b0);
  assign DispatchPlugin_logic_rsHazardChecker_0_onLl_3_onRs_0_hazard = (DispatchPlugin_logic_candidates_0_ctx_hm_RS1_ENABLE && 1'b0);
  assign DispatchPlugin_logic_rsHazardChecker_0_onLl_3_onRs_1_hazard = (DispatchPlugin_logic_candidates_0_ctx_hm_RS2_ENABLE && 1'b0);
  assign DispatchPlugin_logic_rsHazardChecker_1_onLl_0_onRs_0_hazard = (DispatchPlugin_logic_candidates_1_ctx_hm_RS1_ENABLE && (|{((((DispatchPlugin_logic_candidates_1_ctx_hm_DispatchPlugin_logic_hcs_0_onRs_0_ENABLES_0 && toplevel_execute_ctrl2_up_RD_ENABLE_lane1) && (toplevel_execute_ctrl2_up_RD_PHYS_lane1 == DispatchPlugin_logic_candidates_1_ctx_hm_RS1_PHYS)) && 1'b1) && (! toplevel_execute_ctrl2_down_BYPASSED_AT_3_lane1)),{(((_zz_DispatchPlugin_logic_rsHazardChecker_1_onLl_0_onRs_0_hazard && _zz_DispatchPlugin_logic_rsHazardChecker_1_onLl_0_onRs_0_hazard_1) && 1'b1) && (! toplevel_execute_ctrl1_down_BYPASSED_AT_2_lane1)),{((_zz_DispatchPlugin_logic_rsHazardChecker_1_onLl_0_onRs_0_hazard_2 && _zz_DispatchPlugin_logic_rsHazardChecker_1_onLl_0_onRs_0_hazard_3) && (! toplevel_execute_ctrl2_down_BYPASSED_AT_3_lane0)),((_zz_DispatchPlugin_logic_rsHazardChecker_1_onLl_0_onRs_0_hazard_4 && _zz_DispatchPlugin_logic_rsHazardChecker_1_onLl_0_onRs_0_hazard_5) && (! toplevel_execute_ctrl1_down_BYPASSED_AT_2_lane0))}}}));
  assign DispatchPlugin_logic_rsHazardChecker_1_onLl_0_onRs_1_hazard = (DispatchPlugin_logic_candidates_1_ctx_hm_RS2_ENABLE && (|{((((DispatchPlugin_logic_candidates_1_ctx_hm_DispatchPlugin_logic_hcs_0_onRs_1_ENABLES_0 && toplevel_execute_ctrl2_up_RD_ENABLE_lane1) && (toplevel_execute_ctrl2_up_RD_PHYS_lane1 == DispatchPlugin_logic_candidates_1_ctx_hm_RS2_PHYS)) && 1'b1) && (! toplevel_execute_ctrl2_down_BYPASSED_AT_3_lane1)),{(((_zz_DispatchPlugin_logic_rsHazardChecker_1_onLl_0_onRs_1_hazard && _zz_DispatchPlugin_logic_rsHazardChecker_1_onLl_0_onRs_1_hazard_1) && 1'b1) && (! toplevel_execute_ctrl1_down_BYPASSED_AT_2_lane1)),{((_zz_DispatchPlugin_logic_rsHazardChecker_1_onLl_0_onRs_1_hazard_2 && _zz_DispatchPlugin_logic_rsHazardChecker_1_onLl_0_onRs_1_hazard_3) && (! toplevel_execute_ctrl2_down_BYPASSED_AT_3_lane0)),((_zz_DispatchPlugin_logic_rsHazardChecker_1_onLl_0_onRs_1_hazard_4 && _zz_DispatchPlugin_logic_rsHazardChecker_1_onLl_0_onRs_1_hazard_5) && (! toplevel_execute_ctrl1_down_BYPASSED_AT_2_lane0))}}}));
  always @(*) begin
    DispatchPlugin_logic_candidates_1_rsHazards[0] = (|{DispatchPlugin_logic_rsHazardChecker_1_onLl_0_onRs_1_hazard,DispatchPlugin_logic_rsHazardChecker_1_onLl_0_onRs_0_hazard});
    DispatchPlugin_logic_candidates_1_rsHazards[1] = (|{DispatchPlugin_logic_rsHazardChecker_1_onLl_1_onRs_1_hazard,DispatchPlugin_logic_rsHazardChecker_1_onLl_1_onRs_0_hazard});
    DispatchPlugin_logic_candidates_1_rsHazards[2] = (|{DispatchPlugin_logic_rsHazardChecker_1_onLl_2_onRs_1_hazard,DispatchPlugin_logic_rsHazardChecker_1_onLl_2_onRs_0_hazard});
    DispatchPlugin_logic_candidates_1_rsHazards[3] = (|{DispatchPlugin_logic_rsHazardChecker_1_onLl_3_onRs_1_hazard,DispatchPlugin_logic_rsHazardChecker_1_onLl_3_onRs_0_hazard});
  end

  assign DispatchPlugin_logic_rsHazardChecker_1_onLl_1_onRs_0_hazard = (DispatchPlugin_logic_candidates_1_ctx_hm_RS1_ENABLE && (|{((((DispatchPlugin_logic_candidates_1_ctx_hm_DispatchPlugin_logic_hcs_1_onRs_0_ENABLES_0 && toplevel_execute_ctrl2_up_RD_ENABLE_lane1) && (toplevel_execute_ctrl2_up_RD_PHYS_lane1 == DispatchPlugin_logic_candidates_1_ctx_hm_RS1_PHYS)) && 1'b1) && (! toplevel_execute_ctrl2_down_BYPASSED_AT_3_lane1)),{(((_zz_DispatchPlugin_logic_rsHazardChecker_1_onLl_1_onRs_0_hazard && _zz_DispatchPlugin_logic_rsHazardChecker_1_onLl_1_onRs_0_hazard_1) && 1'b1) && (! toplevel_execute_ctrl1_down_BYPASSED_AT_2_lane1)),{((_zz_DispatchPlugin_logic_rsHazardChecker_1_onLl_1_onRs_0_hazard_2 && _zz_DispatchPlugin_logic_rsHazardChecker_1_onLl_1_onRs_0_hazard_3) && (! toplevel_execute_ctrl2_down_BYPASSED_AT_3_lane0)),((_zz_DispatchPlugin_logic_rsHazardChecker_1_onLl_1_onRs_0_hazard_4 && _zz_DispatchPlugin_logic_rsHazardChecker_1_onLl_1_onRs_0_hazard_5) && (! toplevel_execute_ctrl1_down_BYPASSED_AT_2_lane0))}}}));
  assign DispatchPlugin_logic_rsHazardChecker_1_onLl_1_onRs_1_hazard = (DispatchPlugin_logic_candidates_1_ctx_hm_RS2_ENABLE && (|{((((DispatchPlugin_logic_candidates_1_ctx_hm_DispatchPlugin_logic_hcs_1_onRs_1_ENABLES_0 && toplevel_execute_ctrl2_up_RD_ENABLE_lane1) && (toplevel_execute_ctrl2_up_RD_PHYS_lane1 == DispatchPlugin_logic_candidates_1_ctx_hm_RS2_PHYS)) && 1'b1) && (! toplevel_execute_ctrl2_down_BYPASSED_AT_3_lane1)),{(((_zz_DispatchPlugin_logic_rsHazardChecker_1_onLl_1_onRs_1_hazard && _zz_DispatchPlugin_logic_rsHazardChecker_1_onLl_1_onRs_1_hazard_1) && 1'b1) && (! toplevel_execute_ctrl1_down_BYPASSED_AT_2_lane1)),{((_zz_DispatchPlugin_logic_rsHazardChecker_1_onLl_1_onRs_1_hazard_2 && _zz_DispatchPlugin_logic_rsHazardChecker_1_onLl_1_onRs_1_hazard_3) && (! toplevel_execute_ctrl2_down_BYPASSED_AT_3_lane0)),((_zz_DispatchPlugin_logic_rsHazardChecker_1_onLl_1_onRs_1_hazard_4 && _zz_DispatchPlugin_logic_rsHazardChecker_1_onLl_1_onRs_1_hazard_5) && (! toplevel_execute_ctrl1_down_BYPASSED_AT_2_lane0))}}}));
  assign DispatchPlugin_logic_rsHazardChecker_1_onLl_2_onRs_0_hazard = (DispatchPlugin_logic_candidates_1_ctx_hm_RS1_ENABLE && 1'b0);
  assign DispatchPlugin_logic_rsHazardChecker_1_onLl_2_onRs_1_hazard = (DispatchPlugin_logic_candidates_1_ctx_hm_RS2_ENABLE && 1'b0);
  assign DispatchPlugin_logic_rsHazardChecker_1_onLl_3_onRs_0_hazard = (DispatchPlugin_logic_candidates_1_ctx_hm_RS1_ENABLE && 1'b0);
  assign DispatchPlugin_logic_rsHazardChecker_1_onLl_3_onRs_1_hazard = (DispatchPlugin_logic_candidates_1_ctx_hm_RS2_ENABLE && 1'b0);
  assign DispatchPlugin_logic_rsHazardChecker_2_onLl_0_onRs_0_hazard = (DispatchPlugin_logic_candidates_2_ctx_hm_RS1_ENABLE && (|{((((DispatchPlugin_logic_candidates_2_ctx_hm_DispatchPlugin_logic_hcs_0_onRs_0_ENABLES_0 && toplevel_execute_ctrl2_up_RD_ENABLE_lane1) && (toplevel_execute_ctrl2_up_RD_PHYS_lane1 == DispatchPlugin_logic_candidates_2_ctx_hm_RS1_PHYS)) && 1'b1) && (! toplevel_execute_ctrl2_down_BYPASSED_AT_3_lane1)),{(((_zz_DispatchPlugin_logic_rsHazardChecker_2_onLl_0_onRs_0_hazard && _zz_DispatchPlugin_logic_rsHazardChecker_2_onLl_0_onRs_0_hazard_1) && 1'b1) && (! toplevel_execute_ctrl1_down_BYPASSED_AT_2_lane1)),{((_zz_DispatchPlugin_logic_rsHazardChecker_2_onLl_0_onRs_0_hazard_2 && _zz_DispatchPlugin_logic_rsHazardChecker_2_onLl_0_onRs_0_hazard_3) && (! toplevel_execute_ctrl2_down_BYPASSED_AT_3_lane0)),((_zz_DispatchPlugin_logic_rsHazardChecker_2_onLl_0_onRs_0_hazard_4 && _zz_DispatchPlugin_logic_rsHazardChecker_2_onLl_0_onRs_0_hazard_5) && (! toplevel_execute_ctrl1_down_BYPASSED_AT_2_lane0))}}}));
  assign DispatchPlugin_logic_rsHazardChecker_2_onLl_0_onRs_1_hazard = (DispatchPlugin_logic_candidates_2_ctx_hm_RS2_ENABLE && (|{((((DispatchPlugin_logic_candidates_2_ctx_hm_DispatchPlugin_logic_hcs_0_onRs_1_ENABLES_0 && toplevel_execute_ctrl2_up_RD_ENABLE_lane1) && (toplevel_execute_ctrl2_up_RD_PHYS_lane1 == DispatchPlugin_logic_candidates_2_ctx_hm_RS2_PHYS)) && 1'b1) && (! toplevel_execute_ctrl2_down_BYPASSED_AT_3_lane1)),{(((_zz_DispatchPlugin_logic_rsHazardChecker_2_onLl_0_onRs_1_hazard && _zz_DispatchPlugin_logic_rsHazardChecker_2_onLl_0_onRs_1_hazard_1) && 1'b1) && (! toplevel_execute_ctrl1_down_BYPASSED_AT_2_lane1)),{((_zz_DispatchPlugin_logic_rsHazardChecker_2_onLl_0_onRs_1_hazard_2 && _zz_DispatchPlugin_logic_rsHazardChecker_2_onLl_0_onRs_1_hazard_3) && (! toplevel_execute_ctrl2_down_BYPASSED_AT_3_lane0)),((_zz_DispatchPlugin_logic_rsHazardChecker_2_onLl_0_onRs_1_hazard_4 && _zz_DispatchPlugin_logic_rsHazardChecker_2_onLl_0_onRs_1_hazard_5) && (! toplevel_execute_ctrl1_down_BYPASSED_AT_2_lane0))}}}));
  always @(*) begin
    DispatchPlugin_logic_candidates_2_rsHazards[0] = (|{DispatchPlugin_logic_rsHazardChecker_2_onLl_0_onRs_1_hazard,DispatchPlugin_logic_rsHazardChecker_2_onLl_0_onRs_0_hazard});
    DispatchPlugin_logic_candidates_2_rsHazards[1] = (|{DispatchPlugin_logic_rsHazardChecker_2_onLl_1_onRs_1_hazard,DispatchPlugin_logic_rsHazardChecker_2_onLl_1_onRs_0_hazard});
    DispatchPlugin_logic_candidates_2_rsHazards[2] = (|{DispatchPlugin_logic_rsHazardChecker_2_onLl_2_onRs_1_hazard,DispatchPlugin_logic_rsHazardChecker_2_onLl_2_onRs_0_hazard});
    DispatchPlugin_logic_candidates_2_rsHazards[3] = (|{DispatchPlugin_logic_rsHazardChecker_2_onLl_3_onRs_1_hazard,DispatchPlugin_logic_rsHazardChecker_2_onLl_3_onRs_0_hazard});
  end

  assign DispatchPlugin_logic_rsHazardChecker_2_onLl_1_onRs_0_hazard = (DispatchPlugin_logic_candidates_2_ctx_hm_RS1_ENABLE && (|{((((DispatchPlugin_logic_candidates_2_ctx_hm_DispatchPlugin_logic_hcs_1_onRs_0_ENABLES_0 && toplevel_execute_ctrl2_up_RD_ENABLE_lane1) && (toplevel_execute_ctrl2_up_RD_PHYS_lane1 == DispatchPlugin_logic_candidates_2_ctx_hm_RS1_PHYS)) && 1'b1) && (! toplevel_execute_ctrl2_down_BYPASSED_AT_3_lane1)),{(((_zz_DispatchPlugin_logic_rsHazardChecker_2_onLl_1_onRs_0_hazard && _zz_DispatchPlugin_logic_rsHazardChecker_2_onLl_1_onRs_0_hazard_1) && 1'b1) && (! toplevel_execute_ctrl1_down_BYPASSED_AT_2_lane1)),{((_zz_DispatchPlugin_logic_rsHazardChecker_2_onLl_1_onRs_0_hazard_2 && _zz_DispatchPlugin_logic_rsHazardChecker_2_onLl_1_onRs_0_hazard_3) && (! toplevel_execute_ctrl2_down_BYPASSED_AT_3_lane0)),((_zz_DispatchPlugin_logic_rsHazardChecker_2_onLl_1_onRs_0_hazard_4 && _zz_DispatchPlugin_logic_rsHazardChecker_2_onLl_1_onRs_0_hazard_5) && (! toplevel_execute_ctrl1_down_BYPASSED_AT_2_lane0))}}}));
  assign DispatchPlugin_logic_rsHazardChecker_2_onLl_1_onRs_1_hazard = (DispatchPlugin_logic_candidates_2_ctx_hm_RS2_ENABLE && (|{((((DispatchPlugin_logic_candidates_2_ctx_hm_DispatchPlugin_logic_hcs_1_onRs_1_ENABLES_0 && toplevel_execute_ctrl2_up_RD_ENABLE_lane1) && (toplevel_execute_ctrl2_up_RD_PHYS_lane1 == DispatchPlugin_logic_candidates_2_ctx_hm_RS2_PHYS)) && 1'b1) && (! toplevel_execute_ctrl2_down_BYPASSED_AT_3_lane1)),{(((_zz_DispatchPlugin_logic_rsHazardChecker_2_onLl_1_onRs_1_hazard && _zz_DispatchPlugin_logic_rsHazardChecker_2_onLl_1_onRs_1_hazard_1) && 1'b1) && (! toplevel_execute_ctrl1_down_BYPASSED_AT_2_lane1)),{((_zz_DispatchPlugin_logic_rsHazardChecker_2_onLl_1_onRs_1_hazard_2 && _zz_DispatchPlugin_logic_rsHazardChecker_2_onLl_1_onRs_1_hazard_3) && (! toplevel_execute_ctrl2_down_BYPASSED_AT_3_lane0)),((_zz_DispatchPlugin_logic_rsHazardChecker_2_onLl_1_onRs_1_hazard_4 && _zz_DispatchPlugin_logic_rsHazardChecker_2_onLl_1_onRs_1_hazard_5) && (! toplevel_execute_ctrl1_down_BYPASSED_AT_2_lane0))}}}));
  assign DispatchPlugin_logic_rsHazardChecker_2_onLl_2_onRs_0_hazard = (DispatchPlugin_logic_candidates_2_ctx_hm_RS1_ENABLE && 1'b0);
  assign DispatchPlugin_logic_rsHazardChecker_2_onLl_2_onRs_1_hazard = (DispatchPlugin_logic_candidates_2_ctx_hm_RS2_ENABLE && 1'b0);
  assign DispatchPlugin_logic_rsHazardChecker_2_onLl_3_onRs_0_hazard = (DispatchPlugin_logic_candidates_2_ctx_hm_RS1_ENABLE && 1'b0);
  assign DispatchPlugin_logic_rsHazardChecker_2_onLl_3_onRs_1_hazard = (DispatchPlugin_logic_candidates_2_ctx_hm_RS2_ENABLE && 1'b0);
  assign DispatchPlugin_logic_reservationChecker_0_onLl_0_hit = 1'b0;
  always @(*) begin
    DispatchPlugin_logic_candidates_0_reservationHazards[0] = DispatchPlugin_logic_reservationChecker_0_onLl_0_hit;
    DispatchPlugin_logic_candidates_0_reservationHazards[1] = DispatchPlugin_logic_reservationChecker_0_onLl_1_hit;
    DispatchPlugin_logic_candidates_0_reservationHazards[2] = DispatchPlugin_logic_reservationChecker_0_onLl_2_hit;
    DispatchPlugin_logic_candidates_0_reservationHazards[3] = DispatchPlugin_logic_reservationChecker_0_onLl_3_hit;
  end

  assign DispatchPlugin_logic_reservationChecker_0_onLl_1_hit = 1'b0;
  assign DispatchPlugin_logic_reservationChecker_0_onLl_2_hit = 1'b0;
  assign DispatchPlugin_logic_reservationChecker_0_onLl_3_hit = 1'b0;
  assign DispatchPlugin_logic_reservationChecker_1_onLl_0_hit = 1'b0;
  always @(*) begin
    DispatchPlugin_logic_candidates_1_reservationHazards[0] = DispatchPlugin_logic_reservationChecker_1_onLl_0_hit;
    DispatchPlugin_logic_candidates_1_reservationHazards[1] = DispatchPlugin_logic_reservationChecker_1_onLl_1_hit;
    DispatchPlugin_logic_candidates_1_reservationHazards[2] = DispatchPlugin_logic_reservationChecker_1_onLl_2_hit;
    DispatchPlugin_logic_candidates_1_reservationHazards[3] = DispatchPlugin_logic_reservationChecker_1_onLl_3_hit;
  end

  assign DispatchPlugin_logic_reservationChecker_1_onLl_1_hit = 1'b0;
  assign DispatchPlugin_logic_reservationChecker_1_onLl_2_hit = 1'b0;
  assign DispatchPlugin_logic_reservationChecker_1_onLl_3_hit = 1'b0;
  assign DispatchPlugin_logic_reservationChecker_2_onLl_0_hit = 1'b0;
  always @(*) begin
    DispatchPlugin_logic_candidates_2_reservationHazards[0] = DispatchPlugin_logic_reservationChecker_2_onLl_0_hit;
    DispatchPlugin_logic_candidates_2_reservationHazards[1] = DispatchPlugin_logic_reservationChecker_2_onLl_1_hit;
    DispatchPlugin_logic_candidates_2_reservationHazards[2] = DispatchPlugin_logic_reservationChecker_2_onLl_2_hit;
    DispatchPlugin_logic_candidates_2_reservationHazards[3] = DispatchPlugin_logic_reservationChecker_2_onLl_3_hit;
  end

  assign DispatchPlugin_logic_reservationChecker_2_onLl_1_hit = 1'b0;
  assign DispatchPlugin_logic_reservationChecker_2_onLl_2_hit = 1'b0;
  assign DispatchPlugin_logic_reservationChecker_2_onLl_3_hit = 1'b0;
  assign DispatchPlugin_logic_flushChecker_0_executeCheck_0_hits_0 = (|{(((DispatchPlugin_logic_candidates_0_ctx_hm_DONT_FLUSH_PRECISE_4 && toplevel_execute_ctrl1_up_LANE_SEL_lane0) && 1'b1) && toplevel_execute_ctrl1_down_MAY_FLUSH_PRECISE_4_lane0),(((DispatchPlugin_logic_candidates_0_ctx_hm_DONT_FLUSH_PRECISE_3 && toplevel_execute_ctrl1_up_LANE_SEL_lane0) && 1'b1) && toplevel_execute_ctrl1_down_MAY_FLUSH_PRECISE_3_lane0)});
  assign DispatchPlugin_logic_flushChecker_0_executeCheck_0_hits_1 = (|(((DispatchPlugin_logic_candidates_0_ctx_hm_DONT_FLUSH_PRECISE_3 && toplevel_execute_ctrl2_up_LANE_SEL_lane0) && 1'b1) && toplevel_execute_ctrl2_down_MAY_FLUSH_PRECISE_3_lane0));
  assign DispatchPlugin_logic_flushChecker_0_executeCheck_1_hits_0 = (|{(((DispatchPlugin_logic_candidates_0_ctx_hm_DONT_FLUSH_PRECISE_4 && toplevel_execute_ctrl1_up_LANE_SEL_lane1) && 1'b1) && toplevel_execute_ctrl1_down_MAY_FLUSH_PRECISE_4_lane1),(((DispatchPlugin_logic_candidates_0_ctx_hm_DONT_FLUSH_PRECISE_3 && toplevel_execute_ctrl1_up_LANE_SEL_lane1) && 1'b1) && toplevel_execute_ctrl1_down_MAY_FLUSH_PRECISE_3_lane1)});
  assign DispatchPlugin_logic_flushChecker_0_executeCheck_1_hits_1 = (|(((DispatchPlugin_logic_candidates_0_ctx_hm_DONT_FLUSH_PRECISE_3 && toplevel_execute_ctrl2_up_LANE_SEL_lane1) && 1'b1) && toplevel_execute_ctrl2_down_MAY_FLUSH_PRECISE_3_lane1));
  assign DispatchPlugin_logic_flushChecker_0_oldersHazard = 1'b0;
  assign DispatchPlugin_logic_candidates_0_flushHazards = ((|{DispatchPlugin_logic_flushChecker_0_executeCheck_1_hits_1,{DispatchPlugin_logic_flushChecker_0_executeCheck_1_hits_0,{DispatchPlugin_logic_flushChecker_0_executeCheck_0_hits_1,DispatchPlugin_logic_flushChecker_0_executeCheck_0_hits_0}}}) || (DispatchPlugin_logic_candidates_0_ctx_hm_DispatchPlugin_DONT_FLUSH_FROM_LANES && DispatchPlugin_logic_flushChecker_0_oldersHazard));
  assign DispatchPlugin_logic_flushChecker_1_executeCheck_0_hits_0 = (|{(((DispatchPlugin_logic_candidates_1_ctx_hm_DONT_FLUSH_PRECISE_4 && toplevel_execute_ctrl1_up_LANE_SEL_lane0) && 1'b1) && toplevel_execute_ctrl1_down_MAY_FLUSH_PRECISE_4_lane0),(((DispatchPlugin_logic_candidates_1_ctx_hm_DONT_FLUSH_PRECISE_3 && toplevel_execute_ctrl1_up_LANE_SEL_lane0) && 1'b1) && toplevel_execute_ctrl1_down_MAY_FLUSH_PRECISE_3_lane0)});
  assign DispatchPlugin_logic_flushChecker_1_executeCheck_0_hits_1 = (|(((DispatchPlugin_logic_candidates_1_ctx_hm_DONT_FLUSH_PRECISE_3 && toplevel_execute_ctrl2_up_LANE_SEL_lane0) && 1'b1) && toplevel_execute_ctrl2_down_MAY_FLUSH_PRECISE_3_lane0));
  assign DispatchPlugin_logic_flushChecker_1_executeCheck_1_hits_0 = (|{(((DispatchPlugin_logic_candidates_1_ctx_hm_DONT_FLUSH_PRECISE_4 && toplevel_execute_ctrl1_up_LANE_SEL_lane1) && 1'b1) && toplevel_execute_ctrl1_down_MAY_FLUSH_PRECISE_4_lane1),(((DispatchPlugin_logic_candidates_1_ctx_hm_DONT_FLUSH_PRECISE_3 && toplevel_execute_ctrl1_up_LANE_SEL_lane1) && 1'b1) && toplevel_execute_ctrl1_down_MAY_FLUSH_PRECISE_3_lane1)});
  assign DispatchPlugin_logic_flushChecker_1_executeCheck_1_hits_1 = (|(((DispatchPlugin_logic_candidates_1_ctx_hm_DONT_FLUSH_PRECISE_3 && toplevel_execute_ctrl2_up_LANE_SEL_lane1) && 1'b1) && toplevel_execute_ctrl2_down_MAY_FLUSH_PRECISE_3_lane1));
  assign DispatchPlugin_logic_flushChecker_1_oldersHazard = (|(DispatchPlugin_logic_candidates_0_ctx_valid && DispatchPlugin_logic_candidates_0_ctx_hm_DispatchPlugin_MAY_FLUSH));
  assign DispatchPlugin_logic_candidates_1_flushHazards = ((|{DispatchPlugin_logic_flushChecker_1_executeCheck_1_hits_1,{DispatchPlugin_logic_flushChecker_1_executeCheck_1_hits_0,{DispatchPlugin_logic_flushChecker_1_executeCheck_0_hits_1,DispatchPlugin_logic_flushChecker_1_executeCheck_0_hits_0}}}) || (DispatchPlugin_logic_candidates_1_ctx_hm_DispatchPlugin_DONT_FLUSH_FROM_LANES && DispatchPlugin_logic_flushChecker_1_oldersHazard));
  assign DispatchPlugin_logic_flushChecker_2_executeCheck_0_hits_0 = (|{(((DispatchPlugin_logic_candidates_2_ctx_hm_DONT_FLUSH_PRECISE_4 && toplevel_execute_ctrl1_up_LANE_SEL_lane0) && 1'b1) && toplevel_execute_ctrl1_down_MAY_FLUSH_PRECISE_4_lane0),(((DispatchPlugin_logic_candidates_2_ctx_hm_DONT_FLUSH_PRECISE_3 && toplevel_execute_ctrl1_up_LANE_SEL_lane0) && 1'b1) && toplevel_execute_ctrl1_down_MAY_FLUSH_PRECISE_3_lane0)});
  assign DispatchPlugin_logic_flushChecker_2_executeCheck_0_hits_1 = (|(((DispatchPlugin_logic_candidates_2_ctx_hm_DONT_FLUSH_PRECISE_3 && toplevel_execute_ctrl2_up_LANE_SEL_lane0) && 1'b1) && toplevel_execute_ctrl2_down_MAY_FLUSH_PRECISE_3_lane0));
  assign DispatchPlugin_logic_flushChecker_2_executeCheck_1_hits_0 = (|{(((DispatchPlugin_logic_candidates_2_ctx_hm_DONT_FLUSH_PRECISE_4 && toplevel_execute_ctrl1_up_LANE_SEL_lane1) && 1'b1) && toplevel_execute_ctrl1_down_MAY_FLUSH_PRECISE_4_lane1),(((DispatchPlugin_logic_candidates_2_ctx_hm_DONT_FLUSH_PRECISE_3 && toplevel_execute_ctrl1_up_LANE_SEL_lane1) && 1'b1) && toplevel_execute_ctrl1_down_MAY_FLUSH_PRECISE_3_lane1)});
  assign DispatchPlugin_logic_flushChecker_2_executeCheck_1_hits_1 = (|(((DispatchPlugin_logic_candidates_2_ctx_hm_DONT_FLUSH_PRECISE_3 && toplevel_execute_ctrl2_up_LANE_SEL_lane1) && 1'b1) && toplevel_execute_ctrl2_down_MAY_FLUSH_PRECISE_3_lane1));
  assign DispatchPlugin_logic_flushChecker_2_oldersHazard = (|{(DispatchPlugin_logic_candidates_1_ctx_valid && DispatchPlugin_logic_candidates_1_ctx_hm_DispatchPlugin_MAY_FLUSH),(DispatchPlugin_logic_candidates_0_ctx_valid && DispatchPlugin_logic_candidates_0_ctx_hm_DispatchPlugin_MAY_FLUSH)});
  assign DispatchPlugin_logic_candidates_2_flushHazards = ((|{DispatchPlugin_logic_flushChecker_2_executeCheck_1_hits_1,{DispatchPlugin_logic_flushChecker_2_executeCheck_1_hits_0,{DispatchPlugin_logic_flushChecker_2_executeCheck_0_hits_1,DispatchPlugin_logic_flushChecker_2_executeCheck_0_hits_0}}}) || (DispatchPlugin_logic_candidates_2_ctx_hm_DispatchPlugin_DONT_FLUSH_FROM_LANES && DispatchPlugin_logic_flushChecker_2_oldersHazard));
  assign DispatchPlugin_logic_fenceChecker_olderInflights = (|{execute_lane1_api_hartsInflight[0],execute_lane0_api_hartsInflight[0]});
  assign DispatchPlugin_logic_candidates_0_fenceOlderHazards = (DispatchPlugin_logic_candidates_0_ctx_hm_DispatchPlugin_FENCE_OLDER && (DispatchPlugin_logic_fenceChecker_olderInflights[0] || 1'b0));
  assign DispatchPlugin_logic_candidates_1_fenceOlderHazards = (DispatchPlugin_logic_candidates_1_ctx_hm_DispatchPlugin_FENCE_OLDER && (DispatchPlugin_logic_fenceChecker_olderInflights[0] || (|(DispatchPlugin_logic_candidates_0_ctx_valid && 1'b1))));
  assign DispatchPlugin_logic_candidates_2_fenceOlderHazards = (DispatchPlugin_logic_candidates_2_ctx_hm_DispatchPlugin_FENCE_OLDER && (DispatchPlugin_logic_fenceChecker_olderInflights[0] || (|{(DispatchPlugin_logic_candidates_1_ctx_valid && 1'b1),(DispatchPlugin_logic_candidates_0_ctx_valid && 1'b1)})));
  always @(*) begin
    toplevel_decode_ctrls_1_down_ready = 1'b1;
    if(when_DispatchPlugin_l358) begin
      toplevel_decode_ctrls_1_down_ready = 1'b0;
    end
    if(when_DispatchPlugin_l358_1) begin
      toplevel_decode_ctrls_1_down_ready = 1'b0;
    end
    if(DispatchPlugin_logic_slotsFeeds_doIt) begin
      toplevel_decode_ctrls_1_down_ready = 1'b1;
    end
  end

  assign DispatchPlugin_logic_feeds_0_sending = DispatchPlugin_logic_candidates_1_fire;
  assign DispatchPlugin_logic_candidates_1_cancel = toplevel_decode_ctrls_1_lane0_upIsCancel;
  assign DispatchPlugin_logic_candidates_1_ctx_valid = ((toplevel_decode_ctrls_1_up_isValid && toplevel_decode_ctrls_1_up_LANE_SEL_0) && (! DispatchPlugin_logic_feeds_0_sent));
  always @(*) begin
    DispatchPlugin_logic_candidates_1_ctx_laneLayerHits = {toplevel_decode_ctrls_1_down_DispatchPlugin_logic_LANES_LAYER_HIT_3_0,{toplevel_decode_ctrls_1_down_DispatchPlugin_logic_LANES_LAYER_HIT_2_0,{toplevel_decode_ctrls_1_down_DispatchPlugin_logic_LANES_LAYER_HIT_1_0,toplevel_decode_ctrls_1_down_DispatchPlugin_logic_LANES_LAYER_HIT_0_0}}};
    if(toplevel_decode_ctrls_1_down_TRAP_0) begin
      DispatchPlugin_logic_candidates_1_ctx_laneLayerHits = 4'b0010;
    end
  end

  assign DispatchPlugin_logic_candidates_1_ctx_uop = toplevel_decode_ctrls_1_down_Decode_UOP_0;
  assign DispatchPlugin_logic_candidates_1_ctx_hm_Prediction_ALIGNED_JUMPED = toplevel_decode_ctrls_1_down_Prediction_ALIGNED_JUMPED_0;
  assign DispatchPlugin_logic_candidates_1_ctx_hm_Prediction_ALIGNED_JUMPED_PC = toplevel_decode_ctrls_1_down_Prediction_ALIGNED_JUMPED_PC_0;
  assign DispatchPlugin_logic_candidates_1_ctx_hm_Prediction_ALIGNED_SLICES_TAKEN = toplevel_decode_ctrls_1_down_Prediction_ALIGNED_SLICES_TAKEN_0;
  assign DispatchPlugin_logic_candidates_1_ctx_hm_Prediction_ALIGNED_SLICES_BRANCH = toplevel_decode_ctrls_1_down_Prediction_ALIGNED_SLICES_BRANCH_0;
  assign DispatchPlugin_logic_candidates_1_ctx_hm_GSharePlugin_GSHARE_COUNTER_0 = toplevel_decode_ctrls_1_down_GSharePlugin_GSHARE_COUNTER_0_0;
  assign DispatchPlugin_logic_candidates_1_ctx_hm_GSharePlugin_GSHARE_COUNTER_1 = toplevel_decode_ctrls_1_down_GSharePlugin_GSHARE_COUNTER_0_1;
  assign DispatchPlugin_logic_candidates_1_ctx_hm_GSharePlugin_GSHARE_COUNTER_2 = toplevel_decode_ctrls_1_down_GSharePlugin_GSHARE_COUNTER_0_2;
  assign DispatchPlugin_logic_candidates_1_ctx_hm_GSharePlugin_GSHARE_COUNTER_3 = toplevel_decode_ctrls_1_down_GSharePlugin_GSHARE_COUNTER_0_3;
  assign DispatchPlugin_logic_candidates_1_ctx_hm_Prediction_BRANCH_HISTORY = toplevel_decode_ctrls_1_down_Prediction_BRANCH_HISTORY_0;
  assign DispatchPlugin_logic_candidates_1_ctx_hm_DispatchPlugin_FENCE_OLDER = toplevel_decode_ctrls_1_down_DispatchPlugin_FENCE_OLDER_0;
  assign DispatchPlugin_logic_candidates_1_ctx_hm_DispatchPlugin_MAY_FLUSH = toplevel_decode_ctrls_1_down_DispatchPlugin_MAY_FLUSH_0;
  assign DispatchPlugin_logic_candidates_1_ctx_hm_DispatchPlugin_DONT_FLUSH = toplevel_decode_ctrls_1_down_DispatchPlugin_DONT_FLUSH_0;
  assign DispatchPlugin_logic_candidates_1_ctx_hm_DispatchPlugin_DONT_FLUSH_FROM_LANES = toplevel_decode_ctrls_1_down_DispatchPlugin_DONT_FLUSH_FROM_LANES_0;
  assign DispatchPlugin_logic_candidates_1_ctx_hm_Decode_INSTRUCTION_SLICE_COUNT = toplevel_decode_ctrls_1_down_Decode_INSTRUCTION_SLICE_COUNT_0;
  assign DispatchPlugin_logic_candidates_1_ctx_hm_DONT_FLUSH_PRECISE_3 = toplevel_decode_ctrls_1_down_DONT_FLUSH_PRECISE_3_0;
  assign DispatchPlugin_logic_candidates_1_ctx_hm_DONT_FLUSH_PRECISE_4 = toplevel_decode_ctrls_1_down_DONT_FLUSH_PRECISE_4_0;
  assign DispatchPlugin_logic_candidates_1_ctx_hm_PC = toplevel_decode_ctrls_1_down_PC_0;
  assign DispatchPlugin_logic_candidates_1_ctx_hm_TRAP = toplevel_decode_ctrls_1_down_TRAP_0;
  assign DispatchPlugin_logic_candidates_1_ctx_hm_Decode_UOP_ID = toplevel_decode_ctrls_1_down_Decode_UOP_ID_0;
  assign DispatchPlugin_logic_candidates_1_ctx_hm_RS1_ENABLE = toplevel_decode_ctrls_1_down_RS1_ENABLE_0;
  assign DispatchPlugin_logic_candidates_1_ctx_hm_RS1_PHYS = toplevel_decode_ctrls_1_down_RS1_PHYS_0;
  assign DispatchPlugin_logic_candidates_1_ctx_hm_RS2_ENABLE = toplevel_decode_ctrls_1_down_RS2_ENABLE_0;
  assign DispatchPlugin_logic_candidates_1_ctx_hm_RS2_PHYS = toplevel_decode_ctrls_1_down_RS2_PHYS_0;
  assign DispatchPlugin_logic_candidates_1_ctx_hm_RD_ENABLE = toplevel_decode_ctrls_1_down_RD_ENABLE_0;
  assign DispatchPlugin_logic_candidates_1_ctx_hm_RD_PHYS = toplevel_decode_ctrls_1_down_RD_PHYS_0;
  assign DispatchPlugin_logic_candidates_1_ctx_hm_DispatchPlugin_logic_hcs_0_onRs_0_ENABLES_0 = toplevel_decode_ctrls_1_down_DispatchPlugin_logic_hcs_0_onRs_0_ENABLES_0_0;
  assign DispatchPlugin_logic_candidates_1_ctx_hm_DispatchPlugin_logic_hcs_0_onRs_1_ENABLES_0 = toplevel_decode_ctrls_1_down_DispatchPlugin_logic_hcs_0_onRs_1_ENABLES_0_0;
  assign DispatchPlugin_logic_candidates_1_ctx_hm_DispatchPlugin_logic_hcs_1_onRs_0_ENABLES_0 = toplevel_decode_ctrls_1_down_DispatchPlugin_logic_hcs_1_onRs_0_ENABLES_0_0;
  assign DispatchPlugin_logic_candidates_1_ctx_hm_DispatchPlugin_logic_hcs_1_onRs_1_ENABLES_0 = toplevel_decode_ctrls_1_down_DispatchPlugin_logic_hcs_1_onRs_1_ENABLES_0_0;
  assign DispatchPlugin_logic_candidates_1_ctx_hm_DispatchPlugin_logic_hcs_1_onRs_1_ENABLES_1 = toplevel_decode_ctrls_1_down_DispatchPlugin_logic_hcs_1_onRs_1_ENABLES_1_0;
  assign DispatchPlugin_logic_candidates_1_ctx_hm_DispatchPlugin_logic_hcs_2_onRs_0_ENABLES_0 = toplevel_decode_ctrls_1_down_DispatchPlugin_logic_hcs_2_onRs_0_ENABLES_0_0;
  assign DispatchPlugin_logic_candidates_1_ctx_hm_DispatchPlugin_logic_hcs_2_onRs_1_ENABLES_0 = toplevel_decode_ctrls_1_down_DispatchPlugin_logic_hcs_2_onRs_1_ENABLES_0_0;
  assign DispatchPlugin_logic_candidates_1_ctx_hm_DispatchPlugin_logic_hcs_3_onRs_0_ENABLES_0 = toplevel_decode_ctrls_1_down_DispatchPlugin_logic_hcs_3_onRs_0_ENABLES_0_0;
  assign DispatchPlugin_logic_candidates_1_ctx_hm_DispatchPlugin_logic_hcs_3_onRs_1_ENABLES_0 = toplevel_decode_ctrls_1_down_DispatchPlugin_logic_hcs_3_onRs_1_ENABLES_0_0;
  assign when_DispatchPlugin_l358 = ((toplevel_decode_ctrls_1_up_LANE_SEL_0 && (! DispatchPlugin_logic_feeds_0_sent)) && (! DispatchPlugin_logic_candidates_1_fire));
  assign DispatchPlugin_logic_feeds_1_sending = DispatchPlugin_logic_candidates_2_fire;
  assign DispatchPlugin_logic_candidates_2_cancel = toplevel_decode_ctrls_1_lane1_upIsCancel;
  assign DispatchPlugin_logic_candidates_2_ctx_valid = ((toplevel_decode_ctrls_1_up_isValid && toplevel_decode_ctrls_1_up_LANE_SEL_1) && (! DispatchPlugin_logic_feeds_1_sent));
  always @(*) begin
    DispatchPlugin_logic_candidates_2_ctx_laneLayerHits = {toplevel_decode_ctrls_1_down_DispatchPlugin_logic_LANES_LAYER_HIT_3_1,{toplevel_decode_ctrls_1_down_DispatchPlugin_logic_LANES_LAYER_HIT_2_1,{toplevel_decode_ctrls_1_down_DispatchPlugin_logic_LANES_LAYER_HIT_1_1,toplevel_decode_ctrls_1_down_DispatchPlugin_logic_LANES_LAYER_HIT_0_1}}};
    if(toplevel_decode_ctrls_1_down_TRAP_1) begin
      DispatchPlugin_logic_candidates_2_ctx_laneLayerHits = 4'b0010;
    end
  end

  assign DispatchPlugin_logic_candidates_2_ctx_uop = toplevel_decode_ctrls_1_down_Decode_UOP_1;
  assign DispatchPlugin_logic_candidates_2_ctx_hm_Prediction_ALIGNED_JUMPED = toplevel_decode_ctrls_1_down_Prediction_ALIGNED_JUMPED_1;
  assign DispatchPlugin_logic_candidates_2_ctx_hm_Prediction_ALIGNED_JUMPED_PC = toplevel_decode_ctrls_1_down_Prediction_ALIGNED_JUMPED_PC_1;
  assign DispatchPlugin_logic_candidates_2_ctx_hm_Prediction_ALIGNED_SLICES_TAKEN = toplevel_decode_ctrls_1_down_Prediction_ALIGNED_SLICES_TAKEN_1;
  assign DispatchPlugin_logic_candidates_2_ctx_hm_Prediction_ALIGNED_SLICES_BRANCH = toplevel_decode_ctrls_1_down_Prediction_ALIGNED_SLICES_BRANCH_1;
  assign DispatchPlugin_logic_candidates_2_ctx_hm_GSharePlugin_GSHARE_COUNTER_0 = toplevel_decode_ctrls_1_down_GSharePlugin_GSHARE_COUNTER_1_0;
  assign DispatchPlugin_logic_candidates_2_ctx_hm_GSharePlugin_GSHARE_COUNTER_1 = toplevel_decode_ctrls_1_down_GSharePlugin_GSHARE_COUNTER_1_1;
  assign DispatchPlugin_logic_candidates_2_ctx_hm_GSharePlugin_GSHARE_COUNTER_2 = toplevel_decode_ctrls_1_down_GSharePlugin_GSHARE_COUNTER_1_2;
  assign DispatchPlugin_logic_candidates_2_ctx_hm_GSharePlugin_GSHARE_COUNTER_3 = toplevel_decode_ctrls_1_down_GSharePlugin_GSHARE_COUNTER_1_3;
  assign DispatchPlugin_logic_candidates_2_ctx_hm_Prediction_BRANCH_HISTORY = toplevel_decode_ctrls_1_down_Prediction_BRANCH_HISTORY_1;
  assign DispatchPlugin_logic_candidates_2_ctx_hm_DispatchPlugin_FENCE_OLDER = toplevel_decode_ctrls_1_down_DispatchPlugin_FENCE_OLDER_1;
  assign DispatchPlugin_logic_candidates_2_ctx_hm_DispatchPlugin_MAY_FLUSH = toplevel_decode_ctrls_1_down_DispatchPlugin_MAY_FLUSH_1;
  assign DispatchPlugin_logic_candidates_2_ctx_hm_DispatchPlugin_DONT_FLUSH = toplevel_decode_ctrls_1_down_DispatchPlugin_DONT_FLUSH_1;
  assign DispatchPlugin_logic_candidates_2_ctx_hm_DispatchPlugin_DONT_FLUSH_FROM_LANES = toplevel_decode_ctrls_1_down_DispatchPlugin_DONT_FLUSH_FROM_LANES_1;
  assign DispatchPlugin_logic_candidates_2_ctx_hm_Decode_INSTRUCTION_SLICE_COUNT = toplevel_decode_ctrls_1_down_Decode_INSTRUCTION_SLICE_COUNT_1;
  assign DispatchPlugin_logic_candidates_2_ctx_hm_DONT_FLUSH_PRECISE_3 = toplevel_decode_ctrls_1_down_DONT_FLUSH_PRECISE_3_1;
  assign DispatchPlugin_logic_candidates_2_ctx_hm_DONT_FLUSH_PRECISE_4 = toplevel_decode_ctrls_1_down_DONT_FLUSH_PRECISE_4_1;
  assign DispatchPlugin_logic_candidates_2_ctx_hm_PC = toplevel_decode_ctrls_1_down_PC_1;
  assign DispatchPlugin_logic_candidates_2_ctx_hm_TRAP = toplevel_decode_ctrls_1_down_TRAP_1;
  assign DispatchPlugin_logic_candidates_2_ctx_hm_Decode_UOP_ID = toplevel_decode_ctrls_1_down_Decode_UOP_ID_1;
  assign DispatchPlugin_logic_candidates_2_ctx_hm_RS1_ENABLE = toplevel_decode_ctrls_1_down_RS1_ENABLE_1;
  assign DispatchPlugin_logic_candidates_2_ctx_hm_RS1_PHYS = toplevel_decode_ctrls_1_down_RS1_PHYS_1;
  assign DispatchPlugin_logic_candidates_2_ctx_hm_RS2_ENABLE = toplevel_decode_ctrls_1_down_RS2_ENABLE_1;
  assign DispatchPlugin_logic_candidates_2_ctx_hm_RS2_PHYS = toplevel_decode_ctrls_1_down_RS2_PHYS_1;
  assign DispatchPlugin_logic_candidates_2_ctx_hm_RD_ENABLE = toplevel_decode_ctrls_1_down_RD_ENABLE_1;
  assign DispatchPlugin_logic_candidates_2_ctx_hm_RD_PHYS = toplevel_decode_ctrls_1_down_RD_PHYS_1;
  assign DispatchPlugin_logic_candidates_2_ctx_hm_DispatchPlugin_logic_hcs_0_onRs_0_ENABLES_0 = toplevel_decode_ctrls_1_down_DispatchPlugin_logic_hcs_0_onRs_0_ENABLES_0_1;
  assign DispatchPlugin_logic_candidates_2_ctx_hm_DispatchPlugin_logic_hcs_0_onRs_1_ENABLES_0 = toplevel_decode_ctrls_1_down_DispatchPlugin_logic_hcs_0_onRs_1_ENABLES_0_1;
  assign DispatchPlugin_logic_candidates_2_ctx_hm_DispatchPlugin_logic_hcs_1_onRs_0_ENABLES_0 = toplevel_decode_ctrls_1_down_DispatchPlugin_logic_hcs_1_onRs_0_ENABLES_0_1;
  assign DispatchPlugin_logic_candidates_2_ctx_hm_DispatchPlugin_logic_hcs_1_onRs_1_ENABLES_0 = toplevel_decode_ctrls_1_down_DispatchPlugin_logic_hcs_1_onRs_1_ENABLES_0_1;
  assign DispatchPlugin_logic_candidates_2_ctx_hm_DispatchPlugin_logic_hcs_1_onRs_1_ENABLES_1 = toplevel_decode_ctrls_1_down_DispatchPlugin_logic_hcs_1_onRs_1_ENABLES_1_1;
  assign DispatchPlugin_logic_candidates_2_ctx_hm_DispatchPlugin_logic_hcs_2_onRs_0_ENABLES_0 = toplevel_decode_ctrls_1_down_DispatchPlugin_logic_hcs_2_onRs_0_ENABLES_0_1;
  assign DispatchPlugin_logic_candidates_2_ctx_hm_DispatchPlugin_logic_hcs_2_onRs_1_ENABLES_0 = toplevel_decode_ctrls_1_down_DispatchPlugin_logic_hcs_2_onRs_1_ENABLES_0_1;
  assign DispatchPlugin_logic_candidates_2_ctx_hm_DispatchPlugin_logic_hcs_3_onRs_0_ENABLES_0 = toplevel_decode_ctrls_1_down_DispatchPlugin_logic_hcs_3_onRs_0_ENABLES_0_1;
  assign DispatchPlugin_logic_candidates_2_ctx_hm_DispatchPlugin_logic_hcs_3_onRs_1_ENABLES_0 = toplevel_decode_ctrls_1_down_DispatchPlugin_logic_hcs_3_onRs_1_ENABLES_0_1;
  assign when_DispatchPlugin_l358_1 = ((toplevel_decode_ctrls_1_up_LANE_SEL_1 && (! DispatchPlugin_logic_feeds_1_sent)) && (! DispatchPlugin_logic_candidates_2_fire));
  assign DispatchPlugin_logic_candidates_0_ctx_valid = DispatchPlugin_logic_slots_0_ctx_valid;
  assign DispatchPlugin_logic_candidates_0_ctx_laneLayerHits = DispatchPlugin_logic_slots_0_ctx_laneLayerHits;
  assign DispatchPlugin_logic_candidates_0_ctx_uop = DispatchPlugin_logic_slots_0_ctx_uop;
  assign DispatchPlugin_logic_candidates_0_ctx_hm_Prediction_ALIGNED_JUMPED = DispatchPlugin_logic_slots_0_ctx_hm_Prediction_ALIGNED_JUMPED;
  assign DispatchPlugin_logic_candidates_0_ctx_hm_Prediction_ALIGNED_JUMPED_PC = DispatchPlugin_logic_slots_0_ctx_hm_Prediction_ALIGNED_JUMPED_PC;
  assign DispatchPlugin_logic_candidates_0_ctx_hm_Prediction_ALIGNED_SLICES_TAKEN = DispatchPlugin_logic_slots_0_ctx_hm_Prediction_ALIGNED_SLICES_TAKEN;
  assign DispatchPlugin_logic_candidates_0_ctx_hm_Prediction_ALIGNED_SLICES_BRANCH = DispatchPlugin_logic_slots_0_ctx_hm_Prediction_ALIGNED_SLICES_BRANCH;
  assign DispatchPlugin_logic_candidates_0_ctx_hm_GSharePlugin_GSHARE_COUNTER_0 = DispatchPlugin_logic_slots_0_ctx_hm_GSharePlugin_GSHARE_COUNTER_0;
  assign DispatchPlugin_logic_candidates_0_ctx_hm_GSharePlugin_GSHARE_COUNTER_1 = DispatchPlugin_logic_slots_0_ctx_hm_GSharePlugin_GSHARE_COUNTER_1;
  assign DispatchPlugin_logic_candidates_0_ctx_hm_GSharePlugin_GSHARE_COUNTER_2 = DispatchPlugin_logic_slots_0_ctx_hm_GSharePlugin_GSHARE_COUNTER_2;
  assign DispatchPlugin_logic_candidates_0_ctx_hm_GSharePlugin_GSHARE_COUNTER_3 = DispatchPlugin_logic_slots_0_ctx_hm_GSharePlugin_GSHARE_COUNTER_3;
  assign DispatchPlugin_logic_candidates_0_ctx_hm_Prediction_BRANCH_HISTORY = DispatchPlugin_logic_slots_0_ctx_hm_Prediction_BRANCH_HISTORY;
  assign DispatchPlugin_logic_candidates_0_ctx_hm_DispatchPlugin_FENCE_OLDER = DispatchPlugin_logic_slots_0_ctx_hm_DispatchPlugin_FENCE_OLDER;
  assign DispatchPlugin_logic_candidates_0_ctx_hm_DispatchPlugin_MAY_FLUSH = DispatchPlugin_logic_slots_0_ctx_hm_DispatchPlugin_MAY_FLUSH;
  assign DispatchPlugin_logic_candidates_0_ctx_hm_DispatchPlugin_DONT_FLUSH = DispatchPlugin_logic_slots_0_ctx_hm_DispatchPlugin_DONT_FLUSH;
  assign DispatchPlugin_logic_candidates_0_ctx_hm_DispatchPlugin_DONT_FLUSH_FROM_LANES = DispatchPlugin_logic_slots_0_ctx_hm_DispatchPlugin_DONT_FLUSH_FROM_LANES;
  assign DispatchPlugin_logic_candidates_0_ctx_hm_Decode_INSTRUCTION_SLICE_COUNT = DispatchPlugin_logic_slots_0_ctx_hm_Decode_INSTRUCTION_SLICE_COUNT;
  assign DispatchPlugin_logic_candidates_0_ctx_hm_DONT_FLUSH_PRECISE_3 = DispatchPlugin_logic_slots_0_ctx_hm_DONT_FLUSH_PRECISE_3;
  assign DispatchPlugin_logic_candidates_0_ctx_hm_DONT_FLUSH_PRECISE_4 = DispatchPlugin_logic_slots_0_ctx_hm_DONT_FLUSH_PRECISE_4;
  assign DispatchPlugin_logic_candidates_0_ctx_hm_PC = DispatchPlugin_logic_slots_0_ctx_hm_PC;
  assign DispatchPlugin_logic_candidates_0_ctx_hm_TRAP = DispatchPlugin_logic_slots_0_ctx_hm_TRAP;
  assign DispatchPlugin_logic_candidates_0_ctx_hm_Decode_UOP_ID = DispatchPlugin_logic_slots_0_ctx_hm_Decode_UOP_ID;
  assign DispatchPlugin_logic_candidates_0_ctx_hm_RS1_ENABLE = DispatchPlugin_logic_slots_0_ctx_hm_RS1_ENABLE;
  assign DispatchPlugin_logic_candidates_0_ctx_hm_RS1_PHYS = DispatchPlugin_logic_slots_0_ctx_hm_RS1_PHYS;
  assign DispatchPlugin_logic_candidates_0_ctx_hm_RS2_ENABLE = DispatchPlugin_logic_slots_0_ctx_hm_RS2_ENABLE;
  assign DispatchPlugin_logic_candidates_0_ctx_hm_RS2_PHYS = DispatchPlugin_logic_slots_0_ctx_hm_RS2_PHYS;
  assign DispatchPlugin_logic_candidates_0_ctx_hm_RD_ENABLE = DispatchPlugin_logic_slots_0_ctx_hm_RD_ENABLE;
  assign DispatchPlugin_logic_candidates_0_ctx_hm_RD_PHYS = DispatchPlugin_logic_slots_0_ctx_hm_RD_PHYS;
  assign DispatchPlugin_logic_candidates_0_ctx_hm_DispatchPlugin_logic_hcs_0_onRs_0_ENABLES_0 = DispatchPlugin_logic_slots_0_ctx_hm_DispatchPlugin_logic_hcs_0_onRs_0_ENABLES_0;
  assign DispatchPlugin_logic_candidates_0_ctx_hm_DispatchPlugin_logic_hcs_0_onRs_1_ENABLES_0 = DispatchPlugin_logic_slots_0_ctx_hm_DispatchPlugin_logic_hcs_0_onRs_1_ENABLES_0;
  assign DispatchPlugin_logic_candidates_0_ctx_hm_DispatchPlugin_logic_hcs_1_onRs_0_ENABLES_0 = DispatchPlugin_logic_slots_0_ctx_hm_DispatchPlugin_logic_hcs_1_onRs_0_ENABLES_0;
  assign DispatchPlugin_logic_candidates_0_ctx_hm_DispatchPlugin_logic_hcs_1_onRs_1_ENABLES_0 = DispatchPlugin_logic_slots_0_ctx_hm_DispatchPlugin_logic_hcs_1_onRs_1_ENABLES_0;
  assign DispatchPlugin_logic_candidates_0_ctx_hm_DispatchPlugin_logic_hcs_1_onRs_1_ENABLES_1 = DispatchPlugin_logic_slots_0_ctx_hm_DispatchPlugin_logic_hcs_1_onRs_1_ENABLES_1;
  assign DispatchPlugin_logic_candidates_0_ctx_hm_DispatchPlugin_logic_hcs_2_onRs_0_ENABLES_0 = DispatchPlugin_logic_slots_0_ctx_hm_DispatchPlugin_logic_hcs_2_onRs_0_ENABLES_0;
  assign DispatchPlugin_logic_candidates_0_ctx_hm_DispatchPlugin_logic_hcs_2_onRs_1_ENABLES_0 = DispatchPlugin_logic_slots_0_ctx_hm_DispatchPlugin_logic_hcs_2_onRs_1_ENABLES_0;
  assign DispatchPlugin_logic_candidates_0_ctx_hm_DispatchPlugin_logic_hcs_3_onRs_0_ENABLES_0 = DispatchPlugin_logic_slots_0_ctx_hm_DispatchPlugin_logic_hcs_3_onRs_0_ENABLES_0;
  assign DispatchPlugin_logic_candidates_0_ctx_hm_DispatchPlugin_logic_hcs_3_onRs_1_ENABLES_0 = DispatchPlugin_logic_slots_0_ctx_hm_DispatchPlugin_logic_hcs_3_onRs_1_ENABLES_0;
  assign when_DispatchPlugin_l368 = (DispatchPlugin_logic_candidates_0_fire || DispatchPlugin_logic_candidates_0_cancel);
  assign _zz_toplevel_decode_ctrls_1_down_DispatchPlugin_logic_LANES_LAYER_HIT_3_0_1 = ((toplevel_decode_ctrls_1_down_Decode_INSTRUCTION_0 & 32'h02000050) == 32'h00000010);
  assign _zz_toplevel_decode_ctrls_1_down_DispatchPlugin_logic_LANES_LAYER_HIT_3_0_2 = ((toplevel_decode_ctrls_1_down_Decode_INSTRUCTION_0 & 32'h00000030) == 32'h00000010);
  assign toplevel_decode_ctrls_1_down_DispatchPlugin_logic_LANES_LAYER_HIT_0_0 = _zz_toplevel_decode_ctrls_1_down_DispatchPlugin_logic_LANES_LAYER_HIT_0_0_2[0];
  assign _zz_toplevel_decode_ctrls_1_down_DispatchPlugin_logic_hcs_3_onRs_1_ENABLES_0_0 = ((toplevel_decode_ctrls_1_down_Decode_INSTRUCTION_0 & 32'h0) == 32'h0);
  assign toplevel_decode_ctrls_1_down_DispatchPlugin_logic_LANES_LAYER_HIT_1_0 = _zz_toplevel_decode_ctrls_1_down_DispatchPlugin_logic_LANES_LAYER_HIT_1_0[0];
  assign _zz_toplevel_decode_ctrls_1_down_DispatchPlugin_logic_LANES_LAYER_HIT_3_0_3 = ((toplevel_decode_ctrls_1_down_Decode_INSTRUCTION_0 & 32'h00000054) == 32'h00000040);
  assign _zz_toplevel_decode_ctrls_1_down_DispatchPlugin_logic_LANES_LAYER_HIT_3_0_4 = ((toplevel_decode_ctrls_1_down_Decode_INSTRUCTION_0 & 32'h0000004c) == 32'h00000004);
  assign toplevel_decode_ctrls_1_down_DispatchPlugin_logic_LANES_LAYER_HIT_2_0 = _zz_toplevel_decode_ctrls_1_down_DispatchPlugin_logic_LANES_LAYER_HIT_2_0[0];
  assign toplevel_decode_ctrls_1_down_DispatchPlugin_logic_LANES_LAYER_HIT_3_0 = _zz_toplevel_decode_ctrls_1_down_DispatchPlugin_logic_LANES_LAYER_HIT_3_0_5[0];
  assign _zz_toplevel_decode_ctrls_1_down_DispatchPlugin_logic_hcs_1_onRs_1_ENABLES_0_0 = ((toplevel_decode_ctrls_1_down_Decode_INSTRUCTION_0 & 32'h00000040) == 32'h00000040);
  assign toplevel_decode_ctrls_1_down_DispatchPlugin_MAY_FLUSH_0 = _zz_toplevel_decode_ctrls_1_down_DispatchPlugin_MAY_FLUSH_0_1[0];
  assign _zz_toplevel_decode_ctrls_1_down_DONT_FLUSH_PRECISE_4_0 = ((toplevel_decode_ctrls_1_down_Decode_INSTRUCTION_0 & 32'h00002050) == 32'h00002050);
  assign _zz_toplevel_decode_ctrls_1_down_DONT_FLUSH_PRECISE_4_0_1 = ((toplevel_decode_ctrls_1_down_Decode_INSTRUCTION_0 & 32'h00001050) == 32'h00001050);
  assign toplevel_decode_ctrls_1_down_DispatchPlugin_DONT_FLUSH_0 = _zz_toplevel_decode_ctrls_1_down_DispatchPlugin_DONT_FLUSH_0[0];
  assign toplevel_decode_ctrls_1_down_DispatchPlugin_DONT_FLUSH_FROM_LANES_0 = _zz_toplevel_decode_ctrls_1_down_DispatchPlugin_DONT_FLUSH_FROM_LANES_0[0];
  assign toplevel_decode_ctrls_1_down_DispatchPlugin_FENCE_OLDER_0 = _zz_toplevel_decode_ctrls_1_down_DispatchPlugin_FENCE_OLDER_0[0];
  assign toplevel_decode_ctrls_1_down_DONT_FLUSH_PRECISE_3_0 = _zz_toplevel_decode_ctrls_1_down_DONT_FLUSH_PRECISE_3_0[0];
  assign toplevel_decode_ctrls_1_down_DONT_FLUSH_PRECISE_4_0 = _zz_toplevel_decode_ctrls_1_down_DONT_FLUSH_PRECISE_4_0_2[0];
  assign toplevel_decode_ctrls_1_down_DecoderPlugin_logic_NEED_FPU_0 = _zz_toplevel_decode_ctrls_1_down_DecoderPlugin_logic_NEED_FPU_0[0];
  assign toplevel_decode_ctrls_1_down_DecoderPlugin_logic_NEED_RM_0 = _zz_toplevel_decode_ctrls_1_down_DecoderPlugin_logic_NEED_RM_0[0];
  assign toplevel_decode_ctrls_1_down_DispatchPlugin_logic_hcs_0_onRs_0_ENABLES_0_0 = _zz_toplevel_decode_ctrls_1_down_DispatchPlugin_logic_hcs_0_onRs_0_ENABLES_0_0[0];
  assign toplevel_decode_ctrls_1_down_DispatchPlugin_logic_hcs_0_onRs_1_ENABLES_0_0 = _zz_toplevel_decode_ctrls_1_down_DispatchPlugin_logic_hcs_0_onRs_1_ENABLES_0_0[0];
  assign toplevel_decode_ctrls_1_down_DispatchPlugin_logic_hcs_1_onRs_0_ENABLES_0_0 = _zz_toplevel_decode_ctrls_1_down_DispatchPlugin_logic_hcs_1_onRs_0_ENABLES_0_0[0];
  assign toplevel_decode_ctrls_1_down_DispatchPlugin_logic_hcs_1_onRs_1_ENABLES_0_0 = _zz_toplevel_decode_ctrls_1_down_DispatchPlugin_logic_hcs_1_onRs_1_ENABLES_0_0_1[0];
  assign toplevel_decode_ctrls_1_down_DispatchPlugin_logic_hcs_1_onRs_1_ENABLES_1_0 = _zz_toplevel_decode_ctrls_1_down_DispatchPlugin_logic_hcs_1_onRs_1_ENABLES_1_0[0];
  assign toplevel_decode_ctrls_1_down_DispatchPlugin_logic_hcs_2_onRs_0_ENABLES_0_0 = _zz_toplevel_decode_ctrls_1_down_DispatchPlugin_logic_hcs_2_onRs_0_ENABLES_0_0[0];
  assign toplevel_decode_ctrls_1_down_DispatchPlugin_logic_hcs_2_onRs_1_ENABLES_0_0 = _zz_toplevel_decode_ctrls_1_down_DispatchPlugin_logic_hcs_2_onRs_1_ENABLES_0_0[0];
  assign toplevel_decode_ctrls_1_down_DispatchPlugin_logic_hcs_3_onRs_0_ENABLES_0_0 = _zz_toplevel_decode_ctrls_1_down_DispatchPlugin_logic_hcs_3_onRs_0_ENABLES_0_0[0];
  assign toplevel_decode_ctrls_1_down_DispatchPlugin_logic_hcs_3_onRs_1_ENABLES_0_0 = _zz_toplevel_decode_ctrls_1_down_DispatchPlugin_logic_hcs_3_onRs_1_ENABLES_0_0_1[0];
  assign _zz_toplevel_decode_ctrls_1_down_DispatchPlugin_logic_LANES_LAYER_HIT_3_1_1 = ((toplevel_decode_ctrls_1_down_Decode_INSTRUCTION_1 & 32'h02000050) == 32'h00000010);
  assign _zz_toplevel_decode_ctrls_1_down_DispatchPlugin_logic_LANES_LAYER_HIT_3_1_2 = ((toplevel_decode_ctrls_1_down_Decode_INSTRUCTION_1 & 32'h00000030) == 32'h00000010);
  assign toplevel_decode_ctrls_1_down_DispatchPlugin_logic_LANES_LAYER_HIT_0_1 = _zz_toplevel_decode_ctrls_1_down_DispatchPlugin_logic_LANES_LAYER_HIT_0_1_2[0];
  assign _zz_toplevel_decode_ctrls_1_down_DispatchPlugin_logic_hcs_3_onRs_1_ENABLES_0_1 = ((toplevel_decode_ctrls_1_down_Decode_INSTRUCTION_1 & 32'h0) == 32'h0);
  assign toplevel_decode_ctrls_1_down_DispatchPlugin_logic_LANES_LAYER_HIT_1_1 = _zz_toplevel_decode_ctrls_1_down_DispatchPlugin_logic_LANES_LAYER_HIT_1_1[0];
  assign _zz_toplevel_decode_ctrls_1_down_DispatchPlugin_logic_LANES_LAYER_HIT_3_1_3 = ((toplevel_decode_ctrls_1_down_Decode_INSTRUCTION_1 & 32'h00000054) == 32'h00000040);
  assign _zz_toplevel_decode_ctrls_1_down_DispatchPlugin_logic_LANES_LAYER_HIT_3_1_4 = ((toplevel_decode_ctrls_1_down_Decode_INSTRUCTION_1 & 32'h0000004c) == 32'h00000004);
  assign toplevel_decode_ctrls_1_down_DispatchPlugin_logic_LANES_LAYER_HIT_2_1 = _zz_toplevel_decode_ctrls_1_down_DispatchPlugin_logic_LANES_LAYER_HIT_2_1[0];
  assign toplevel_decode_ctrls_1_down_DispatchPlugin_logic_LANES_LAYER_HIT_3_1 = _zz_toplevel_decode_ctrls_1_down_DispatchPlugin_logic_LANES_LAYER_HIT_3_1_5[0];
  assign _zz_toplevel_decode_ctrls_1_down_DispatchPlugin_logic_hcs_1_onRs_1_ENABLES_0_1 = ((toplevel_decode_ctrls_1_down_Decode_INSTRUCTION_1 & 32'h00000040) == 32'h00000040);
  assign toplevel_decode_ctrls_1_down_DispatchPlugin_MAY_FLUSH_1 = _zz_toplevel_decode_ctrls_1_down_DispatchPlugin_MAY_FLUSH_1_1[0];
  assign _zz_toplevel_decode_ctrls_1_down_DONT_FLUSH_PRECISE_4_1 = ((toplevel_decode_ctrls_1_down_Decode_INSTRUCTION_1 & 32'h00002050) == 32'h00002050);
  assign _zz_toplevel_decode_ctrls_1_down_DONT_FLUSH_PRECISE_4_1_1 = ((toplevel_decode_ctrls_1_down_Decode_INSTRUCTION_1 & 32'h00001050) == 32'h00001050);
  assign toplevel_decode_ctrls_1_down_DispatchPlugin_DONT_FLUSH_1 = _zz_toplevel_decode_ctrls_1_down_DispatchPlugin_DONT_FLUSH_1[0];
  assign toplevel_decode_ctrls_1_down_DispatchPlugin_DONT_FLUSH_FROM_LANES_1 = _zz_toplevel_decode_ctrls_1_down_DispatchPlugin_DONT_FLUSH_FROM_LANES_1[0];
  assign toplevel_decode_ctrls_1_down_DispatchPlugin_FENCE_OLDER_1 = _zz_toplevel_decode_ctrls_1_down_DispatchPlugin_FENCE_OLDER_1[0];
  assign toplevel_decode_ctrls_1_down_DONT_FLUSH_PRECISE_3_1 = _zz_toplevel_decode_ctrls_1_down_DONT_FLUSH_PRECISE_3_1[0];
  assign toplevel_decode_ctrls_1_down_DONT_FLUSH_PRECISE_4_1 = _zz_toplevel_decode_ctrls_1_down_DONT_FLUSH_PRECISE_4_1_2[0];
  assign toplevel_decode_ctrls_1_down_DecoderPlugin_logic_NEED_FPU_1 = _zz_toplevel_decode_ctrls_1_down_DecoderPlugin_logic_NEED_FPU_1[0];
  assign toplevel_decode_ctrls_1_down_DecoderPlugin_logic_NEED_RM_1 = _zz_toplevel_decode_ctrls_1_down_DecoderPlugin_logic_NEED_RM_1[0];
  assign toplevel_decode_ctrls_1_down_DispatchPlugin_logic_hcs_0_onRs_0_ENABLES_0_1 = _zz_toplevel_decode_ctrls_1_down_DispatchPlugin_logic_hcs_0_onRs_0_ENABLES_0_1[0];
  assign toplevel_decode_ctrls_1_down_DispatchPlugin_logic_hcs_0_onRs_1_ENABLES_0_1 = _zz_toplevel_decode_ctrls_1_down_DispatchPlugin_logic_hcs_0_onRs_1_ENABLES_0_1[0];
  assign toplevel_decode_ctrls_1_down_DispatchPlugin_logic_hcs_1_onRs_0_ENABLES_0_1 = _zz_toplevel_decode_ctrls_1_down_DispatchPlugin_logic_hcs_1_onRs_0_ENABLES_0_1[0];
  assign toplevel_decode_ctrls_1_down_DispatchPlugin_logic_hcs_1_onRs_1_ENABLES_0_1 = _zz_toplevel_decode_ctrls_1_down_DispatchPlugin_logic_hcs_1_onRs_1_ENABLES_0_1_1[0];
  assign toplevel_decode_ctrls_1_down_DispatchPlugin_logic_hcs_1_onRs_1_ENABLES_1_1 = _zz_toplevel_decode_ctrls_1_down_DispatchPlugin_logic_hcs_1_onRs_1_ENABLES_1_1[0];
  assign toplevel_decode_ctrls_1_down_DispatchPlugin_logic_hcs_2_onRs_0_ENABLES_0_1 = _zz_toplevel_decode_ctrls_1_down_DispatchPlugin_logic_hcs_2_onRs_0_ENABLES_0_1[0];
  assign toplevel_decode_ctrls_1_down_DispatchPlugin_logic_hcs_2_onRs_1_ENABLES_0_1 = _zz_toplevel_decode_ctrls_1_down_DispatchPlugin_logic_hcs_2_onRs_1_ENABLES_0_1[0];
  assign toplevel_decode_ctrls_1_down_DispatchPlugin_logic_hcs_3_onRs_0_ENABLES_0_1 = _zz_toplevel_decode_ctrls_1_down_DispatchPlugin_logic_hcs_3_onRs_0_ENABLES_0_1[0];
  assign toplevel_decode_ctrls_1_down_DispatchPlugin_logic_hcs_3_onRs_1_ENABLES_0_1 = _zz_toplevel_decode_ctrls_1_down_DispatchPlugin_logic_hcs_3_onRs_1_ENABLES_0_1_1[0];
  assign when_CtrlLaneApi_l46_4 = (toplevel_decode_ctrls_1_up_isReady || toplevel_decode_ctrls_1_lane0_upIsCancel);
  assign WhiteboxerPlugin_logic_serializeds_0_fire = (toplevel_decode_ctrls_1_up_LANE_SEL_0 && (! toplevel_decode_ctrls_1_up_LANE_SEL_0_regNext_1));
  assign WhiteboxerPlugin_logic_serializeds_0_decodeId = toplevel_decode_ctrls_1_down_Decode_DOP_ID_0;
  assign WhiteboxerPlugin_logic_serializeds_0_microOpId = toplevel_decode_ctrls_1_down_Decode_UOP_ID_0;
  assign WhiteboxerPlugin_logic_serializeds_0_microOp = toplevel_decode_ctrls_1_down_Decode_UOP_0;
  assign when_CtrlLaneApi_l46_5 = (toplevel_decode_ctrls_1_up_isReady || toplevel_decode_ctrls_1_lane1_upIsCancel);
  assign WhiteboxerPlugin_logic_serializeds_1_fire = (toplevel_decode_ctrls_1_up_LANE_SEL_1 && (! toplevel_decode_ctrls_1_up_LANE_SEL_1_regNext_1));
  assign WhiteboxerPlugin_logic_serializeds_1_decodeId = toplevel_decode_ctrls_1_down_Decode_DOP_ID_1;
  assign WhiteboxerPlugin_logic_serializeds_1_microOpId = toplevel_decode_ctrls_1_down_Decode_UOP_ID_1;
  assign WhiteboxerPlugin_logic_serializeds_1_microOp = toplevel_decode_ctrls_1_down_Decode_UOP_1;
  assign when_CtrlLaneApi_l46_6 = (toplevel_execute_ctrl0_down_isReady || toplevel_execute_lane0_ctrls_0_downIsCancel);
  assign WhiteboxerPlugin_logic_dispatches_0_fire = (toplevel_execute_ctrl0_down_LANE_SEL_lane0 && (! toplevel_execute_ctrl0_down_LANE_SEL_lane0_regNext));
  assign WhiteboxerPlugin_logic_dispatches_0_microOpId = toplevel_execute_ctrl0_down_Decode_UOP_ID_lane0;
  assign when_CtrlLaneApi_l46_7 = (toplevel_execute_ctrl0_down_isReady || toplevel_execute_lane1_ctrls_0_downIsCancel);
  assign WhiteboxerPlugin_logic_dispatches_1_fire = (toplevel_execute_ctrl0_down_LANE_SEL_lane1 && (! toplevel_execute_ctrl0_down_LANE_SEL_lane1_regNext));
  assign WhiteboxerPlugin_logic_dispatches_1_microOpId = toplevel_execute_ctrl0_down_Decode_UOP_ID_lane1;
  assign when_CtrlLaneApi_l46_8 = (toplevel_execute_ctrl2_down_isReady || toplevel_execute_lane0_ctrls_2_downIsCancel);
  assign WhiteboxerPlugin_logic_executes_0_fire = ((toplevel_execute_ctrl2_down_LANE_SEL_lane0 && (! toplevel_execute_ctrl2_down_LANE_SEL_lane0_regNext)) && toplevel_execute_ctrl2_down_COMMIT_lane0);
  assign WhiteboxerPlugin_logic_executes_0_microOpId = toplevel_execute_ctrl2_down_Decode_UOP_ID_lane0;
  assign when_CtrlLaneApi_l46_9 = (toplevel_execute_ctrl2_down_isReady || toplevel_execute_lane1_ctrls_2_downIsCancel);
  assign WhiteboxerPlugin_logic_executes_1_fire = ((toplevel_execute_ctrl2_down_LANE_SEL_lane1 && (! toplevel_execute_ctrl2_down_LANE_SEL_lane1_regNext)) && toplevel_execute_ctrl2_down_COMMIT_lane1);
  assign WhiteboxerPlugin_logic_executes_1_microOpId = toplevel_execute_ctrl2_down_Decode_UOP_ID_lane1;
  assign BtbPlugin_logic_onForget_hash = DecoderPlugin_logic_forgetPort_payload_pcOnLastSlice[26 : 11];
  assign _zz_BtbPlugin_logic_readPort_rsp_0_hash = BtbPlugin_logic_mem_spinal_port1;
  assign _zz_BtbPlugin_logic_readPort_rsp_0_hash_1 = _zz_BtbPlugin_logic_readPort_rsp_0_hash[50 : 0];
  assign _zz_BtbPlugin_logic_readPort_rsp_1_hash = _zz_BtbPlugin_logic_readPort_rsp_0_hash[101 : 51];
  assign BtbPlugin_logic_readPort_rsp_0_hash = _zz_BtbPlugin_logic_readPort_rsp_0_hash_1[15 : 0];
  assign BtbPlugin_logic_readPort_rsp_0_sliceLow = _zz_BtbPlugin_logic_readPort_rsp_0_hash_1[16 : 16];
  assign BtbPlugin_logic_readPort_rsp_0_pcTarget = _zz_BtbPlugin_logic_readPort_rsp_0_hash_1[47 : 17];
  assign BtbPlugin_logic_readPort_rsp_0_isBranch = _zz_BtbPlugin_logic_readPort_rsp_0_hash_1[48];
  assign BtbPlugin_logic_readPort_rsp_0_isPush = _zz_BtbPlugin_logic_readPort_rsp_0_hash_1[49];
  assign BtbPlugin_logic_readPort_rsp_0_isPop = _zz_BtbPlugin_logic_readPort_rsp_0_hash_1[50];
  assign BtbPlugin_logic_readPort_rsp_1_hash = _zz_BtbPlugin_logic_readPort_rsp_1_hash[15 : 0];
  assign BtbPlugin_logic_readPort_rsp_1_sliceLow = _zz_BtbPlugin_logic_readPort_rsp_1_hash[16 : 16];
  assign BtbPlugin_logic_readPort_rsp_1_pcTarget = _zz_BtbPlugin_logic_readPort_rsp_1_hash[47 : 17];
  assign BtbPlugin_logic_readPort_rsp_1_isBranch = _zz_BtbPlugin_logic_readPort_rsp_1_hash[48];
  assign BtbPlugin_logic_readPort_rsp_1_isPush = _zz_BtbPlugin_logic_readPort_rsp_1_hash[49];
  assign BtbPlugin_logic_readPort_rsp_1_isPop = _zz_BtbPlugin_logic_readPort_rsp_1_hash[50];
  assign BtbPlugin_logic_readPort_cmd_valid = fetch_logic_ctrls_0_down_isReady;
  assign BtbPlugin_logic_readPort_cmd_payload = _zz_BtbPlugin_logic_readPort_cmd_payload[7:0];
  assign fetch_logic_ctrls_0_down_BtbPlugin_logic_readCmd_HAZARDS = ((BtbPlugin_logic_onLearn_port_valid && (BtbPlugin_logic_onLearn_port_payload_address == BtbPlugin_logic_readPort_cmd_payload)) ? BtbPlugin_logic_onLearn_port_payload_mask : 2'b00);
  assign fetch_logic_ctrls_0_haltRequest_BtbPlugin_l171 = BtbPlugin_logic_onLearn_port_valid;
  assign BtbPlugin_logic_predictions = {fetch_logic_ctrls_2_down_GSharePlugin_GSHARE_COUNTER_3[1],{fetch_logic_ctrls_2_down_GSharePlugin_GSHARE_COUNTER_2[1],{fetch_logic_ctrls_2_down_GSharePlugin_GSHARE_COUNTER_1[1],fetch_logic_ctrls_2_down_GSharePlugin_GSHARE_COUNTER_0[1]}}};
  assign fetch_logic_ctrls_1_down_BtbPlugin_logic_chunksLogic_0_readRsp_ENTRY_hash = BtbPlugin_logic_readPort_rsp_0_hash;
  assign fetch_logic_ctrls_1_down_BtbPlugin_logic_chunksLogic_0_readRsp_ENTRY_sliceLow = BtbPlugin_logic_readPort_rsp_0_sliceLow;
  assign fetch_logic_ctrls_1_down_BtbPlugin_logic_chunksLogic_0_readRsp_ENTRY_pcTarget = BtbPlugin_logic_readPort_rsp_0_pcTarget;
  assign fetch_logic_ctrls_1_down_BtbPlugin_logic_chunksLogic_0_readRsp_ENTRY_isBranch = BtbPlugin_logic_readPort_rsp_0_isBranch;
  assign fetch_logic_ctrls_1_down_BtbPlugin_logic_chunksLogic_0_readRsp_ENTRY_isPush = BtbPlugin_logic_readPort_rsp_0_isPush;
  assign fetch_logic_ctrls_1_down_BtbPlugin_logic_chunksLogic_0_readRsp_ENTRY_isPop = BtbPlugin_logic_readPort_rsp_0_isPop;
  assign fetch_logic_ctrls_1_down_BtbPlugin_logic_chunksLogic_0_hitCalc_HIT = ((fetch_logic_ctrls_1_down_BtbPlugin_logic_chunksLogic_0_readRsp_ENTRY_hash == fetch_logic_ctrls_1_down_Fetch_WORD_PC[26 : 11]) && (fetch_logic_ctrls_1_down_Fetch_WORD_PC[2 : 1] <= {1'b0,fetch_logic_ctrls_1_down_BtbPlugin_logic_chunksLogic_0_readRsp_ENTRY_sliceLow}));
  assign fetch_logic_ctrls_2_down_BtbPlugin_logic_chunksLogic_0_predict_TAKEN = ((! fetch_logic_ctrls_2_down_BtbPlugin_logic_chunksLogic_0_readRsp_ENTRY_isBranch) || BtbPlugin_logic_predictions[{1'b0,fetch_logic_ctrls_2_down_BtbPlugin_logic_chunksLogic_0_readRsp_ENTRY_sliceLow}]);
  assign fetch_logic_ctrls_1_down_BtbPlugin_logic_chunksLogic_1_readRsp_ENTRY_hash = BtbPlugin_logic_readPort_rsp_1_hash;
  assign fetch_logic_ctrls_1_down_BtbPlugin_logic_chunksLogic_1_readRsp_ENTRY_sliceLow = BtbPlugin_logic_readPort_rsp_1_sliceLow;
  assign fetch_logic_ctrls_1_down_BtbPlugin_logic_chunksLogic_1_readRsp_ENTRY_pcTarget = BtbPlugin_logic_readPort_rsp_1_pcTarget;
  assign fetch_logic_ctrls_1_down_BtbPlugin_logic_chunksLogic_1_readRsp_ENTRY_isBranch = BtbPlugin_logic_readPort_rsp_1_isBranch;
  assign fetch_logic_ctrls_1_down_BtbPlugin_logic_chunksLogic_1_readRsp_ENTRY_isPush = BtbPlugin_logic_readPort_rsp_1_isPush;
  assign fetch_logic_ctrls_1_down_BtbPlugin_logic_chunksLogic_1_readRsp_ENTRY_isPop = BtbPlugin_logic_readPort_rsp_1_isPop;
  assign fetch_logic_ctrls_1_down_BtbPlugin_logic_chunksLogic_1_hitCalc_HIT = ((fetch_logic_ctrls_1_down_BtbPlugin_logic_chunksLogic_1_readRsp_ENTRY_hash == fetch_logic_ctrls_1_down_Fetch_WORD_PC[26 : 11]) && (fetch_logic_ctrls_1_down_Fetch_WORD_PC[2 : 1] <= {1'b1,fetch_logic_ctrls_1_down_BtbPlugin_logic_chunksLogic_1_readRsp_ENTRY_sliceLow}));
  assign fetch_logic_ctrls_2_down_BtbPlugin_logic_chunksLogic_1_predict_TAKEN = ((! fetch_logic_ctrls_2_down_BtbPlugin_logic_chunksLogic_1_readRsp_ENTRY_isBranch) || BtbPlugin_logic_predictions[{1'b1,fetch_logic_ctrls_2_down_BtbPlugin_logic_chunksLogic_1_readRsp_ENTRY_sliceLow}]);
  assign BtbPlugin_logic_ras_readIt = fetch_logic_ctrls_1_down_isReady;
  assign BtbPlugin_logic_applyIt_chunksMask = {(fetch_logic_ctrls_2_down_BtbPlugin_logic_chunksLogic_1_hitCalc_HIT && ((fetch_logic_ctrls_2_down_BtbPlugin_logic_chunksLogic_0_hitCalc_HIT && fetch_logic_ctrls_2_down_BtbPlugin_logic_chunksLogic_0_predict_TAKEN) == 1'b0)),(fetch_logic_ctrls_2_down_BtbPlugin_logic_chunksLogic_0_hitCalc_HIT && 1'b1)};
  assign BtbPlugin_logic_applyIt_chunksTakenOh = ({fetch_logic_ctrls_2_down_BtbPlugin_logic_chunksLogic_1_predict_TAKEN,fetch_logic_ctrls_2_down_BtbPlugin_logic_chunksLogic_0_predict_TAKEN} & BtbPlugin_logic_applyIt_chunksMask);
  assign BtbPlugin_logic_applyIt_needIt = (fetch_logic_ctrls_2_up_isValid && (|BtbPlugin_logic_applyIt_chunksTakenOh));
  assign when_BtbPlugin_l205 = (fetch_logic_ctrls_2_up_isReady || fetch_logic_ctrls_2_up_isCancel);
  assign BtbPlugin_logic_applyIt_doIt = (BtbPlugin_logic_applyIt_needIt && (! BtbPlugin_logic_applyIt_correctionSent));
  assign _zz_BtbPlugin_logic_applyIt_doItSlice = BtbPlugin_logic_applyIt_chunksTakenOh[1];
  assign _zz_BtbPlugin_logic_applyIt_entry_hash = ((BtbPlugin_logic_applyIt_chunksTakenOh[0] ? {fetch_logic_ctrls_2_down_BtbPlugin_logic_chunksLogic_0_readRsp_ENTRY_isPop,{fetch_logic_ctrls_2_down_BtbPlugin_logic_chunksLogic_0_readRsp_ENTRY_isPush,{fetch_logic_ctrls_2_down_BtbPlugin_logic_chunksLogic_0_readRsp_ENTRY_isBranch,{_zz__zz_BtbPlugin_logic_applyIt_entry_hash,_zz__zz_BtbPlugin_logic_applyIt_entry_hash_1}}}} : 51'h0) | (_zz_BtbPlugin_logic_applyIt_doItSlice ? {fetch_logic_ctrls_2_down_BtbPlugin_logic_chunksLogic_1_readRsp_ENTRY_isPop,{fetch_logic_ctrls_2_down_BtbPlugin_logic_chunksLogic_1_readRsp_ENTRY_isPush,{fetch_logic_ctrls_2_down_BtbPlugin_logic_chunksLogic_1_readRsp_ENTRY_isBranch,{_zz__zz_BtbPlugin_logic_applyIt_entry_hash_2,_zz__zz_BtbPlugin_logic_applyIt_entry_hash_3}}}} : 51'h0));
  assign BtbPlugin_logic_applyIt_entry_hash = _zz_BtbPlugin_logic_applyIt_entry_hash[15 : 0];
  assign BtbPlugin_logic_applyIt_entry_sliceLow = _zz_BtbPlugin_logic_applyIt_entry_hash[16 : 16];
  assign BtbPlugin_logic_applyIt_entry_pcTarget = _zz_BtbPlugin_logic_applyIt_entry_hash[47 : 17];
  assign BtbPlugin_logic_applyIt_entry_isBranch = _zz_BtbPlugin_logic_applyIt_entry_hash[48];
  assign BtbPlugin_logic_applyIt_entry_isPush = _zz_BtbPlugin_logic_applyIt_entry_hash[49];
  assign BtbPlugin_logic_applyIt_entry_isPop = _zz_BtbPlugin_logic_applyIt_entry_hash[50];
  always @(*) begin
    BtbPlugin_logic_applyIt_pcTarget = BtbPlugin_logic_applyIt_entry_pcTarget;
    if(BtbPlugin_logic_applyIt_entry_isPop) begin
      BtbPlugin_logic_applyIt_pcTarget = BtbPlugin_logic_ras_read;
    end
  end

  assign BtbPlugin_logic_applyIt_doItSlice = {_zz_BtbPlugin_logic_applyIt_doItSlice,BtbPlugin_logic_applyIt_entry_sliceLow};
  assign BtbPlugin_logic_applyIt_rasLogic_pushValid = (BtbPlugin_logic_applyIt_doIt && BtbPlugin_logic_applyIt_entry_isPush);
  always @(*) begin
    BtbPlugin_logic_applyIt_rasLogic_pushPc = fetch_logic_ctrls_2_down_Fetch_WORD_PC;
    BtbPlugin_logic_applyIt_rasLogic_pushPc[2 : 1] = BtbPlugin_logic_applyIt_doItSlice;
  end

  assign when_BtbPlugin_l218 = (BtbPlugin_logic_applyIt_doIt && BtbPlugin_logic_applyIt_entry_isPop);
  assign BtbPlugin_logic_flushPort_valid = BtbPlugin_logic_applyIt_doIt;
  assign BtbPlugin_logic_flushPort_payload_self = 1'b0;
  assign BtbPlugin_logic_pcPort_valid = BtbPlugin_logic_applyIt_doIt;
  assign BtbPlugin_logic_pcPort_payload_fault = 1'b0;
  assign BtbPlugin_logic_pcPort_payload_pc = ({1'd0,BtbPlugin_logic_applyIt_pcTarget} <<< 1'd1);
  assign fetch_logic_ctrls_2_down_Prediction_WORD_JUMPED = BtbPlugin_logic_applyIt_needIt;
  assign fetch_logic_ctrls_2_down_Prediction_WORD_JUMP_SLICE = BtbPlugin_logic_applyIt_doItSlice;
  assign fetch_logic_ctrls_2_down_Prediction_WORD_JUMP_PC = ({1'd0,BtbPlugin_logic_applyIt_pcTarget} <<< 1'd1);
  assign BtbPlugin_logic_applyIt_history_layers_0_history = fetch_logic_ctrls_2_down_Prediction_BRANCH_HISTORY;
  assign BtbPlugin_logic_applyIt_history_layersLogic_0_doIt = (BtbPlugin_logic_applyIt_chunksMask[0] && fetch_logic_ctrls_2_down_BtbPlugin_logic_chunksLogic_0_readRsp_ENTRY_isBranch);
  assign BtbPlugin_logic_applyIt_history_layersLogic_0_shifted = {BtbPlugin_logic_applyIt_history_layers_0_history[10 : 0],fetch_logic_ctrls_2_down_BtbPlugin_logic_chunksLogic_0_predict_TAKEN};
  assign BtbPlugin_logic_applyIt_history_layers_1_history = (BtbPlugin_logic_applyIt_history_layersLogic_0_doIt ? BtbPlugin_logic_applyIt_history_layersLogic_0_shifted : BtbPlugin_logic_applyIt_history_layers_0_history);
  assign BtbPlugin_logic_applyIt_history_layersLogic_1_doIt = (BtbPlugin_logic_applyIt_chunksMask[1] && fetch_logic_ctrls_2_down_BtbPlugin_logic_chunksLogic_1_readRsp_ENTRY_isBranch);
  assign BtbPlugin_logic_applyIt_history_layersLogic_1_shifted = {BtbPlugin_logic_applyIt_history_layers_1_history[10 : 0],fetch_logic_ctrls_2_down_BtbPlugin_logic_chunksLogic_1_predict_TAKEN};
  assign BtbPlugin_logic_applyIt_history_layers_2_history = (BtbPlugin_logic_applyIt_history_layersLogic_1_doIt ? BtbPlugin_logic_applyIt_history_layersLogic_1_shifted : BtbPlugin_logic_applyIt_history_layers_1_history);
  assign BtbPlugin_logic_historyPort_valid = ((fetch_logic_ctrls_2_up_isValid && (! BtbPlugin_logic_applyIt_correctionSent)) && (|{fetch_logic_ctrls_2_down_BtbPlugin_logic_chunksLogic_1_hitCalc_HIT,fetch_logic_ctrls_2_down_BtbPlugin_logic_chunksLogic_0_hitCalc_HIT}));
  assign BtbPlugin_logic_historyPort_payload_history = BtbPlugin_logic_applyIt_history_layers_2_history;
  always @(*) begin
    fetch_logic_ctrls_2_down_Prediction_WORD_SLICES_BRANCH[0] = ((fetch_logic_ctrls_2_down_BtbPlugin_logic_chunksLogic_0_hitCalc_HIT && fetch_logic_ctrls_2_down_BtbPlugin_logic_chunksLogic_0_readRsp_ENTRY_isBranch) && (fetch_logic_ctrls_2_down_BtbPlugin_logic_chunksLogic_0_readRsp_ENTRY_sliceLow == 1'b0));
    fetch_logic_ctrls_2_down_Prediction_WORD_SLICES_BRANCH[1] = ((fetch_logic_ctrls_2_down_BtbPlugin_logic_chunksLogic_0_hitCalc_HIT && fetch_logic_ctrls_2_down_BtbPlugin_logic_chunksLogic_0_readRsp_ENTRY_isBranch) && (fetch_logic_ctrls_2_down_BtbPlugin_logic_chunksLogic_0_readRsp_ENTRY_sliceLow == 1'b1));
    fetch_logic_ctrls_2_down_Prediction_WORD_SLICES_BRANCH[2] = ((fetch_logic_ctrls_2_down_BtbPlugin_logic_chunksLogic_1_hitCalc_HIT && fetch_logic_ctrls_2_down_BtbPlugin_logic_chunksLogic_1_readRsp_ENTRY_isBranch) && (fetch_logic_ctrls_2_down_BtbPlugin_logic_chunksLogic_1_readRsp_ENTRY_sliceLow == 1'b0));
    fetch_logic_ctrls_2_down_Prediction_WORD_SLICES_BRANCH[3] = ((fetch_logic_ctrls_2_down_BtbPlugin_logic_chunksLogic_1_hitCalc_HIT && fetch_logic_ctrls_2_down_BtbPlugin_logic_chunksLogic_1_readRsp_ENTRY_isBranch) && (fetch_logic_ctrls_2_down_BtbPlugin_logic_chunksLogic_1_readRsp_ENTRY_sliceLow == 1'b1));
  end

  always @(*) begin
    fetch_logic_ctrls_2_down_Prediction_WORD_SLICES_TAKEN[0] = fetch_logic_ctrls_2_down_BtbPlugin_logic_chunksLogic_0_predict_TAKEN;
    fetch_logic_ctrls_2_down_Prediction_WORD_SLICES_TAKEN[1] = fetch_logic_ctrls_2_down_BtbPlugin_logic_chunksLogic_0_predict_TAKEN;
    fetch_logic_ctrls_2_down_Prediction_WORD_SLICES_TAKEN[2] = fetch_logic_ctrls_2_down_BtbPlugin_logic_chunksLogic_1_predict_TAKEN;
    fetch_logic_ctrls_2_down_Prediction_WORD_SLICES_TAKEN[3] = fetch_logic_ctrls_2_down_BtbPlugin_logic_chunksLogic_1_predict_TAKEN;
  end

  assign BtbPlugin_logic_initializer_busy = (! BtbPlugin_logic_initializer_counter[8]);
  assign AlignerPlugin_logic_buffer_flushIt = (|{(DecoderPlugin_logic_laneLogic_1_flushPort_valid && 1'b1),{(DecoderPlugin_logic_laneLogic_0_flushPort_valid && 1'b1),{(late1_BranchPlugin_logic_flushPort_valid && 1'b1),{(early1_BranchPlugin_logic_flushPort_valid && 1'b1),{(late0_BranchPlugin_logic_flushPort_valid && _zz_AlignerPlugin_logic_buffer_flushIt),{_zz_AlignerPlugin_logic_buffer_flushIt_1,{_zz_AlignerPlugin_logic_buffer_flushIt_2,_zz_AlignerPlugin_logic_buffer_flushIt_3}}}}}}});
  assign AlignerPlugin_logic_buffer_readers_0_firstFromBuffer = (|{_zz_AlignerPlugin_logic_extractors_0_redo_3,{_zz_AlignerPlugin_logic_extractors_0_redo_2,{_zz_AlignerPlugin_logic_extractors_0_redo_1,_zz_AlignerPlugin_logic_extractors_0_redo}}});
  assign AlignerPlugin_logic_buffer_readers_0_lastFromBuffer = ({AlignerPlugin_logic_extractors_0_usageMask[7],{AlignerPlugin_logic_extractors_0_usageMask[6],{AlignerPlugin_logic_extractors_0_usageMask[5],AlignerPlugin_logic_extractors_0_usageMask[4]}}} == 4'b0000);
  assign _zz_AlignerPlugin_logic_extractors_0_ctx_instruction = {_zz_AlignerPlugin_logic_extractors_0_redo_7,{_zz_AlignerPlugin_logic_extractors_0_redo_6,{_zz_AlignerPlugin_logic_extractors_0_redo_5,{_zz_AlignerPlugin_logic_extractors_0_redo_4,{_zz_AlignerPlugin_logic_extractors_0_redo_3,{_zz_AlignerPlugin_logic_extractors_0_redo_2,{_zz_AlignerPlugin_logic_extractors_0_redo_1,_zz_AlignerPlugin_logic_extractors_0_redo}}}}}}};
  assign AlignerPlugin_logic_extractors_0_ctx_instruction = ((((_zz_AlignerPlugin_logic_extractors_0_ctx_instruction_1 ? AlignerPlugin_logic_slicesInstructions_0 : _zz_AlignerPlugin_logic_extractors_0_ctx_instruction_2) | (_zz_AlignerPlugin_logic_extractors_0_ctx_instruction_3 ? AlignerPlugin_logic_slicesInstructions_1 : _zz_AlignerPlugin_logic_extractors_0_ctx_instruction_4)) | ((_zz_AlignerPlugin_logic_extractors_0_ctx_instruction_5 ? AlignerPlugin_logic_slicesInstructions_2 : _zz_AlignerPlugin_logic_extractors_0_ctx_instruction_6) | (_zz_AlignerPlugin_logic_extractors_0_ctx_instruction_7 ? AlignerPlugin_logic_slicesInstructions_3 : _zz_AlignerPlugin_logic_extractors_0_ctx_instruction_8))) | (((_zz_AlignerPlugin_logic_extractors_0_ctx_instruction_9 ? AlignerPlugin_logic_slicesInstructions_4 : _zz_AlignerPlugin_logic_extractors_0_ctx_instruction_10) | (_zz_AlignerPlugin_logic_extractors_0_ctx_instruction_11 ? AlignerPlugin_logic_slicesInstructions_5 : _zz_AlignerPlugin_logic_extractors_0_ctx_instruction_12)) | ((_zz_AlignerPlugin_logic_extractors_0_ctx_instruction_13 ? AlignerPlugin_logic_slicesInstructions_6 : _zz_AlignerPlugin_logic_extractors_0_ctx_instruction_14) | (_zz_AlignerPlugin_logic_extractors_0_ctx_instruction_15 ? AlignerPlugin_logic_slicesInstructions_7 : _zz_AlignerPlugin_logic_extractors_0_ctx_instruction_16))));
  always @(*) begin
    AlignerPlugin_logic_extractors_0_ctx_pc = (AlignerPlugin_logic_buffer_readers_0_firstFromBuffer ? AlignerPlugin_logic_buffer_pc : fetch_logic_ctrls_2_down_Fetch_WORD_PC);
    AlignerPlugin_logic_extractors_0_ctx_pc[2 : 1] = {_zz_AlignerPlugin_logic_extractors_0_ctx_pc_2,_zz_AlignerPlugin_logic_extractors_0_ctx_pc_1};
  end

  assign _zz_AlignerPlugin_logic_extractors_0_ctx_pc = (|{_zz_AlignerPlugin_logic_extractors_0_redo_7,_zz_AlignerPlugin_logic_extractors_0_redo_3});
  assign _zz_AlignerPlugin_logic_extractors_0_ctx_pc_1 = ((|{_zz_AlignerPlugin_logic_extractors_0_redo_5,_zz_AlignerPlugin_logic_extractors_0_redo_1}) || _zz_AlignerPlugin_logic_extractors_0_ctx_pc);
  assign _zz_AlignerPlugin_logic_extractors_0_ctx_pc_2 = ((|{_zz_AlignerPlugin_logic_extractors_0_redo_6,_zz_AlignerPlugin_logic_extractors_0_redo_2}) || _zz_AlignerPlugin_logic_extractors_0_ctx_pc);
  assign AlignerPlugin_logic_extractors_0_ctx_trap = ((AlignerPlugin_logic_buffer_readers_0_firstFromBuffer && AlignerPlugin_logic_buffer_trap) || ((! AlignerPlugin_logic_buffer_readers_0_lastFromBuffer) && fetch_logic_ctrls_2_down_TRAP));
  assign AlignerPlugin_logic_extractors_0_ctx_hm_Fetch_ID = (AlignerPlugin_logic_buffer_readers_0_firstFromBuffer ? AlignerPlugin_logic_buffer_hm_Fetch_ID : fetch_logic_ctrls_2_down_Fetch_ID);
  assign AlignerPlugin_logic_extractors_0_ctx_hm_GSharePlugin_GSHARE_COUNTER_0 = (AlignerPlugin_logic_buffer_readers_0_lastFromBuffer ? AlignerPlugin_logic_buffer_hm_GSharePlugin_GSHARE_COUNTER_0 : fetch_logic_ctrls_2_down_GSharePlugin_GSHARE_COUNTER_0);
  assign AlignerPlugin_logic_extractors_0_ctx_hm_GSharePlugin_GSHARE_COUNTER_1 = (AlignerPlugin_logic_buffer_readers_0_lastFromBuffer ? AlignerPlugin_logic_buffer_hm_GSharePlugin_GSHARE_COUNTER_1 : fetch_logic_ctrls_2_down_GSharePlugin_GSHARE_COUNTER_1);
  assign AlignerPlugin_logic_extractors_0_ctx_hm_GSharePlugin_GSHARE_COUNTER_2 = (AlignerPlugin_logic_buffer_readers_0_lastFromBuffer ? AlignerPlugin_logic_buffer_hm_GSharePlugin_GSHARE_COUNTER_2 : fetch_logic_ctrls_2_down_GSharePlugin_GSHARE_COUNTER_2);
  assign AlignerPlugin_logic_extractors_0_ctx_hm_GSharePlugin_GSHARE_COUNTER_3 = (AlignerPlugin_logic_buffer_readers_0_lastFromBuffer ? AlignerPlugin_logic_buffer_hm_GSharePlugin_GSHARE_COUNTER_3 : fetch_logic_ctrls_2_down_GSharePlugin_GSHARE_COUNTER_3);
  assign AlignerPlugin_logic_extractors_0_ctx_hm_Prediction_BRANCH_HISTORY = (AlignerPlugin_logic_buffer_readers_0_lastFromBuffer ? AlignerPlugin_logic_buffer_hm_Prediction_BRANCH_HISTORY : fetch_logic_ctrls_2_down_Prediction_BRANCH_HISTORY);
  assign AlignerPlugin_logic_extractors_0_ctx_hm_Prediction_WORD_SLICES_BRANCH = (AlignerPlugin_logic_buffer_readers_0_lastFromBuffer ? AlignerPlugin_logic_buffer_hm_Prediction_WORD_SLICES_BRANCH : fetch_logic_ctrls_2_down_Prediction_WORD_SLICES_BRANCH);
  assign AlignerPlugin_logic_extractors_0_ctx_hm_Prediction_WORD_SLICES_TAKEN = (AlignerPlugin_logic_buffer_readers_0_lastFromBuffer ? AlignerPlugin_logic_buffer_hm_Prediction_WORD_SLICES_TAKEN : fetch_logic_ctrls_2_down_Prediction_WORD_SLICES_TAKEN);
  assign AlignerPlugin_logic_extractors_0_ctx_hm_Prediction_WORD_JUMP_PC = (AlignerPlugin_logic_buffer_readers_0_lastFromBuffer ? AlignerPlugin_logic_buffer_hm_Prediction_WORD_JUMP_PC : fetch_logic_ctrls_2_down_Prediction_WORD_JUMP_PC);
  assign AlignerPlugin_logic_extractors_0_ctx_hm_Prediction_WORD_JUMPED = (AlignerPlugin_logic_buffer_readers_0_lastFromBuffer ? AlignerPlugin_logic_buffer_hm_Prediction_WORD_JUMPED : fetch_logic_ctrls_2_down_Prediction_WORD_JUMPED);
  assign AlignerPlugin_logic_extractors_0_ctx_hm_Prediction_WORD_JUMP_SLICE = (AlignerPlugin_logic_buffer_readers_0_lastFromBuffer ? AlignerPlugin_logic_buffer_hm_Prediction_WORD_JUMP_SLICE : fetch_logic_ctrls_2_down_Prediction_WORD_JUMP_SLICE);
  assign AlignerPlugin_logic_buffer_readers_1_firstFromBuffer = (|{_zz_AlignerPlugin_logic_extractors_1_redo_2,{_zz_AlignerPlugin_logic_extractors_1_redo_1,_zz_AlignerPlugin_logic_extractors_1_redo}});
  assign AlignerPlugin_logic_buffer_readers_1_lastFromBuffer = ({AlignerPlugin_logic_extractors_1_usageMask[7],{AlignerPlugin_logic_extractors_1_usageMask[6],{AlignerPlugin_logic_extractors_1_usageMask[5],AlignerPlugin_logic_extractors_1_usageMask[4]}}} == 4'b0000);
  assign _zz_AlignerPlugin_logic_extractors_1_ctx_instruction = {_zz_AlignerPlugin_logic_extractors_1_redo_6,{_zz_AlignerPlugin_logic_extractors_1_redo_5,{_zz_AlignerPlugin_logic_extractors_1_redo_4,{_zz_AlignerPlugin_logic_extractors_1_redo_3,{_zz_AlignerPlugin_logic_extractors_1_redo_2,{_zz_AlignerPlugin_logic_extractors_1_redo_1,_zz_AlignerPlugin_logic_extractors_1_redo}}}}}};
  assign AlignerPlugin_logic_extractors_1_ctx_instruction = ((((_zz_AlignerPlugin_logic_extractors_1_ctx_instruction[0] ? AlignerPlugin_logic_slicesInstructions_1 : 32'h0) | (_zz_AlignerPlugin_logic_extractors_1_ctx_instruction[1] ? AlignerPlugin_logic_slicesInstructions_2 : 32'h0)) | ((_zz_AlignerPlugin_logic_extractors_1_ctx_instruction[2] ? AlignerPlugin_logic_slicesInstructions_3 : 32'h0) | (_zz_AlignerPlugin_logic_extractors_1_ctx_instruction[3] ? AlignerPlugin_logic_slicesInstructions_4 : 32'h0))) | (((_zz_AlignerPlugin_logic_extractors_1_ctx_instruction[4] ? AlignerPlugin_logic_slicesInstructions_5 : 32'h0) | (_zz_AlignerPlugin_logic_extractors_1_ctx_instruction[5] ? AlignerPlugin_logic_slicesInstructions_6 : 32'h0)) | (_zz_AlignerPlugin_logic_extractors_1_ctx_instruction[6] ? AlignerPlugin_logic_slicesInstructions_7 : 32'h0)));
  always @(*) begin
    AlignerPlugin_logic_extractors_1_ctx_pc = (AlignerPlugin_logic_buffer_readers_1_firstFromBuffer ? AlignerPlugin_logic_buffer_pc : fetch_logic_ctrls_2_down_Fetch_WORD_PC);
    AlignerPlugin_logic_extractors_1_ctx_pc[2 : 1] = {_zz_AlignerPlugin_logic_extractors_1_ctx_pc_2,_zz_AlignerPlugin_logic_extractors_1_ctx_pc_1};
  end

  assign _zz_AlignerPlugin_logic_extractors_1_ctx_pc = (|{_zz_AlignerPlugin_logic_extractors_1_redo_6,_zz_AlignerPlugin_logic_extractors_1_redo_2});
  assign _zz_AlignerPlugin_logic_extractors_1_ctx_pc_1 = ((|{_zz_AlignerPlugin_logic_extractors_1_redo_4,_zz_AlignerPlugin_logic_extractors_1_redo}) || _zz_AlignerPlugin_logic_extractors_1_ctx_pc);
  assign _zz_AlignerPlugin_logic_extractors_1_ctx_pc_2 = ((|{_zz_AlignerPlugin_logic_extractors_1_redo_5,_zz_AlignerPlugin_logic_extractors_1_redo_1}) || _zz_AlignerPlugin_logic_extractors_1_ctx_pc);
  assign AlignerPlugin_logic_extractors_1_ctx_trap = ((AlignerPlugin_logic_buffer_readers_1_firstFromBuffer && AlignerPlugin_logic_buffer_trap) || ((! AlignerPlugin_logic_buffer_readers_1_lastFromBuffer) && fetch_logic_ctrls_2_down_TRAP));
  assign AlignerPlugin_logic_extractors_1_ctx_hm_Fetch_ID = (AlignerPlugin_logic_buffer_readers_1_firstFromBuffer ? AlignerPlugin_logic_buffer_hm_Fetch_ID : fetch_logic_ctrls_2_down_Fetch_ID);
  assign AlignerPlugin_logic_extractors_1_ctx_hm_GSharePlugin_GSHARE_COUNTER_0 = (AlignerPlugin_logic_buffer_readers_1_lastFromBuffer ? AlignerPlugin_logic_buffer_hm_GSharePlugin_GSHARE_COUNTER_0 : fetch_logic_ctrls_2_down_GSharePlugin_GSHARE_COUNTER_0);
  assign AlignerPlugin_logic_extractors_1_ctx_hm_GSharePlugin_GSHARE_COUNTER_1 = (AlignerPlugin_logic_buffer_readers_1_lastFromBuffer ? AlignerPlugin_logic_buffer_hm_GSharePlugin_GSHARE_COUNTER_1 : fetch_logic_ctrls_2_down_GSharePlugin_GSHARE_COUNTER_1);
  assign AlignerPlugin_logic_extractors_1_ctx_hm_GSharePlugin_GSHARE_COUNTER_2 = (AlignerPlugin_logic_buffer_readers_1_lastFromBuffer ? AlignerPlugin_logic_buffer_hm_GSharePlugin_GSHARE_COUNTER_2 : fetch_logic_ctrls_2_down_GSharePlugin_GSHARE_COUNTER_2);
  assign AlignerPlugin_logic_extractors_1_ctx_hm_GSharePlugin_GSHARE_COUNTER_3 = (AlignerPlugin_logic_buffer_readers_1_lastFromBuffer ? AlignerPlugin_logic_buffer_hm_GSharePlugin_GSHARE_COUNTER_3 : fetch_logic_ctrls_2_down_GSharePlugin_GSHARE_COUNTER_3);
  assign AlignerPlugin_logic_extractors_1_ctx_hm_Prediction_BRANCH_HISTORY = (AlignerPlugin_logic_buffer_readers_1_lastFromBuffer ? AlignerPlugin_logic_buffer_hm_Prediction_BRANCH_HISTORY : fetch_logic_ctrls_2_down_Prediction_BRANCH_HISTORY);
  assign AlignerPlugin_logic_extractors_1_ctx_hm_Prediction_WORD_SLICES_BRANCH = (AlignerPlugin_logic_buffer_readers_1_lastFromBuffer ? AlignerPlugin_logic_buffer_hm_Prediction_WORD_SLICES_BRANCH : fetch_logic_ctrls_2_down_Prediction_WORD_SLICES_BRANCH);
  assign AlignerPlugin_logic_extractors_1_ctx_hm_Prediction_WORD_SLICES_TAKEN = (AlignerPlugin_logic_buffer_readers_1_lastFromBuffer ? AlignerPlugin_logic_buffer_hm_Prediction_WORD_SLICES_TAKEN : fetch_logic_ctrls_2_down_Prediction_WORD_SLICES_TAKEN);
  assign AlignerPlugin_logic_extractors_1_ctx_hm_Prediction_WORD_JUMP_PC = (AlignerPlugin_logic_buffer_readers_1_lastFromBuffer ? AlignerPlugin_logic_buffer_hm_Prediction_WORD_JUMP_PC : fetch_logic_ctrls_2_down_Prediction_WORD_JUMP_PC);
  assign AlignerPlugin_logic_extractors_1_ctx_hm_Prediction_WORD_JUMPED = (AlignerPlugin_logic_buffer_readers_1_lastFromBuffer ? AlignerPlugin_logic_buffer_hm_Prediction_WORD_JUMPED : fetch_logic_ctrls_2_down_Prediction_WORD_JUMPED);
  assign AlignerPlugin_logic_extractors_1_ctx_hm_Prediction_WORD_JUMP_SLICE = (AlignerPlugin_logic_buffer_readers_1_lastFromBuffer ? AlignerPlugin_logic_buffer_hm_Prediction_WORD_JUMP_SLICE : fetch_logic_ctrls_2_down_Prediction_WORD_JUMP_SLICE);
  assign AlignerPlugin_api_downMoving = toplevel_decode_ctrls_0_up_isMoving;
  assign DispatchPlugin_logic_candidates_0_cancel = (|{(late1_BranchPlugin_logic_flushPort_valid && 1'b1),{(early1_BranchPlugin_logic_flushPort_valid && 1'b1),{(late0_BranchPlugin_logic_flushPort_valid && 1'b1),{(early0_EnvPlugin_logic_flushPort_valid && 1'b1),{(CsrAccessPlugin_logic_flushPort_valid && 1'b1),{(early0_BranchPlugin_logic_flushPort_valid && _zz_DispatchPlugin_logic_candidates_0_cancel),(LsuPlugin_logic_flushPort_valid && _zz_DispatchPlugin_logic_candidates_0_cancel_1)}}}}}});
  assign DispatchPlugin_logic_slotsFeeds_free = (&DispatchPlugin_logic_candidates_0_moving);
  assign DispatchPlugin_logic_slotsFeeds_fit = (_zz_DispatchPlugin_logic_slotsFeeds_fit <= 2'b01);
  assign DispatchPlugin_logic_slotsFeeds_doIt = (DispatchPlugin_logic_slotsFeeds_free && DispatchPlugin_logic_slotsFeeds_fit);
  assign _zz_DispatchPlugin_logic_slots_0_ctx_valid = {(! DispatchPlugin_logic_candidates_2_moving),(! DispatchPlugin_logic_candidates_1_moving)};
  assign _zz_DispatchPlugin_logic_slots_0_ctx_valid_1 = _zz_DispatchPlugin_logic_slots_0_ctx_valid[0];
  always @(*) begin
    _zz_DispatchPlugin_logic_slots_0_ctx_valid_2[0] = (_zz_DispatchPlugin_logic_slots_0_ctx_valid_1 && (! 1'b0));
    _zz_DispatchPlugin_logic_slots_0_ctx_valid_2[1] = (_zz_DispatchPlugin_logic_slots_0_ctx_valid[1] && (! _zz_DispatchPlugin_logic_slots_0_ctx_valid_1));
  end

  assign _zz_DispatchPlugin_logic_slots_0_ctx_valid_3 = _zz_DispatchPlugin_logic_slots_0_ctx_valid_2;
  assign _zz_DispatchPlugin_logic_slots_0_ctx_valid_4 = ((_zz_DispatchPlugin_logic_slots_0_ctx_valid_3[0] ? {{DispatchPlugin_logic_candidates_1_ctx_hm_DispatchPlugin_logic_hcs_3_onRs_1_ENABLES_0,{_zz__zz_DispatchPlugin_logic_slots_0_ctx_valid_4,_zz__zz_DispatchPlugin_logic_slots_0_ctx_valid_4_1}},{DispatchPlugin_logic_candidates_1_ctx_uop,{DispatchPlugin_logic_candidates_1_ctx_laneLayerHits,_zz__zz_DispatchPlugin_logic_slots_0_ctx_valid_4_10}}} : 181'h0) | (_zz_DispatchPlugin_logic_slots_0_ctx_valid_3[1] ? {{DispatchPlugin_logic_candidates_2_ctx_hm_DispatchPlugin_logic_hcs_3_onRs_1_ENABLES_0,{_zz__zz_DispatchPlugin_logic_slots_0_ctx_valid_4_11,_zz__zz_DispatchPlugin_logic_slots_0_ctx_valid_4_12}},{DispatchPlugin_logic_candidates_2_ctx_uop,{DispatchPlugin_logic_candidates_2_ctx_laneLayerHits,_zz__zz_DispatchPlugin_logic_slots_0_ctx_valid_4_21}}} : 181'h0));
  assign _zz_DispatchPlugin_logic_slots_0_ctx_hm_Prediction_ALIGNED_JUMPED = _zz_DispatchPlugin_logic_slots_0_ctx_valid_4[180 : 37];
  assign _zz_DispatchPlugin_logic_slots_0_ctx_hm_GSharePlugin_GSHARE_COUNTER_0 = _zz_DispatchPlugin_logic_slots_0_ctx_hm_Prediction_ALIGNED_JUMPED[48 : 41];
  assign DispatchPlugin_logic_scheduler_eusFree_0 = 2'b11;
  assign DispatchPlugin_logic_scheduler_hartFree_0 = 1'b1;
  assign DispatchPlugin_logic_scheduler_arbiters_0_candHazard = 1'b0;
  assign DispatchPlugin_logic_scheduler_arbiters_0_layersHits = (((DispatchPlugin_logic_candidates_0_ctx_laneLayerHits & (~ DispatchPlugin_logic_candidates_0_rsHazards)) & (~ DispatchPlugin_logic_candidates_0_reservationHazards)) & {DispatchPlugin_logic_scheduler_eusFree_0[0],{DispatchPlugin_logic_scheduler_eusFree_0[1],{DispatchPlugin_logic_scheduler_eusFree_0[0],DispatchPlugin_logic_scheduler_eusFree_0[1]}}});
  assign _zz_DispatchPlugin_logic_scheduler_arbiters_0_layersHits_bools_0 = DispatchPlugin_logic_scheduler_arbiters_0_layersHits;
  assign DispatchPlugin_logic_scheduler_arbiters_0_layersHits_bools_0 = _zz_DispatchPlugin_logic_scheduler_arbiters_0_layersHits_bools_0[0];
  assign DispatchPlugin_logic_scheduler_arbiters_0_layersHits_bools_1 = _zz_DispatchPlugin_logic_scheduler_arbiters_0_layersHits_bools_0[1];
  assign DispatchPlugin_logic_scheduler_arbiters_0_layersHits_bools_2 = _zz_DispatchPlugin_logic_scheduler_arbiters_0_layersHits_bools_0[2];
  assign DispatchPlugin_logic_scheduler_arbiters_0_layersHits_bools_3 = _zz_DispatchPlugin_logic_scheduler_arbiters_0_layersHits_bools_0[3];
  always @(*) begin
    _zz_DispatchPlugin_logic_scheduler_arbiters_0_layerOh[0] = (DispatchPlugin_logic_scheduler_arbiters_0_layersHits_bools_0 && (! 1'b0));
    _zz_DispatchPlugin_logic_scheduler_arbiters_0_layerOh[1] = (DispatchPlugin_logic_scheduler_arbiters_0_layersHits_bools_1 && (! DispatchPlugin_logic_scheduler_arbiters_0_layersHits_bools_0));
    _zz_DispatchPlugin_logic_scheduler_arbiters_0_layerOh[2] = (DispatchPlugin_logic_scheduler_arbiters_0_layersHits_bools_2 && (! DispatchPlugin_logic_scheduler_arbiters_0_layersHits_range_0_to_1));
    _zz_DispatchPlugin_logic_scheduler_arbiters_0_layerOh[3] = (DispatchPlugin_logic_scheduler_arbiters_0_layersHits_bools_3 && (! DispatchPlugin_logic_scheduler_arbiters_0_layersHits_range_0_to_2));
  end

  assign DispatchPlugin_logic_scheduler_arbiters_0_layersHits_range_0_to_1 = (|{DispatchPlugin_logic_scheduler_arbiters_0_layersHits_bools_1,DispatchPlugin_logic_scheduler_arbiters_0_layersHits_bools_0});
  assign DispatchPlugin_logic_scheduler_arbiters_0_layersHits_range_0_to_2 = (|{DispatchPlugin_logic_scheduler_arbiters_0_layersHits_bools_2,{DispatchPlugin_logic_scheduler_arbiters_0_layersHits_bools_1,DispatchPlugin_logic_scheduler_arbiters_0_layersHits_bools_0}});
  assign DispatchPlugin_logic_scheduler_arbiters_0_layerOh = _zz_DispatchPlugin_logic_scheduler_arbiters_0_layerOh;
  assign DispatchPlugin_logic_scheduler_arbiters_0_eusOh = {(|{DispatchPlugin_logic_scheduler_arbiters_0_layerOh[2],DispatchPlugin_logic_scheduler_arbiters_0_layerOh[0]}),(|{DispatchPlugin_logic_scheduler_arbiters_0_layerOh[3],DispatchPlugin_logic_scheduler_arbiters_0_layerOh[1]})};
  assign DispatchPlugin_logic_scheduler_arbiters_0_doIt = (((((DispatchPlugin_logic_candidates_0_ctx_valid && (! DispatchPlugin_logic_candidates_0_flushHazards)) && (! DispatchPlugin_logic_candidates_0_fenceOlderHazards)) && (|DispatchPlugin_logic_scheduler_arbiters_0_layerOh)) && DispatchPlugin_logic_scheduler_hartFree_0[0]) && (! DispatchPlugin_logic_scheduler_arbiters_0_candHazard));
  assign DispatchPlugin_logic_scheduler_eusFree_1 = (DispatchPlugin_logic_scheduler_eusFree_0 & ((! DispatchPlugin_logic_scheduler_arbiters_0_doIt) ? 2'b11 : (~ DispatchPlugin_logic_scheduler_arbiters_0_eusOh)));
  assign DispatchPlugin_logic_scheduler_hartFree_1 = (DispatchPlugin_logic_scheduler_hartFree_0 & (((! DispatchPlugin_logic_candidates_0_ctx_valid) || DispatchPlugin_logic_scheduler_arbiters_0_doIt) ? 1'b1 : (~ 1'b1)));
  assign DispatchPlugin_logic_candidates_0_fire = ((DispatchPlugin_logic_scheduler_arbiters_0_doIt && (! execute_freeze_valid)) && (! DispatchPlugin_api_haltDispatch));
  assign DispatchPlugin_logic_scheduler_arbiters_1_candHazards_0_doWrite = ((DispatchPlugin_logic_candidates_0_ctx_valid && 1'b1) && DispatchPlugin_logic_candidates_0_ctx_hm_RD_ENABLE);
  assign DispatchPlugin_logic_scheduler_arbiters_1_candHazards_0_rfas_0 = ((DispatchPlugin_logic_candidates_1_ctx_hm_RS1_ENABLE && (DispatchPlugin_logic_candidates_0_ctx_hm_RD_PHYS == DispatchPlugin_logic_candidates_1_ctx_hm_RS1_PHYS)) && 1'b1);
  assign DispatchPlugin_logic_scheduler_arbiters_1_candHazards_0_rfas_1 = ((DispatchPlugin_logic_candidates_1_ctx_hm_RS2_ENABLE && (DispatchPlugin_logic_candidates_0_ctx_hm_RD_PHYS == DispatchPlugin_logic_candidates_1_ctx_hm_RS2_PHYS)) && 1'b1);
  assign DispatchPlugin_logic_scheduler_arbiters_1_candHazards_0_rfas_2 = ((DispatchPlugin_logic_candidates_1_ctx_hm_RD_ENABLE && (DispatchPlugin_logic_candidates_0_ctx_hm_RD_PHYS == DispatchPlugin_logic_candidates_1_ctx_hm_RD_PHYS)) && 1'b1);
  assign DispatchPlugin_logic_scheduler_arbiters_1_candHazards_0_hit = (DispatchPlugin_logic_scheduler_arbiters_1_candHazards_0_doWrite && (|{DispatchPlugin_logic_scheduler_arbiters_1_candHazards_0_rfas_2,{DispatchPlugin_logic_scheduler_arbiters_1_candHazards_0_rfas_1,DispatchPlugin_logic_scheduler_arbiters_1_candHazards_0_rfas_0}}));
  assign DispatchPlugin_logic_scheduler_arbiters_1_candHazard = (|DispatchPlugin_logic_scheduler_arbiters_1_candHazards_0_hit);
  assign DispatchPlugin_logic_scheduler_arbiters_1_layersHits = (((DispatchPlugin_logic_candidates_1_ctx_laneLayerHits & (~ DispatchPlugin_logic_candidates_1_rsHazards)) & (~ DispatchPlugin_logic_candidates_1_reservationHazards)) & {DispatchPlugin_logic_scheduler_eusFree_1[0],{DispatchPlugin_logic_scheduler_eusFree_1[1],{DispatchPlugin_logic_scheduler_eusFree_1[0],DispatchPlugin_logic_scheduler_eusFree_1[1]}}});
  assign _zz_DispatchPlugin_logic_scheduler_arbiters_1_layersHits_bools_0 = DispatchPlugin_logic_scheduler_arbiters_1_layersHits;
  assign DispatchPlugin_logic_scheduler_arbiters_1_layersHits_bools_0 = _zz_DispatchPlugin_logic_scheduler_arbiters_1_layersHits_bools_0[0];
  assign DispatchPlugin_logic_scheduler_arbiters_1_layersHits_bools_1 = _zz_DispatchPlugin_logic_scheduler_arbiters_1_layersHits_bools_0[1];
  assign DispatchPlugin_logic_scheduler_arbiters_1_layersHits_bools_2 = _zz_DispatchPlugin_logic_scheduler_arbiters_1_layersHits_bools_0[2];
  assign DispatchPlugin_logic_scheduler_arbiters_1_layersHits_bools_3 = _zz_DispatchPlugin_logic_scheduler_arbiters_1_layersHits_bools_0[3];
  always @(*) begin
    _zz_DispatchPlugin_logic_scheduler_arbiters_1_layerOh[0] = (DispatchPlugin_logic_scheduler_arbiters_1_layersHits_bools_0 && (! 1'b0));
    _zz_DispatchPlugin_logic_scheduler_arbiters_1_layerOh[1] = (DispatchPlugin_logic_scheduler_arbiters_1_layersHits_bools_1 && (! DispatchPlugin_logic_scheduler_arbiters_1_layersHits_bools_0));
    _zz_DispatchPlugin_logic_scheduler_arbiters_1_layerOh[2] = (DispatchPlugin_logic_scheduler_arbiters_1_layersHits_bools_2 && (! DispatchPlugin_logic_scheduler_arbiters_1_layersHits_range_0_to_1));
    _zz_DispatchPlugin_logic_scheduler_arbiters_1_layerOh[3] = (DispatchPlugin_logic_scheduler_arbiters_1_layersHits_bools_3 && (! DispatchPlugin_logic_scheduler_arbiters_1_layersHits_range_0_to_2));
  end

  assign DispatchPlugin_logic_scheduler_arbiters_1_layersHits_range_0_to_1 = (|{DispatchPlugin_logic_scheduler_arbiters_1_layersHits_bools_1,DispatchPlugin_logic_scheduler_arbiters_1_layersHits_bools_0});
  assign DispatchPlugin_logic_scheduler_arbiters_1_layersHits_range_0_to_2 = (|{DispatchPlugin_logic_scheduler_arbiters_1_layersHits_bools_2,{DispatchPlugin_logic_scheduler_arbiters_1_layersHits_bools_1,DispatchPlugin_logic_scheduler_arbiters_1_layersHits_bools_0}});
  assign DispatchPlugin_logic_scheduler_arbiters_1_layerOh = _zz_DispatchPlugin_logic_scheduler_arbiters_1_layerOh;
  assign DispatchPlugin_logic_scheduler_arbiters_1_eusOh = {(|{DispatchPlugin_logic_scheduler_arbiters_1_layerOh[2],DispatchPlugin_logic_scheduler_arbiters_1_layerOh[0]}),(|{DispatchPlugin_logic_scheduler_arbiters_1_layerOh[3],DispatchPlugin_logic_scheduler_arbiters_1_layerOh[1]})};
  assign DispatchPlugin_logic_scheduler_arbiters_1_doIt = (((((DispatchPlugin_logic_candidates_1_ctx_valid && (! DispatchPlugin_logic_candidates_1_flushHazards)) && (! DispatchPlugin_logic_candidates_1_fenceOlderHazards)) && (|DispatchPlugin_logic_scheduler_arbiters_1_layerOh)) && DispatchPlugin_logic_scheduler_hartFree_1[0]) && (! DispatchPlugin_logic_scheduler_arbiters_1_candHazard));
  assign DispatchPlugin_logic_scheduler_eusFree_2 = (DispatchPlugin_logic_scheduler_eusFree_1 & ((! DispatchPlugin_logic_scheduler_arbiters_1_doIt) ? 2'b11 : (~ DispatchPlugin_logic_scheduler_arbiters_1_eusOh)));
  assign DispatchPlugin_logic_scheduler_hartFree_2 = (DispatchPlugin_logic_scheduler_hartFree_1 & (((! DispatchPlugin_logic_candidates_1_ctx_valid) || DispatchPlugin_logic_scheduler_arbiters_1_doIt) ? 1'b1 : (~ 1'b1)));
  assign DispatchPlugin_logic_candidates_1_fire = ((DispatchPlugin_logic_scheduler_arbiters_1_doIt && (! execute_freeze_valid)) && (! DispatchPlugin_api_haltDispatch));
  assign DispatchPlugin_logic_scheduler_arbiters_2_candHazards_0_doWrite = ((DispatchPlugin_logic_candidates_0_ctx_valid && 1'b1) && DispatchPlugin_logic_candidates_0_ctx_hm_RD_ENABLE);
  assign DispatchPlugin_logic_scheduler_arbiters_2_candHazards_0_rfas_0 = ((DispatchPlugin_logic_candidates_2_ctx_hm_RS1_ENABLE && (DispatchPlugin_logic_candidates_0_ctx_hm_RD_PHYS == DispatchPlugin_logic_candidates_2_ctx_hm_RS1_PHYS)) && 1'b1);
  assign DispatchPlugin_logic_scheduler_arbiters_2_candHazards_0_rfas_1 = ((DispatchPlugin_logic_candidates_2_ctx_hm_RS2_ENABLE && (DispatchPlugin_logic_candidates_0_ctx_hm_RD_PHYS == DispatchPlugin_logic_candidates_2_ctx_hm_RS2_PHYS)) && 1'b1);
  assign DispatchPlugin_logic_scheduler_arbiters_2_candHazards_0_rfas_2 = ((DispatchPlugin_logic_candidates_2_ctx_hm_RD_ENABLE && (DispatchPlugin_logic_candidates_0_ctx_hm_RD_PHYS == DispatchPlugin_logic_candidates_2_ctx_hm_RD_PHYS)) && 1'b1);
  assign DispatchPlugin_logic_scheduler_arbiters_2_candHazards_0_hit = (DispatchPlugin_logic_scheduler_arbiters_2_candHazards_0_doWrite && (|{DispatchPlugin_logic_scheduler_arbiters_2_candHazards_0_rfas_2,{DispatchPlugin_logic_scheduler_arbiters_2_candHazards_0_rfas_1,DispatchPlugin_logic_scheduler_arbiters_2_candHazards_0_rfas_0}}));
  assign DispatchPlugin_logic_scheduler_arbiters_2_candHazards_1_doWrite = ((DispatchPlugin_logic_candidates_1_ctx_valid && 1'b1) && DispatchPlugin_logic_candidates_1_ctx_hm_RD_ENABLE);
  assign DispatchPlugin_logic_scheduler_arbiters_2_candHazards_1_rfas_0 = ((DispatchPlugin_logic_candidates_2_ctx_hm_RS1_ENABLE && (DispatchPlugin_logic_candidates_1_ctx_hm_RD_PHYS == DispatchPlugin_logic_candidates_2_ctx_hm_RS1_PHYS)) && 1'b1);
  assign DispatchPlugin_logic_scheduler_arbiters_2_candHazards_1_rfas_1 = ((DispatchPlugin_logic_candidates_2_ctx_hm_RS2_ENABLE && (DispatchPlugin_logic_candidates_1_ctx_hm_RD_PHYS == DispatchPlugin_logic_candidates_2_ctx_hm_RS2_PHYS)) && 1'b1);
  assign DispatchPlugin_logic_scheduler_arbiters_2_candHazards_1_rfas_2 = ((DispatchPlugin_logic_candidates_2_ctx_hm_RD_ENABLE && (DispatchPlugin_logic_candidates_1_ctx_hm_RD_PHYS == DispatchPlugin_logic_candidates_2_ctx_hm_RD_PHYS)) && 1'b1);
  assign DispatchPlugin_logic_scheduler_arbiters_2_candHazards_1_hit = (DispatchPlugin_logic_scheduler_arbiters_2_candHazards_1_doWrite && (|{DispatchPlugin_logic_scheduler_arbiters_2_candHazards_1_rfas_2,{DispatchPlugin_logic_scheduler_arbiters_2_candHazards_1_rfas_1,DispatchPlugin_logic_scheduler_arbiters_2_candHazards_1_rfas_0}}));
  assign DispatchPlugin_logic_scheduler_arbiters_2_candHazard = (|{DispatchPlugin_logic_scheduler_arbiters_2_candHazards_1_hit,DispatchPlugin_logic_scheduler_arbiters_2_candHazards_0_hit});
  assign DispatchPlugin_logic_scheduler_arbiters_2_layersHits = (((DispatchPlugin_logic_candidates_2_ctx_laneLayerHits & (~ DispatchPlugin_logic_candidates_2_rsHazards)) & (~ DispatchPlugin_logic_candidates_2_reservationHazards)) & {DispatchPlugin_logic_scheduler_eusFree_2[0],{DispatchPlugin_logic_scheduler_eusFree_2[1],{DispatchPlugin_logic_scheduler_eusFree_2[0],DispatchPlugin_logic_scheduler_eusFree_2[1]}}});
  assign _zz_DispatchPlugin_logic_scheduler_arbiters_2_layersHits_bools_0 = DispatchPlugin_logic_scheduler_arbiters_2_layersHits;
  assign DispatchPlugin_logic_scheduler_arbiters_2_layersHits_bools_0 = _zz_DispatchPlugin_logic_scheduler_arbiters_2_layersHits_bools_0[0];
  assign DispatchPlugin_logic_scheduler_arbiters_2_layersHits_bools_1 = _zz_DispatchPlugin_logic_scheduler_arbiters_2_layersHits_bools_0[1];
  assign DispatchPlugin_logic_scheduler_arbiters_2_layersHits_bools_2 = _zz_DispatchPlugin_logic_scheduler_arbiters_2_layersHits_bools_0[2];
  assign DispatchPlugin_logic_scheduler_arbiters_2_layersHits_bools_3 = _zz_DispatchPlugin_logic_scheduler_arbiters_2_layersHits_bools_0[3];
  always @(*) begin
    _zz_DispatchPlugin_logic_scheduler_arbiters_2_layerOh[0] = (DispatchPlugin_logic_scheduler_arbiters_2_layersHits_bools_0 && (! 1'b0));
    _zz_DispatchPlugin_logic_scheduler_arbiters_2_layerOh[1] = (DispatchPlugin_logic_scheduler_arbiters_2_layersHits_bools_1 && (! DispatchPlugin_logic_scheduler_arbiters_2_layersHits_bools_0));
    _zz_DispatchPlugin_logic_scheduler_arbiters_2_layerOh[2] = (DispatchPlugin_logic_scheduler_arbiters_2_layersHits_bools_2 && (! DispatchPlugin_logic_scheduler_arbiters_2_layersHits_range_0_to_1));
    _zz_DispatchPlugin_logic_scheduler_arbiters_2_layerOh[3] = (DispatchPlugin_logic_scheduler_arbiters_2_layersHits_bools_3 && (! DispatchPlugin_logic_scheduler_arbiters_2_layersHits_range_0_to_2));
  end

  assign DispatchPlugin_logic_scheduler_arbiters_2_layersHits_range_0_to_1 = (|{DispatchPlugin_logic_scheduler_arbiters_2_layersHits_bools_1,DispatchPlugin_logic_scheduler_arbiters_2_layersHits_bools_0});
  assign DispatchPlugin_logic_scheduler_arbiters_2_layersHits_range_0_to_2 = (|{DispatchPlugin_logic_scheduler_arbiters_2_layersHits_bools_2,{DispatchPlugin_logic_scheduler_arbiters_2_layersHits_bools_1,DispatchPlugin_logic_scheduler_arbiters_2_layersHits_bools_0}});
  assign DispatchPlugin_logic_scheduler_arbiters_2_layerOh = _zz_DispatchPlugin_logic_scheduler_arbiters_2_layerOh;
  assign DispatchPlugin_logic_scheduler_arbiters_2_eusOh = {(|{DispatchPlugin_logic_scheduler_arbiters_2_layerOh[2],DispatchPlugin_logic_scheduler_arbiters_2_layerOh[0]}),(|{DispatchPlugin_logic_scheduler_arbiters_2_layerOh[3],DispatchPlugin_logic_scheduler_arbiters_2_layerOh[1]})};
  assign DispatchPlugin_logic_scheduler_arbiters_2_doIt = (((((DispatchPlugin_logic_candidates_2_ctx_valid && (! DispatchPlugin_logic_candidates_2_flushHazards)) && (! DispatchPlugin_logic_candidates_2_fenceOlderHazards)) && (|DispatchPlugin_logic_scheduler_arbiters_2_layerOh)) && DispatchPlugin_logic_scheduler_hartFree_2[0]) && (! DispatchPlugin_logic_scheduler_arbiters_2_candHazard));
  assign DispatchPlugin_logic_scheduler_eusFree_3 = (DispatchPlugin_logic_scheduler_eusFree_2 & ((! DispatchPlugin_logic_scheduler_arbiters_2_doIt) ? 2'b11 : (~ DispatchPlugin_logic_scheduler_arbiters_2_eusOh)));
  assign DispatchPlugin_logic_scheduler_hartFree_3 = (DispatchPlugin_logic_scheduler_hartFree_2 & (((! DispatchPlugin_logic_candidates_2_ctx_valid) || DispatchPlugin_logic_scheduler_arbiters_2_doIt) ? 1'b1 : (~ 1'b1)));
  assign DispatchPlugin_logic_candidates_2_fire = ((DispatchPlugin_logic_scheduler_arbiters_2_doIt && (! execute_freeze_valid)) && (! DispatchPlugin_api_haltDispatch));
  assign DispatchPlugin_logic_inserter_0_oh = {(DispatchPlugin_logic_scheduler_arbiters_2_doIt && DispatchPlugin_logic_scheduler_arbiters_2_eusOh[0]),{(DispatchPlugin_logic_scheduler_arbiters_1_doIt && DispatchPlugin_logic_scheduler_arbiters_1_eusOh[0]),(DispatchPlugin_logic_scheduler_arbiters_0_doIt && DispatchPlugin_logic_scheduler_arbiters_0_eusOh[0])}};
  assign _zz_toplevel_execute_ctrl0_up_LANE_AGE_lane0 = DispatchPlugin_logic_inserter_0_oh[0];
  assign _zz_toplevel_execute_ctrl0_up_LANE_AGE_lane0_1 = DispatchPlugin_logic_inserter_0_oh[1];
  assign _zz_toplevel_execute_ctrl0_up_LANE_AGE_lane0_2 = DispatchPlugin_logic_inserter_0_oh[2];
  assign DispatchPlugin_logic_inserter_0_trap = _zz_DispatchPlugin_logic_inserter_0_trap[0];
  assign toplevel_execute_ctrl0_up_LANE_SEL_lane0 = (((|DispatchPlugin_logic_inserter_0_oh) && (! _zz_toplevel_execute_ctrl0_up_LANE_SEL_lane0[0])) && (! DispatchPlugin_api_haltDispatch));
  assign toplevel_execute_ctrl0_up_Decode_UOP_lane0 = (((_zz_toplevel_execute_ctrl0_up_LANE_AGE_lane0 ? DispatchPlugin_logic_candidates_0_ctx_uop : 32'h0) | (_zz_toplevel_execute_ctrl0_up_LANE_AGE_lane0_1 ? DispatchPlugin_logic_candidates_1_ctx_uop : 32'h0)) | (_zz_toplevel_execute_ctrl0_up_LANE_AGE_lane0_2 ? DispatchPlugin_logic_candidates_2_ctx_uop : 32'h0));
  assign toplevel_execute_ctrl0_up_Prediction_ALIGNED_JUMPED_lane0 = _zz_toplevel_execute_ctrl0_up_Prediction_ALIGNED_JUMPED_lane0[0];
  assign toplevel_execute_ctrl0_up_Prediction_ALIGNED_JUMPED_PC_lane0 = (((_zz_toplevel_execute_ctrl0_up_LANE_AGE_lane0 ? DispatchPlugin_logic_candidates_0_ctx_hm_Prediction_ALIGNED_JUMPED_PC : 32'h0) | (_zz_toplevel_execute_ctrl0_up_LANE_AGE_lane0_1 ? DispatchPlugin_logic_candidates_1_ctx_hm_Prediction_ALIGNED_JUMPED_PC : 32'h0)) | (_zz_toplevel_execute_ctrl0_up_LANE_AGE_lane0_2 ? DispatchPlugin_logic_candidates_2_ctx_hm_Prediction_ALIGNED_JUMPED_PC : 32'h0));
  assign toplevel_execute_ctrl0_up_Prediction_ALIGNED_SLICES_TAKEN_lane0 = (((_zz_toplevel_execute_ctrl0_up_LANE_AGE_lane0 ? DispatchPlugin_logic_candidates_0_ctx_hm_Prediction_ALIGNED_SLICES_TAKEN : 4'b0000) | (_zz_toplevel_execute_ctrl0_up_LANE_AGE_lane0_1 ? DispatchPlugin_logic_candidates_1_ctx_hm_Prediction_ALIGNED_SLICES_TAKEN : 4'b0000)) | (_zz_toplevel_execute_ctrl0_up_LANE_AGE_lane0_2 ? DispatchPlugin_logic_candidates_2_ctx_hm_Prediction_ALIGNED_SLICES_TAKEN : 4'b0000));
  assign toplevel_execute_ctrl0_up_Prediction_ALIGNED_SLICES_BRANCH_lane0 = (((_zz_toplevel_execute_ctrl0_up_LANE_AGE_lane0 ? DispatchPlugin_logic_candidates_0_ctx_hm_Prediction_ALIGNED_SLICES_BRANCH : 4'b0000) | (_zz_toplevel_execute_ctrl0_up_LANE_AGE_lane0_1 ? DispatchPlugin_logic_candidates_1_ctx_hm_Prediction_ALIGNED_SLICES_BRANCH : 4'b0000)) | (_zz_toplevel_execute_ctrl0_up_LANE_AGE_lane0_2 ? DispatchPlugin_logic_candidates_2_ctx_hm_Prediction_ALIGNED_SLICES_BRANCH : 4'b0000));
  assign _zz_toplevel_execute_ctrl0_up_GSharePlugin_GSHARE_COUNTER_lane0_0 = (((_zz_toplevel_execute_ctrl0_up_LANE_AGE_lane0 ? {DispatchPlugin_logic_candidates_0_ctx_hm_GSharePlugin_GSHARE_COUNTER_3,{_zz__zz_toplevel_execute_ctrl0_up_GSharePlugin_GSHARE_COUNTER_lane0_0,_zz__zz_toplevel_execute_ctrl0_up_GSharePlugin_GSHARE_COUNTER_lane0_0_1}} : 8'h0) | (_zz_toplevel_execute_ctrl0_up_LANE_AGE_lane0_1 ? {DispatchPlugin_logic_candidates_1_ctx_hm_GSharePlugin_GSHARE_COUNTER_3,{_zz__zz_toplevel_execute_ctrl0_up_GSharePlugin_GSHARE_COUNTER_lane0_0_2,_zz__zz_toplevel_execute_ctrl0_up_GSharePlugin_GSHARE_COUNTER_lane0_0_3}} : 8'h0)) | (_zz_toplevel_execute_ctrl0_up_LANE_AGE_lane0_2 ? {DispatchPlugin_logic_candidates_2_ctx_hm_GSharePlugin_GSHARE_COUNTER_3,{DispatchPlugin_logic_candidates_2_ctx_hm_GSharePlugin_GSHARE_COUNTER_2,{_zz__zz_toplevel_execute_ctrl0_up_GSharePlugin_GSHARE_COUNTER_lane0_0_4,_zz__zz_toplevel_execute_ctrl0_up_GSharePlugin_GSHARE_COUNTER_lane0_0_5}}} : 8'h0));
  assign toplevel_execute_ctrl0_up_GSharePlugin_GSHARE_COUNTER_lane0_0 = _zz_toplevel_execute_ctrl0_up_GSharePlugin_GSHARE_COUNTER_lane0_0[1 : 0];
  assign toplevel_execute_ctrl0_up_GSharePlugin_GSHARE_COUNTER_lane0_1 = _zz_toplevel_execute_ctrl0_up_GSharePlugin_GSHARE_COUNTER_lane0_0[3 : 2];
  assign toplevel_execute_ctrl0_up_GSharePlugin_GSHARE_COUNTER_lane0_2 = _zz_toplevel_execute_ctrl0_up_GSharePlugin_GSHARE_COUNTER_lane0_0[5 : 4];
  assign toplevel_execute_ctrl0_up_GSharePlugin_GSHARE_COUNTER_lane0_3 = _zz_toplevel_execute_ctrl0_up_GSharePlugin_GSHARE_COUNTER_lane0_0[7 : 6];
  assign toplevel_execute_ctrl0_up_Prediction_BRANCH_HISTORY_lane0 = (((_zz_toplevel_execute_ctrl0_up_LANE_AGE_lane0 ? DispatchPlugin_logic_candidates_0_ctx_hm_Prediction_BRANCH_HISTORY : 12'h0) | (_zz_toplevel_execute_ctrl0_up_LANE_AGE_lane0_1 ? DispatchPlugin_logic_candidates_1_ctx_hm_Prediction_BRANCH_HISTORY : 12'h0)) | (_zz_toplevel_execute_ctrl0_up_LANE_AGE_lane0_2 ? DispatchPlugin_logic_candidates_2_ctx_hm_Prediction_BRANCH_HISTORY : 12'h0));
  assign toplevel_execute_ctrl0_up_DispatchPlugin_FENCE_OLDER_lane0 = _zz_toplevel_execute_ctrl0_up_DispatchPlugin_FENCE_OLDER_lane0[0];
  always @(*) begin
    toplevel_execute_ctrl0_up_DispatchPlugin_MAY_FLUSH_lane0 = _zz_toplevel_execute_ctrl0_up_DispatchPlugin_MAY_FLUSH_lane0[0];
    if(when_DispatchPlugin_l427) begin
      toplevel_execute_ctrl0_up_DispatchPlugin_MAY_FLUSH_lane0 = 1'b0;
    end
  end

  assign toplevel_execute_ctrl0_up_DispatchPlugin_DONT_FLUSH_lane0 = _zz_toplevel_execute_ctrl0_up_DispatchPlugin_DONT_FLUSH_lane0[0];
  assign toplevel_execute_ctrl0_up_DispatchPlugin_DONT_FLUSH_FROM_LANES_lane0 = _zz_toplevel_execute_ctrl0_up_DispatchPlugin_DONT_FLUSH_FROM_LANES_lane0[0];
  assign toplevel_execute_ctrl0_up_Decode_INSTRUCTION_SLICE_COUNT_lane0 = (((_zz_toplevel_execute_ctrl0_up_LANE_AGE_lane0 ? DispatchPlugin_logic_candidates_0_ctx_hm_Decode_INSTRUCTION_SLICE_COUNT : 1'b0) | (_zz_toplevel_execute_ctrl0_up_LANE_AGE_lane0_1 ? DispatchPlugin_logic_candidates_1_ctx_hm_Decode_INSTRUCTION_SLICE_COUNT : 1'b0)) | (_zz_toplevel_execute_ctrl0_up_LANE_AGE_lane0_2 ? DispatchPlugin_logic_candidates_2_ctx_hm_Decode_INSTRUCTION_SLICE_COUNT : 1'b0));
  assign toplevel_execute_ctrl0_up_DONT_FLUSH_PRECISE_3_lane0 = _zz_toplevel_execute_ctrl0_up_DONT_FLUSH_PRECISE_3_lane0[0];
  assign toplevel_execute_ctrl0_up_DONT_FLUSH_PRECISE_4_lane0 = _zz_toplevel_execute_ctrl0_up_DONT_FLUSH_PRECISE_4_lane0[0];
  assign toplevel_execute_ctrl0_up_PC_lane0 = (((_zz_toplevel_execute_ctrl0_up_LANE_AGE_lane0 ? DispatchPlugin_logic_candidates_0_ctx_hm_PC : 32'h0) | (_zz_toplevel_execute_ctrl0_up_LANE_AGE_lane0_1 ? DispatchPlugin_logic_candidates_1_ctx_hm_PC : 32'h0)) | (_zz_toplevel_execute_ctrl0_up_LANE_AGE_lane0_2 ? DispatchPlugin_logic_candidates_2_ctx_hm_PC : 32'h0));
  assign toplevel_execute_ctrl0_up_TRAP_lane0 = _zz_toplevel_execute_ctrl0_up_TRAP_lane0[0];
  assign toplevel_execute_ctrl0_up_Decode_UOP_ID_lane0 = (((_zz_toplevel_execute_ctrl0_up_LANE_AGE_lane0 ? DispatchPlugin_logic_candidates_0_ctx_hm_Decode_UOP_ID : 16'h0) | (_zz_toplevel_execute_ctrl0_up_LANE_AGE_lane0_1 ? DispatchPlugin_logic_candidates_1_ctx_hm_Decode_UOP_ID : 16'h0)) | (_zz_toplevel_execute_ctrl0_up_LANE_AGE_lane0_2 ? DispatchPlugin_logic_candidates_2_ctx_hm_Decode_UOP_ID : 16'h0));
  assign toplevel_execute_ctrl0_up_RS1_ENABLE_lane0 = _zz_toplevel_execute_ctrl0_up_RS1_ENABLE_lane0[0];
  assign toplevel_execute_ctrl0_up_RS1_PHYS_lane0 = (((_zz_toplevel_execute_ctrl0_up_LANE_AGE_lane0 ? DispatchPlugin_logic_candidates_0_ctx_hm_RS1_PHYS : 5'h0) | (_zz_toplevel_execute_ctrl0_up_LANE_AGE_lane0_1 ? DispatchPlugin_logic_candidates_1_ctx_hm_RS1_PHYS : 5'h0)) | (_zz_toplevel_execute_ctrl0_up_LANE_AGE_lane0_2 ? DispatchPlugin_logic_candidates_2_ctx_hm_RS1_PHYS : 5'h0));
  assign toplevel_execute_ctrl0_up_RS2_ENABLE_lane0 = _zz_toplevel_execute_ctrl0_up_RS2_ENABLE_lane0[0];
  assign toplevel_execute_ctrl0_up_RS2_PHYS_lane0 = (((_zz_toplevel_execute_ctrl0_up_LANE_AGE_lane0 ? DispatchPlugin_logic_candidates_0_ctx_hm_RS2_PHYS : 5'h0) | (_zz_toplevel_execute_ctrl0_up_LANE_AGE_lane0_1 ? DispatchPlugin_logic_candidates_1_ctx_hm_RS2_PHYS : 5'h0)) | (_zz_toplevel_execute_ctrl0_up_LANE_AGE_lane0_2 ? DispatchPlugin_logic_candidates_2_ctx_hm_RS2_PHYS : 5'h0));
  always @(*) begin
    toplevel_execute_ctrl0_up_RD_ENABLE_lane0 = _zz_toplevel_execute_ctrl0_up_RD_ENABLE_lane0[0];
    if(when_DispatchPlugin_l427) begin
      toplevel_execute_ctrl0_up_RD_ENABLE_lane0 = 1'b0;
    end
  end

  assign toplevel_execute_ctrl0_up_RD_PHYS_lane0 = (((_zz_toplevel_execute_ctrl0_up_LANE_AGE_lane0 ? DispatchPlugin_logic_candidates_0_ctx_hm_RD_PHYS : 5'h0) | (_zz_toplevel_execute_ctrl0_up_LANE_AGE_lane0_1 ? DispatchPlugin_logic_candidates_1_ctx_hm_RD_PHYS : 5'h0)) | (_zz_toplevel_execute_ctrl0_up_LANE_AGE_lane0_2 ? DispatchPlugin_logic_candidates_2_ctx_hm_RD_PHYS : 5'h0));
  assign toplevel_execute_ctrl0_up_DispatchPlugin_logic_hcs_0_onRs_0_ENABLES_0_lane0 = _zz_toplevel_execute_ctrl0_up_DispatchPlugin_logic_hcs_0_onRs_0_ENABLES_0_lane0[0];
  assign toplevel_execute_ctrl0_up_DispatchPlugin_logic_hcs_0_onRs_1_ENABLES_0_lane0 = _zz_toplevel_execute_ctrl0_up_DispatchPlugin_logic_hcs_0_onRs_1_ENABLES_0_lane0[0];
  assign toplevel_execute_ctrl0_up_DispatchPlugin_logic_hcs_1_onRs_0_ENABLES_0_lane0 = _zz_toplevel_execute_ctrl0_up_DispatchPlugin_logic_hcs_1_onRs_0_ENABLES_0_lane0[0];
  assign toplevel_execute_ctrl0_up_DispatchPlugin_logic_hcs_1_onRs_1_ENABLES_0_lane0 = _zz_toplevel_execute_ctrl0_up_DispatchPlugin_logic_hcs_1_onRs_1_ENABLES_0_lane0[0];
  assign toplevel_execute_ctrl0_up_DispatchPlugin_logic_hcs_1_onRs_1_ENABLES_1_lane0 = _zz_toplevel_execute_ctrl0_up_DispatchPlugin_logic_hcs_1_onRs_1_ENABLES_1_lane0[0];
  assign toplevel_execute_ctrl0_up_DispatchPlugin_logic_hcs_2_onRs_0_ENABLES_0_lane0 = _zz_toplevel_execute_ctrl0_up_DispatchPlugin_logic_hcs_2_onRs_0_ENABLES_0_lane0[0];
  assign toplevel_execute_ctrl0_up_DispatchPlugin_logic_hcs_2_onRs_1_ENABLES_0_lane0 = _zz_toplevel_execute_ctrl0_up_DispatchPlugin_logic_hcs_2_onRs_1_ENABLES_0_lane0[0];
  assign toplevel_execute_ctrl0_up_DispatchPlugin_logic_hcs_3_onRs_0_ENABLES_0_lane0 = _zz_toplevel_execute_ctrl0_up_DispatchPlugin_logic_hcs_3_onRs_0_ENABLES_0_lane0[0];
  assign toplevel_execute_ctrl0_up_DispatchPlugin_logic_hcs_3_onRs_1_ENABLES_0_lane0 = _zz_toplevel_execute_ctrl0_up_DispatchPlugin_logic_hcs_3_onRs_1_ENABLES_0_lane0[0];
  assign when_DispatchPlugin_l427 = ((! toplevel_execute_ctrl0_up_LANE_SEL_lane0) || DispatchPlugin_logic_inserter_0_trap);
  assign toplevel_execute_ctrl0_up_LANE_AGE_lane0 = (((_zz_toplevel_execute_ctrl0_up_LANE_AGE_lane0 ? DispatchPlugin_logic_candidates_0_age : 1'b0) | (_zz_toplevel_execute_ctrl0_up_LANE_AGE_lane0_1 ? DispatchPlugin_logic_candidates_1_age : 1'b0)) | (_zz_toplevel_execute_ctrl0_up_LANE_AGE_lane0_2 ? DispatchPlugin_logic_candidates_2_age : 1'b0));
  assign toplevel_execute_ctrl0_up_COMPLETED_lane0 = DispatchPlugin_logic_inserter_0_trap;
  assign DispatchPlugin_logic_inserter_0_layerOhUnfiltred = (((_zz_toplevel_execute_ctrl0_up_LANE_AGE_lane0 ? DispatchPlugin_logic_scheduler_arbiters_0_layerOh : 4'b0000) | (_zz_toplevel_execute_ctrl0_up_LANE_AGE_lane0_1 ? DispatchPlugin_logic_scheduler_arbiters_1_layerOh : 4'b0000)) | (_zz_toplevel_execute_ctrl0_up_LANE_AGE_lane0_2 ? DispatchPlugin_logic_scheduler_arbiters_2_layerOh : 4'b0000));
  assign DispatchPlugin_logic_inserter_0_layer_0_0 = 1'b1;
  assign DispatchPlugin_logic_inserter_0_layer_0_1 = DispatchPlugin_logic_inserter_0_layerOhUnfiltred[1];
  assign DispatchPlugin_logic_inserter_0_layer_1_0 = 1'b0;
  assign DispatchPlugin_logic_inserter_0_layer_1_1 = DispatchPlugin_logic_inserter_0_layerOhUnfiltred[3];
  assign _zz_toplevel_execute_ctrl0_up_execute_lane0_LAYER_SEL_lane0 = {DispatchPlugin_logic_inserter_0_layer_1_1,DispatchPlugin_logic_inserter_0_layer_0_1};
  assign toplevel_execute_ctrl0_up_execute_lane0_LAYER_SEL_lane0 = ((_zz_toplevel_execute_ctrl0_up_execute_lane0_LAYER_SEL_lane0[0] ? DispatchPlugin_logic_inserter_0_layer_0_0 : 1'b0) | (_zz_toplevel_execute_ctrl0_up_execute_lane0_LAYER_SEL_lane0[1] ? DispatchPlugin_logic_inserter_0_layer_1_0 : 1'b0));
  assign DispatchPlugin_logic_inserter_1_oh = {(DispatchPlugin_logic_scheduler_arbiters_2_doIt && DispatchPlugin_logic_scheduler_arbiters_2_eusOh[1]),{(DispatchPlugin_logic_scheduler_arbiters_1_doIt && DispatchPlugin_logic_scheduler_arbiters_1_eusOh[1]),(DispatchPlugin_logic_scheduler_arbiters_0_doIt && DispatchPlugin_logic_scheduler_arbiters_0_eusOh[1])}};
  assign _zz_toplevel_execute_ctrl0_up_LANE_AGE_lane1 = DispatchPlugin_logic_inserter_1_oh[0];
  assign _zz_toplevel_execute_ctrl0_up_LANE_AGE_lane1_1 = DispatchPlugin_logic_inserter_1_oh[1];
  assign _zz_toplevel_execute_ctrl0_up_LANE_AGE_lane1_2 = DispatchPlugin_logic_inserter_1_oh[2];
  assign DispatchPlugin_logic_inserter_1_trap = _zz_DispatchPlugin_logic_inserter_1_trap[0];
  assign toplevel_execute_ctrl0_up_LANE_SEL_lane1 = (((|DispatchPlugin_logic_inserter_1_oh) && (! _zz_toplevel_execute_ctrl0_up_LANE_SEL_lane1[0])) && (! DispatchPlugin_api_haltDispatch));
  assign toplevel_execute_ctrl0_up_Decode_UOP_lane1 = (((_zz_toplevel_execute_ctrl0_up_LANE_AGE_lane1 ? DispatchPlugin_logic_candidates_0_ctx_uop : 32'h0) | (_zz_toplevel_execute_ctrl0_up_LANE_AGE_lane1_1 ? DispatchPlugin_logic_candidates_1_ctx_uop : 32'h0)) | (_zz_toplevel_execute_ctrl0_up_LANE_AGE_lane1_2 ? DispatchPlugin_logic_candidates_2_ctx_uop : 32'h0));
  assign toplevel_execute_ctrl0_up_Prediction_ALIGNED_JUMPED_lane1 = _zz_toplevel_execute_ctrl0_up_Prediction_ALIGNED_JUMPED_lane1[0];
  assign toplevel_execute_ctrl0_up_Prediction_ALIGNED_JUMPED_PC_lane1 = (((_zz_toplevel_execute_ctrl0_up_LANE_AGE_lane1 ? DispatchPlugin_logic_candidates_0_ctx_hm_Prediction_ALIGNED_JUMPED_PC : 32'h0) | (_zz_toplevel_execute_ctrl0_up_LANE_AGE_lane1_1 ? DispatchPlugin_logic_candidates_1_ctx_hm_Prediction_ALIGNED_JUMPED_PC : 32'h0)) | (_zz_toplevel_execute_ctrl0_up_LANE_AGE_lane1_2 ? DispatchPlugin_logic_candidates_2_ctx_hm_Prediction_ALIGNED_JUMPED_PC : 32'h0));
  assign toplevel_execute_ctrl0_up_Prediction_ALIGNED_SLICES_TAKEN_lane1 = (((_zz_toplevel_execute_ctrl0_up_LANE_AGE_lane1 ? DispatchPlugin_logic_candidates_0_ctx_hm_Prediction_ALIGNED_SLICES_TAKEN : 4'b0000) | (_zz_toplevel_execute_ctrl0_up_LANE_AGE_lane1_1 ? DispatchPlugin_logic_candidates_1_ctx_hm_Prediction_ALIGNED_SLICES_TAKEN : 4'b0000)) | (_zz_toplevel_execute_ctrl0_up_LANE_AGE_lane1_2 ? DispatchPlugin_logic_candidates_2_ctx_hm_Prediction_ALIGNED_SLICES_TAKEN : 4'b0000));
  assign toplevel_execute_ctrl0_up_Prediction_ALIGNED_SLICES_BRANCH_lane1 = (((_zz_toplevel_execute_ctrl0_up_LANE_AGE_lane1 ? DispatchPlugin_logic_candidates_0_ctx_hm_Prediction_ALIGNED_SLICES_BRANCH : 4'b0000) | (_zz_toplevel_execute_ctrl0_up_LANE_AGE_lane1_1 ? DispatchPlugin_logic_candidates_1_ctx_hm_Prediction_ALIGNED_SLICES_BRANCH : 4'b0000)) | (_zz_toplevel_execute_ctrl0_up_LANE_AGE_lane1_2 ? DispatchPlugin_logic_candidates_2_ctx_hm_Prediction_ALIGNED_SLICES_BRANCH : 4'b0000));
  assign _zz_toplevel_execute_ctrl0_up_GSharePlugin_GSHARE_COUNTER_lane1_0 = (((_zz_toplevel_execute_ctrl0_up_LANE_AGE_lane1 ? {DispatchPlugin_logic_candidates_0_ctx_hm_GSharePlugin_GSHARE_COUNTER_3,{DispatchPlugin_logic_candidates_0_ctx_hm_GSharePlugin_GSHARE_COUNTER_2,{_zz__zz_toplevel_execute_ctrl0_up_GSharePlugin_GSHARE_COUNTER_lane1_0,_zz__zz_toplevel_execute_ctrl0_up_GSharePlugin_GSHARE_COUNTER_lane1_0_1}}} : 8'h0) | (_zz_toplevel_execute_ctrl0_up_LANE_AGE_lane1_1 ? {DispatchPlugin_logic_candidates_1_ctx_hm_GSharePlugin_GSHARE_COUNTER_3,{DispatchPlugin_logic_candidates_1_ctx_hm_GSharePlugin_GSHARE_COUNTER_2,{_zz__zz_toplevel_execute_ctrl0_up_GSharePlugin_GSHARE_COUNTER_lane1_0_2,_zz__zz_toplevel_execute_ctrl0_up_GSharePlugin_GSHARE_COUNTER_lane1_0_3}}} : 8'h0)) | (_zz_toplevel_execute_ctrl0_up_LANE_AGE_lane1_2 ? {DispatchPlugin_logic_candidates_2_ctx_hm_GSharePlugin_GSHARE_COUNTER_3,{DispatchPlugin_logic_candidates_2_ctx_hm_GSharePlugin_GSHARE_COUNTER_2,{DispatchPlugin_logic_candidates_2_ctx_hm_GSharePlugin_GSHARE_COUNTER_1,DispatchPlugin_logic_candidates_2_ctx_hm_GSharePlugin_GSHARE_COUNTER_0}}} : 8'h0));
  assign toplevel_execute_ctrl0_up_GSharePlugin_GSHARE_COUNTER_lane1_0 = _zz_toplevel_execute_ctrl0_up_GSharePlugin_GSHARE_COUNTER_lane1_0[1 : 0];
  assign toplevel_execute_ctrl0_up_GSharePlugin_GSHARE_COUNTER_lane1_1 = _zz_toplevel_execute_ctrl0_up_GSharePlugin_GSHARE_COUNTER_lane1_0[3 : 2];
  assign toplevel_execute_ctrl0_up_GSharePlugin_GSHARE_COUNTER_lane1_2 = _zz_toplevel_execute_ctrl0_up_GSharePlugin_GSHARE_COUNTER_lane1_0[5 : 4];
  assign toplevel_execute_ctrl0_up_GSharePlugin_GSHARE_COUNTER_lane1_3 = _zz_toplevel_execute_ctrl0_up_GSharePlugin_GSHARE_COUNTER_lane1_0[7 : 6];
  assign toplevel_execute_ctrl0_up_Prediction_BRANCH_HISTORY_lane1 = (((_zz_toplevel_execute_ctrl0_up_LANE_AGE_lane1 ? DispatchPlugin_logic_candidates_0_ctx_hm_Prediction_BRANCH_HISTORY : 12'h0) | (_zz_toplevel_execute_ctrl0_up_LANE_AGE_lane1_1 ? DispatchPlugin_logic_candidates_1_ctx_hm_Prediction_BRANCH_HISTORY : 12'h0)) | (_zz_toplevel_execute_ctrl0_up_LANE_AGE_lane1_2 ? DispatchPlugin_logic_candidates_2_ctx_hm_Prediction_BRANCH_HISTORY : 12'h0));
  assign toplevel_execute_ctrl0_up_DispatchPlugin_FENCE_OLDER_lane1 = _zz_toplevel_execute_ctrl0_up_DispatchPlugin_FENCE_OLDER_lane1[0];
  always @(*) begin
    toplevel_execute_ctrl0_up_DispatchPlugin_MAY_FLUSH_lane1 = _zz_toplevel_execute_ctrl0_up_DispatchPlugin_MAY_FLUSH_lane1[0];
    if(when_DispatchPlugin_l427_1) begin
      toplevel_execute_ctrl0_up_DispatchPlugin_MAY_FLUSH_lane1 = 1'b0;
    end
  end

  assign toplevel_execute_ctrl0_up_DispatchPlugin_DONT_FLUSH_lane1 = _zz_toplevel_execute_ctrl0_up_DispatchPlugin_DONT_FLUSH_lane1[0];
  assign toplevel_execute_ctrl0_up_DispatchPlugin_DONT_FLUSH_FROM_LANES_lane1 = _zz_toplevel_execute_ctrl0_up_DispatchPlugin_DONT_FLUSH_FROM_LANES_lane1[0];
  assign toplevel_execute_ctrl0_up_Decode_INSTRUCTION_SLICE_COUNT_lane1 = (((_zz_toplevel_execute_ctrl0_up_LANE_AGE_lane1 ? DispatchPlugin_logic_candidates_0_ctx_hm_Decode_INSTRUCTION_SLICE_COUNT : 1'b0) | (_zz_toplevel_execute_ctrl0_up_LANE_AGE_lane1_1 ? DispatchPlugin_logic_candidates_1_ctx_hm_Decode_INSTRUCTION_SLICE_COUNT : 1'b0)) | (_zz_toplevel_execute_ctrl0_up_LANE_AGE_lane1_2 ? DispatchPlugin_logic_candidates_2_ctx_hm_Decode_INSTRUCTION_SLICE_COUNT : 1'b0));
  assign toplevel_execute_ctrl0_up_DONT_FLUSH_PRECISE_3_lane1 = _zz_toplevel_execute_ctrl0_up_DONT_FLUSH_PRECISE_3_lane1[0];
  assign toplevel_execute_ctrl0_up_DONT_FLUSH_PRECISE_4_lane1 = _zz_toplevel_execute_ctrl0_up_DONT_FLUSH_PRECISE_4_lane1[0];
  assign toplevel_execute_ctrl0_up_PC_lane1 = (((_zz_toplevel_execute_ctrl0_up_LANE_AGE_lane1 ? DispatchPlugin_logic_candidates_0_ctx_hm_PC : 32'h0) | (_zz_toplevel_execute_ctrl0_up_LANE_AGE_lane1_1 ? DispatchPlugin_logic_candidates_1_ctx_hm_PC : 32'h0)) | (_zz_toplevel_execute_ctrl0_up_LANE_AGE_lane1_2 ? DispatchPlugin_logic_candidates_2_ctx_hm_PC : 32'h0));
  assign toplevel_execute_ctrl0_up_TRAP_lane1 = _zz_toplevel_execute_ctrl0_up_TRAP_lane1[0];
  assign toplevel_execute_ctrl0_up_Decode_UOP_ID_lane1 = (((_zz_toplevel_execute_ctrl0_up_LANE_AGE_lane1 ? DispatchPlugin_logic_candidates_0_ctx_hm_Decode_UOP_ID : 16'h0) | (_zz_toplevel_execute_ctrl0_up_LANE_AGE_lane1_1 ? DispatchPlugin_logic_candidates_1_ctx_hm_Decode_UOP_ID : 16'h0)) | (_zz_toplevel_execute_ctrl0_up_LANE_AGE_lane1_2 ? DispatchPlugin_logic_candidates_2_ctx_hm_Decode_UOP_ID : 16'h0));
  assign toplevel_execute_ctrl0_up_RS1_ENABLE_lane1 = _zz_toplevel_execute_ctrl0_up_RS1_ENABLE_lane1[0];
  assign toplevel_execute_ctrl0_up_RS1_PHYS_lane1 = (((_zz_toplevel_execute_ctrl0_up_LANE_AGE_lane1 ? DispatchPlugin_logic_candidates_0_ctx_hm_RS1_PHYS : 5'h0) | (_zz_toplevel_execute_ctrl0_up_LANE_AGE_lane1_1 ? DispatchPlugin_logic_candidates_1_ctx_hm_RS1_PHYS : 5'h0)) | (_zz_toplevel_execute_ctrl0_up_LANE_AGE_lane1_2 ? DispatchPlugin_logic_candidates_2_ctx_hm_RS1_PHYS : 5'h0));
  assign toplevel_execute_ctrl0_up_RS2_ENABLE_lane1 = _zz_toplevel_execute_ctrl0_up_RS2_ENABLE_lane1[0];
  assign toplevel_execute_ctrl0_up_RS2_PHYS_lane1 = (((_zz_toplevel_execute_ctrl0_up_LANE_AGE_lane1 ? DispatchPlugin_logic_candidates_0_ctx_hm_RS2_PHYS : 5'h0) | (_zz_toplevel_execute_ctrl0_up_LANE_AGE_lane1_1 ? DispatchPlugin_logic_candidates_1_ctx_hm_RS2_PHYS : 5'h0)) | (_zz_toplevel_execute_ctrl0_up_LANE_AGE_lane1_2 ? DispatchPlugin_logic_candidates_2_ctx_hm_RS2_PHYS : 5'h0));
  always @(*) begin
    toplevel_execute_ctrl0_up_RD_ENABLE_lane1 = _zz_toplevel_execute_ctrl0_up_RD_ENABLE_lane1[0];
    if(when_DispatchPlugin_l427_1) begin
      toplevel_execute_ctrl0_up_RD_ENABLE_lane1 = 1'b0;
    end
  end

  assign toplevel_execute_ctrl0_up_RD_PHYS_lane1 = (((_zz_toplevel_execute_ctrl0_up_LANE_AGE_lane1 ? DispatchPlugin_logic_candidates_0_ctx_hm_RD_PHYS : 5'h0) | (_zz_toplevel_execute_ctrl0_up_LANE_AGE_lane1_1 ? DispatchPlugin_logic_candidates_1_ctx_hm_RD_PHYS : 5'h0)) | (_zz_toplevel_execute_ctrl0_up_LANE_AGE_lane1_2 ? DispatchPlugin_logic_candidates_2_ctx_hm_RD_PHYS : 5'h0));
  assign toplevel_execute_ctrl0_up_DispatchPlugin_logic_hcs_0_onRs_0_ENABLES_0_lane1 = _zz_toplevel_execute_ctrl0_up_DispatchPlugin_logic_hcs_0_onRs_0_ENABLES_0_lane1[0];
  assign toplevel_execute_ctrl0_up_DispatchPlugin_logic_hcs_0_onRs_1_ENABLES_0_lane1 = _zz_toplevel_execute_ctrl0_up_DispatchPlugin_logic_hcs_0_onRs_1_ENABLES_0_lane1[0];
  assign toplevel_execute_ctrl0_up_DispatchPlugin_logic_hcs_1_onRs_0_ENABLES_0_lane1 = _zz_toplevel_execute_ctrl0_up_DispatchPlugin_logic_hcs_1_onRs_0_ENABLES_0_lane1[0];
  assign toplevel_execute_ctrl0_up_DispatchPlugin_logic_hcs_1_onRs_1_ENABLES_0_lane1 = _zz_toplevel_execute_ctrl0_up_DispatchPlugin_logic_hcs_1_onRs_1_ENABLES_0_lane1[0];
  assign toplevel_execute_ctrl0_up_DispatchPlugin_logic_hcs_1_onRs_1_ENABLES_1_lane1 = _zz_toplevel_execute_ctrl0_up_DispatchPlugin_logic_hcs_1_onRs_1_ENABLES_1_lane1[0];
  assign toplevel_execute_ctrl0_up_DispatchPlugin_logic_hcs_2_onRs_0_ENABLES_0_lane1 = _zz_toplevel_execute_ctrl0_up_DispatchPlugin_logic_hcs_2_onRs_0_ENABLES_0_lane1[0];
  assign toplevel_execute_ctrl0_up_DispatchPlugin_logic_hcs_2_onRs_1_ENABLES_0_lane1 = _zz_toplevel_execute_ctrl0_up_DispatchPlugin_logic_hcs_2_onRs_1_ENABLES_0_lane1[0];
  assign toplevel_execute_ctrl0_up_DispatchPlugin_logic_hcs_3_onRs_0_ENABLES_0_lane1 = _zz_toplevel_execute_ctrl0_up_DispatchPlugin_logic_hcs_3_onRs_0_ENABLES_0_lane1[0];
  assign toplevel_execute_ctrl0_up_DispatchPlugin_logic_hcs_3_onRs_1_ENABLES_0_lane1 = _zz_toplevel_execute_ctrl0_up_DispatchPlugin_logic_hcs_3_onRs_1_ENABLES_0_lane1[0];
  assign when_DispatchPlugin_l427_1 = ((! toplevel_execute_ctrl0_up_LANE_SEL_lane1) || DispatchPlugin_logic_inserter_1_trap);
  assign toplevel_execute_ctrl0_up_LANE_AGE_lane1 = (((_zz_toplevel_execute_ctrl0_up_LANE_AGE_lane1 ? DispatchPlugin_logic_candidates_0_age : 1'b0) | (_zz_toplevel_execute_ctrl0_up_LANE_AGE_lane1_1 ? DispatchPlugin_logic_candidates_1_age : 1'b0)) | (_zz_toplevel_execute_ctrl0_up_LANE_AGE_lane1_2 ? DispatchPlugin_logic_candidates_2_age : 1'b0));
  assign toplevel_execute_ctrl0_up_COMPLETED_lane1 = DispatchPlugin_logic_inserter_1_trap;
  assign DispatchPlugin_logic_inserter_1_layerOhUnfiltred = (((_zz_toplevel_execute_ctrl0_up_LANE_AGE_lane1 ? DispatchPlugin_logic_scheduler_arbiters_0_layerOh : 4'b0000) | (_zz_toplevel_execute_ctrl0_up_LANE_AGE_lane1_1 ? DispatchPlugin_logic_scheduler_arbiters_1_layerOh : 4'b0000)) | (_zz_toplevel_execute_ctrl0_up_LANE_AGE_lane1_2 ? DispatchPlugin_logic_scheduler_arbiters_2_layerOh : 4'b0000));
  assign DispatchPlugin_logic_inserter_1_layer_0_0 = 1'b1;
  assign DispatchPlugin_logic_inserter_1_layer_0_1 = DispatchPlugin_logic_inserter_1_layerOhUnfiltred[0];
  assign DispatchPlugin_logic_inserter_1_layer_1_0 = 1'b0;
  assign DispatchPlugin_logic_inserter_1_layer_1_1 = DispatchPlugin_logic_inserter_1_layerOhUnfiltred[2];
  assign _zz_toplevel_execute_ctrl0_up_execute_lane1_LAYER_SEL_lane1 = {DispatchPlugin_logic_inserter_1_layer_1_1,DispatchPlugin_logic_inserter_1_layer_0_1};
  assign toplevel_execute_ctrl0_up_execute_lane1_LAYER_SEL_lane1 = ((_zz_toplevel_execute_ctrl0_up_execute_lane1_LAYER_SEL_lane1[0] ? DispatchPlugin_logic_inserter_1_layer_0_0 : 1'b0) | (_zz_toplevel_execute_ctrl0_up_execute_lane1_LAYER_SEL_lane1[1] ? DispatchPlugin_logic_inserter_1_layer_1_0 : 1'b0));
  always @(*) begin
    TrapPlugin_logic_harts_0_crsPorts_read_valid = 1'b0;
    case(TrapPlugin_logic_harts_0_trap_fsm_stateReg)
      TrapPlugin_logic_harts_0_trap_fsm_enumDef_RUNNING : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_enumDef_PROCESS_1 : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_enumDef_TRAP_EPC : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_enumDef_TRAP_TVAL : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_enumDef_TRAP_TVEC : begin
        TrapPlugin_logic_harts_0_crsPorts_read_valid = 1'b1;
      end
      TrapPlugin_logic_harts_0_trap_fsm_enumDef_TRAP_APPLY : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_enumDef_XRET_EPC : begin
        TrapPlugin_logic_harts_0_crsPorts_read_valid = 1'b1;
      end
      TrapPlugin_logic_harts_0_trap_fsm_enumDef_XRET_APPLY : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_enumDef_ATS_RSP : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_enumDef_JUMP : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_enumDef_LSU_FLUSH : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_enumDef_FETCH_FLUSH : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    TrapPlugin_logic_harts_0_crsPorts_read_address = 3'bxxx;
    case(TrapPlugin_logic_harts_0_trap_fsm_stateReg)
      TrapPlugin_logic_harts_0_trap_fsm_enumDef_RUNNING : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_enumDef_PROCESS_1 : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_enumDef_TRAP_EPC : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_enumDef_TRAP_TVAL : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_enumDef_TRAP_TVEC : begin
        TrapPlugin_logic_harts_0_crsPorts_read_address = _zz_TrapPlugin_logic_harts_0_crsPorts_read_address;
      end
      TrapPlugin_logic_harts_0_trap_fsm_enumDef_TRAP_APPLY : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_enumDef_XRET_EPC : begin
        TrapPlugin_logic_harts_0_crsPorts_read_address = _zz_TrapPlugin_logic_harts_0_crsPorts_read_address_1;
      end
      TrapPlugin_logic_harts_0_trap_fsm_enumDef_XRET_APPLY : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_enumDef_ATS_RSP : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_enumDef_JUMP : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_enumDef_LSU_FLUSH : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_enumDef_FETCH_FLUSH : begin
      end
      default : begin
      end
    endcase
  end

  assign decode_logic_flushes_0_onLanes_0_doIt = (|{(DecoderPlugin_logic_laneLogic_1_flushPort_valid && 1'b1),{(DecoderPlugin_logic_laneLogic_0_flushPort_valid && 1'b1),{(late1_BranchPlugin_logic_flushPort_valid && 1'b1),{(early1_BranchPlugin_logic_flushPort_valid && 1'b1),{(late0_BranchPlugin_logic_flushPort_valid && 1'b1),{(early0_EnvPlugin_logic_flushPort_valid && _zz_decode_logic_flushes_0_onLanes_0_doIt),{_zz_decode_logic_flushes_0_onLanes_0_doIt_1,{_zz_decode_logic_flushes_0_onLanes_0_doIt_2,_zz_decode_logic_flushes_0_onLanes_0_doIt_3}}}}}}}});
  assign toplevel_decode_ctrls_0_lane0_downIsCancel = 1'b0;
  assign toplevel_decode_ctrls_0_lane0_upIsCancel = decode_logic_flushes_0_onLanes_0_doIt;
  assign decode_logic_flushes_0_onLanes_1_doIt = (|{(DecoderPlugin_logic_laneLogic_1_flushPort_valid && 1'b1),{(DecoderPlugin_logic_laneLogic_0_flushPort_valid && 1'b1),{(late1_BranchPlugin_logic_flushPort_valid && 1'b1),{(early1_BranchPlugin_logic_flushPort_valid && 1'b1),{(late0_BranchPlugin_logic_flushPort_valid && 1'b1),{(early0_EnvPlugin_logic_flushPort_valid && _zz_decode_logic_flushes_0_onLanes_1_doIt),{_zz_decode_logic_flushes_0_onLanes_1_doIt_1,{_zz_decode_logic_flushes_0_onLanes_1_doIt_2,_zz_decode_logic_flushes_0_onLanes_1_doIt_3}}}}}}}});
  assign toplevel_decode_ctrls_0_lane1_downIsCancel = 1'b0;
  assign toplevel_decode_ctrls_0_lane1_upIsCancel = decode_logic_flushes_0_onLanes_1_doIt;
  assign decode_logic_flushes_1_onLanes_0_doIt = (|{((DecoderPlugin_logic_laneLogic_1_flushPort_valid && 1'b1) && ((DecoderPlugin_logic_laneLogic_1_flushPort_payload_laneAge < _zz_decode_logic_flushes_1_onLanes_0_doIt) || (_zz_decode_logic_flushes_1_onLanes_0_doIt_1 && DecoderPlugin_logic_laneLogic_1_flushPort_payload_self))),{((DecoderPlugin_logic_laneLogic_0_flushPort_valid && _zz_decode_logic_flushes_1_onLanes_0_doIt_2) && (_zz_decode_logic_flushes_1_onLanes_0_doIt_3 || _zz_decode_logic_flushes_1_onLanes_0_doIt_4)),{(late1_BranchPlugin_logic_flushPort_valid && _zz_decode_logic_flushes_1_onLanes_0_doIt_5),{_zz_decode_logic_flushes_1_onLanes_0_doIt_6,{_zz_decode_logic_flushes_1_onLanes_0_doIt_7,_zz_decode_logic_flushes_1_onLanes_0_doIt_8}}}}});
  assign toplevel_decode_ctrls_1_lane0_downIsCancel = 1'b0;
  assign toplevel_decode_ctrls_1_lane0_upIsCancel = decode_logic_flushes_1_onLanes_0_doIt;
  assign _zz_decode_logic_flushes_1_onLanes_1_doIt = 1'b1;
  assign decode_logic_flushes_1_onLanes_1_doIt = (|{((DecoderPlugin_logic_laneLogic_1_flushPort_valid && 1'b1) && ((DecoderPlugin_logic_laneLogic_1_flushPort_payload_laneAge < _zz_decode_logic_flushes_1_onLanes_1_doIt) || ((DecoderPlugin_logic_laneLogic_1_flushPort_payload_laneAge == _zz_decode_logic_flushes_1_onLanes_1_doIt) && DecoderPlugin_logic_laneLogic_1_flushPort_payload_self))),{((DecoderPlugin_logic_laneLogic_0_flushPort_valid && 1'b1) && ((DecoderPlugin_logic_laneLogic_0_flushPort_payload_laneAge < _zz_decode_logic_flushes_1_onLanes_1_doIt) || (_zz_decode_logic_flushes_1_onLanes_1_doIt_1 && DecoderPlugin_logic_laneLogic_0_flushPort_payload_self))),{(late1_BranchPlugin_logic_flushPort_valid && 1'b1),{(early1_BranchPlugin_logic_flushPort_valid && _zz_decode_logic_flushes_1_onLanes_1_doIt_2),{_zz_decode_logic_flushes_1_onLanes_1_doIt_3,{_zz_decode_logic_flushes_1_onLanes_1_doIt_4,_zz_decode_logic_flushes_1_onLanes_1_doIt_5}}}}}});
  assign toplevel_decode_ctrls_1_lane1_downIsCancel = 1'b0;
  assign toplevel_decode_ctrls_1_lane1_upIsCancel = decode_logic_flushes_1_onLanes_1_doIt;
  assign decode_logic_trapPending[0] = (|{((toplevel_decode_ctrls_1_up_LANE_SEL_1 && 1'b1) && toplevel_decode_ctrls_1_down_TRAP_1),{((toplevel_decode_ctrls_1_up_LANE_SEL_0 && 1'b1) && toplevel_decode_ctrls_1_down_TRAP_0),{((toplevel_decode_ctrls_0_up_LANE_SEL_1 && 1'b1) && toplevel_decode_ctrls_0_down_TRAP_1),((toplevel_decode_ctrls_0_up_LANE_SEL_0 && 1'b1) && toplevel_decode_ctrls_0_down_TRAP_0)}}});
  assign toplevel_execute_lane1_bypasser_integer_RS1_port_valid = (! execute_freeze_valid);
  assign toplevel_execute_lane1_bypasser_integer_RS1_port_address = toplevel_execute_ctrl0_down_RS1_PHYS_lane1;
  always @(*) begin
    LsuL1Plugin_logic_banksWrite_address = 9'bxxxxxxxxx;
    LsuL1Plugin_logic_banksWrite_address = {LsuL1Plugin_logic_refill_read_rspAddress[11 : 6],LsuL1Plugin_logic_refill_read_wordIndex};
    if(LsuL1Plugin_logic_ls_ctrl_bankWriteReservation_win) begin
      LsuL1Plugin_logic_banksWrite_address = toplevel_execute_ctrl4_down_LsuL1_PHYSICAL_ADDRESS_lane0[11 : 3];
    end
    if(LsuL1Plugin_logic_initializerMem_busy) begin
      LsuL1Plugin_logic_banksWrite_address = LsuL1Plugin_logic_initializerMem_counter[8:0];
    end
  end

  always @(*) begin
    LsuL1Plugin_logic_banksWrite_writeData = 64'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
    LsuL1Plugin_logic_banksWrite_writeData = LsuL1Plugin_logic_bus_read_rsp_payload_data;
    if(LsuL1Plugin_logic_ls_ctrl_bankWriteReservation_win) begin
      LsuL1Plugin_logic_banksWrite_writeData[31 : 0] = toplevel_execute_ctrl4_down_LsuL1_WRITE_DATA_lane0;
      LsuL1Plugin_logic_banksWrite_writeData[63 : 32] = toplevel_execute_ctrl4_down_LsuL1_WRITE_DATA_lane0;
    end
    if(LsuL1Plugin_logic_initializerMem_busy) begin
      LsuL1Plugin_logic_banksWrite_writeData = 64'h0;
    end
  end

  always @(*) begin
    LsuL1Plugin_logic_banksWrite_writeMask = 8'bxxxxxxxx;
    LsuL1Plugin_logic_banksWrite_writeMask = 8'hff;
    if(LsuL1Plugin_logic_ls_ctrl_bankWriteReservation_win) begin
      LsuL1Plugin_logic_banksWrite_writeMask = 8'h0;
      if(_zz_39[0]) begin
        LsuL1Plugin_logic_banksWrite_writeMask[3 : 0] = toplevel_execute_ctrl4_down_LsuL1_MASK_lane0;
      end
      if(_zz_39[1]) begin
        LsuL1Plugin_logic_banksWrite_writeMask[7 : 4] = toplevel_execute_ctrl4_down_LsuL1_MASK_lane0;
      end
    end
    if(LsuL1Plugin_logic_ls_ctrl_preventSideEffects) begin
      if(LsuL1Plugin_logic_ls_ctrl_bankWriteReservation_win) begin
        LsuL1Plugin_logic_banksWrite_writeMask = 8'h0;
      end
    end
    if(LsuL1Plugin_logic_initializerMem_busy) begin
      LsuL1Plugin_logic_banksWrite_writeMask = 8'hff;
    end
  end

  always @(*) begin
    LsuL1Plugin_logic_waysWrite_mask = 2'b00;
    if(LsuL1Plugin_logic_bus_read_rsp_valid) begin
      if(when_LsuL1Plugin_l446) begin
        LsuL1Plugin_logic_waysWrite_mask[LsuL1Plugin_logic_refill_read_way] = 1'b1;
      end
    end
    if(LsuL1Plugin_logic_ls_ctrl_doFlush) begin
      LsuL1Plugin_logic_waysWrite_mask = LsuL1Plugin_logic_ls_ctrl_needFlushOh;
    end
    if(LsuL1Plugin_logic_ls_ctrl_preventSideEffects) begin
      if(LsuL1Plugin_logic_ls_ctrl_wayWriteReservation_win) begin
        LsuL1Plugin_logic_waysWrite_mask = 2'b00;
      end
    end
    if(when_LsuL1Plugin_l1160) begin
      LsuL1Plugin_logic_waysWrite_mask = 2'b11;
    end
  end

  always @(*) begin
    LsuL1Plugin_logic_waysWrite_address = 6'bxxxxxx;
    if(LsuL1Plugin_logic_bus_read_rsp_valid) begin
      if(when_LsuL1Plugin_l446) begin
        LsuL1Plugin_logic_waysWrite_address = LsuL1Plugin_logic_refill_read_rspAddress[11 : 6];
      end
    end
    if(LsuL1Plugin_logic_ls_ctrl_doFlush) begin
      LsuL1Plugin_logic_waysWrite_address = toplevel_execute_ctrl4_down_LsuL1_MIXED_ADDRESS_lane0[11 : 6];
    end
    if(when_LsuL1Plugin_l1160) begin
      LsuL1Plugin_logic_waysWrite_address = LsuL1Plugin_logic_initializer_counter[5:0];
    end
  end

  always @(*) begin
    LsuL1Plugin_logic_waysWrite_tag_loaded = 1'bx;
    if(LsuL1Plugin_logic_bus_read_rsp_valid) begin
      if(when_LsuL1Plugin_l446) begin
        LsuL1Plugin_logic_waysWrite_tag_loaded = 1'b1;
      end
    end
    if(LsuL1Plugin_logic_ls_ctrl_doFlush) begin
      LsuL1Plugin_logic_waysWrite_tag_loaded = 1'b1;
    end
    if(when_LsuL1Plugin_l1160) begin
      LsuL1Plugin_logic_waysWrite_tag_loaded = 1'b0;
    end
  end

  always @(*) begin
    LsuL1Plugin_logic_waysWrite_tag_address = 20'bxxxxxxxxxxxxxxxxxxxx;
    if(LsuL1Plugin_logic_bus_read_rsp_valid) begin
      if(when_LsuL1Plugin_l446) begin
        LsuL1Plugin_logic_waysWrite_tag_address = LsuL1Plugin_logic_refill_read_rspAddress[31 : 12];
      end
    end
    if(LsuL1Plugin_logic_ls_ctrl_doFlush) begin
      LsuL1Plugin_logic_waysWrite_tag_address = _zz_LsuL1Plugin_logic_waysWrite_tag_address;
    end
  end

  always @(*) begin
    LsuL1Plugin_logic_waysWrite_tag_fault = 1'bx;
    if(LsuL1Plugin_logic_bus_read_rsp_valid) begin
      if(when_LsuL1Plugin_l446) begin
        LsuL1Plugin_logic_waysWrite_tag_fault = LsuL1Plugin_logic_refill_read_faulty;
      end
    end
    if(LsuL1Plugin_logic_ls_ctrl_doFlush) begin
      LsuL1Plugin_logic_waysWrite_tag_fault = _zz_LsuL1Plugin_logic_waysWrite_tag_fault;
    end
  end

  assign LsuL1Plugin_logic_waysWrite_valid = (|LsuL1Plugin_logic_waysWrite_mask);
  assign LsuL1Plugin_logic_banks_0_write_valid = LsuL1Plugin_logic_banksWrite_mask[0];
  assign LsuL1Plugin_logic_banks_0_write_payload_address = LsuL1Plugin_logic_banksWrite_address;
  assign LsuL1Plugin_logic_banks_0_write_payload_data = LsuL1Plugin_logic_banksWrite_writeData;
  assign LsuL1Plugin_logic_banks_0_write_payload_mask = LsuL1Plugin_logic_banksWrite_writeMask;
  assign LsuL1Plugin_logic_banks_0_read_rsp = LsuL1Plugin_logic_banks_0_mem_spinal_port1;
  assign LsuL1Plugin_logic_banks_1_write_valid = LsuL1Plugin_logic_banksWrite_mask[1];
  assign LsuL1Plugin_logic_banks_1_write_payload_address = LsuL1Plugin_logic_banksWrite_address;
  assign LsuL1Plugin_logic_banks_1_write_payload_data = LsuL1Plugin_logic_banksWrite_writeData;
  assign LsuL1Plugin_logic_banks_1_write_payload_mask = LsuL1Plugin_logic_banksWrite_writeMask;
  assign LsuL1Plugin_logic_banks_1_read_rsp = LsuL1Plugin_logic_banks_1_mem_spinal_port1;
  assign _zz_LsuL1Plugin_logic_ways_0_lsuRead_rsp_loaded = LsuL1Plugin_logic_ways_0_mem_spinal_port1;
  assign LsuL1Plugin_logic_ways_0_lsuRead_rsp_loaded = _zz_LsuL1Plugin_logic_ways_0_lsuRead_rsp_loaded[0];
  assign LsuL1Plugin_logic_ways_0_lsuRead_rsp_address = _zz_LsuL1Plugin_logic_ways_0_lsuRead_rsp_loaded[20 : 1];
  assign LsuL1Plugin_logic_ways_0_lsuRead_rsp_fault = _zz_LsuL1Plugin_logic_ways_0_lsuRead_rsp_loaded[21];
  assign _zz_LsuL1Plugin_logic_ways_1_lsuRead_rsp_loaded = LsuL1Plugin_logic_ways_1_mem_spinal_port1;
  assign LsuL1Plugin_logic_ways_1_lsuRead_rsp_loaded = _zz_LsuL1Plugin_logic_ways_1_lsuRead_rsp_loaded[0];
  assign LsuL1Plugin_logic_ways_1_lsuRead_rsp_address = _zz_LsuL1Plugin_logic_ways_1_lsuRead_rsp_loaded[20 : 1];
  assign LsuL1Plugin_logic_ways_1_lsuRead_rsp_fault = _zz_LsuL1Plugin_logic_ways_1_lsuRead_rsp_loaded[21];
  assign _zz_LsuL1Plugin_logic_shared_lsuRead_rsp_plru_0 = LsuL1Plugin_logic_shared_mem_spinal_port1;
  assign LsuL1Plugin_logic_shared_lsuRead_rsp_plru_0 = _zz_LsuL1Plugin_logic_shared_lsuRead_rsp_plru_0_1[0 : 0];
  assign LsuL1Plugin_logic_shared_lsuRead_rsp_dirty = _zz_LsuL1Plugin_logic_shared_lsuRead_rsp_plru_0[2 : 1];
  always @(*) begin
    LsuL1Plugin_logic_refill_slots_0_loadedSet = 1'b0;
    if(LsuL1Plugin_logic_bus_read_rsp_valid) begin
      if(when_LsuL1Plugin_l446) begin
        LsuL1Plugin_logic_refill_slots_0_loadedSet = 1'b1;
      end
    end
  end

  assign LsuL1Plugin_logic_refill_slots_0_loadedDone = (LsuL1Plugin_logic_refill_slots_0_loadedCounter == 1'b1);
  assign LsuL1Plugin_logic_refill_slots_0_fire = ((! execute_freeze_valid) && LsuL1Plugin_logic_refill_slots_0_loadedDone);
  assign LsuL1Plugin_logic_refill_slots_0_free = ((! LsuL1Plugin_logic_refill_slots_0_valid) && 1'b1);
  assign LsuL1Plugin_logic_refill_free = LsuL1Plugin_logic_refill_slots_0_free;
  assign LsuL1Plugin_logic_refill_full = (&(! LsuL1Plugin_logic_refill_slots_0_free));
  assign when_LsuL1Plugin_l358 = LsuL1Plugin_logic_refill_free[0];
  assign LsuL1Plugin_logic_refill_read_arbiter_slotsWithId_0_0 = ((LsuL1Plugin_logic_refill_slots_0_valid && (! LsuL1Plugin_logic_refill_slots_0_cmdSent)) && (LsuL1Plugin_logic_refill_slots_0_victim == 1'b0));
  assign LsuL1Plugin_logic_refill_read_arbiter_hits = LsuL1Plugin_logic_refill_read_arbiter_slotsWithId_0_0;
  assign LsuL1Plugin_logic_refill_read_arbiter_hit = (|LsuL1Plugin_logic_refill_read_arbiter_hits);
  always @(*) begin
    LsuL1Plugin_logic_refill_read_arbiter_oh = (LsuL1Plugin_logic_refill_read_arbiter_hits & 1'b1);
    if(when_LsuL1Plugin_l288) begin
      LsuL1Plugin_logic_refill_read_arbiter_oh = LsuL1Plugin_logic_refill_read_arbiter_lock;
    end
  end

  assign when_LsuL1Plugin_l288 = (|LsuL1Plugin_logic_refill_read_arbiter_lock);
  assign LsuL1Plugin_logic_bus_read_cmd_fire = (LsuL1Plugin_logic_bus_read_cmd_valid && LsuL1Plugin_logic_bus_read_cmd_ready);
  assign LsuL1Plugin_logic_refill_read_cmdAddress = {LsuL1Plugin_logic_refill_slots_0_address[31 : 6],6'h0};
  assign LsuL1Plugin_logic_bus_read_cmd_valid = LsuL1Plugin_logic_refill_read_arbiter_hit;
  assign LsuL1Plugin_logic_bus_read_cmd_payload_address = LsuL1Plugin_logic_refill_read_cmdAddress;
  assign LsuL1Plugin_logic_refill_read_rspAddress = LsuL1Plugin_logic_refill_slots_0_address;
  assign LsuL1Plugin_logic_refill_read_dirty = LsuL1Plugin_logic_refill_slots_0_dirty;
  assign LsuL1Plugin_logic_refill_read_way = LsuL1Plugin_logic_refill_slots_0_way;
  assign LsuL1Plugin_logic_refill_read_rspWithData = 1'b1;
  always @(*) begin
    LsuL1Plugin_logic_refill_read_writeReservation_take = 1'b0;
    if(LsuL1Plugin_logic_bus_read_rsp_valid) begin
      LsuL1Plugin_logic_refill_read_writeReservation_take = 1'b1;
    end
  end

  always @(*) begin
    LsuL1Plugin_logic_refill_read_bankWriteNotif[0] = ((LsuL1Plugin_logic_bus_read_rsp_valid && LsuL1Plugin_logic_refill_read_rspWithData) && (LsuL1Plugin_logic_refill_read_way == 1'b0));
    LsuL1Plugin_logic_refill_read_bankWriteNotif[1] = ((LsuL1Plugin_logic_bus_read_rsp_valid && LsuL1Plugin_logic_refill_read_rspWithData) && (LsuL1Plugin_logic_refill_read_way == 1'b1));
  end

  always @(*) begin
    LsuL1Plugin_logic_banksWrite_mask[0] = LsuL1Plugin_logic_refill_read_bankWriteNotif[0];
    LsuL1Plugin_logic_banksWrite_mask[1] = LsuL1Plugin_logic_refill_read_bankWriteNotif[1];
    if(LsuL1Plugin_logic_ls_ctrl_bankWriteReservation_win) begin
      if(when_LsuL1Plugin_l890) begin
        LsuL1Plugin_logic_banksWrite_mask[0] = ((1'b0 == LsuL1Plugin_logic_ls_ctrl_wayId) && LsuL1Plugin_logic_ls_ctrl_doWrite);
      end
      if(when_LsuL1Plugin_l890_1) begin
        LsuL1Plugin_logic_banksWrite_mask[1] = ((1'b1 == LsuL1Plugin_logic_ls_ctrl_wayId) && LsuL1Plugin_logic_ls_ctrl_doWrite);
      end
    end
    if(LsuL1Plugin_logic_initializerMem_busy) begin
      LsuL1Plugin_logic_banksWrite_mask = 2'b11;
    end
  end

  assign when_LsuL1Plugin_l434 = (LsuL1Plugin_logic_bus_read_rsp_valid && LsuL1Plugin_logic_bus_read_rsp_payload_error);
  always @(*) begin
    LsuL1Plugin_logic_refill_read_fire = 1'b0;
    if(LsuL1Plugin_logic_bus_read_rsp_valid) begin
      if(when_LsuL1Plugin_l446) begin
        LsuL1Plugin_logic_refill_read_fire = 1'b1;
      end
    end
  end

  always @(*) begin
    LsuL1Plugin_logic_refill_read_reservation_take = 1'b0;
    if(LsuL1Plugin_logic_bus_read_rsp_valid) begin
      if(when_LsuL1Plugin_l446) begin
        LsuL1Plugin_logic_refill_read_reservation_take = 1'b1;
      end
    end
  end

  assign LsuL1Plugin_logic_refill_read_faulty = (LsuL1Plugin_logic_refill_read_hadError || LsuL1Plugin_logic_bus_read_rsp_payload_error);
  always @(*) begin
    LsuL1Plugin_logic_refillCompletions = 1'b0;
    if(LsuL1Plugin_logic_bus_read_rsp_valid) begin
      if(when_LsuL1Plugin_l446) begin
        LsuL1Plugin_logic_refillCompletions[0] = 1'b1;
      end
    end
  end

  assign LsuL1Plugin_logic_bus_read_rsp_ready = 1'b1;
  assign when_LsuL1Plugin_l446 = ((LsuL1Plugin_logic_refill_read_wordIndex == 3'b111) || (! LsuL1Plugin_logic_refill_read_rspWithData));
  assign LsuL1_REFILL_BUSY = ((! LsuL1Plugin_logic_refill_slots_0_loaded) && (! LsuL1Plugin_logic_refill_slots_0_loadedSet));
  always @(*) begin
    LsuL1Plugin_logic_writeback_slots_0_fire = 1'b0;
    if(LsuL1Plugin_logic_bus_write_rsp_valid) begin
      LsuL1Plugin_logic_writeback_slots_0_fire = 1'b1;
    end
  end

  assign LsuL1Plugin_logic_writeback_slots_0_timer_done = (LsuL1Plugin_logic_writeback_slots_0_timer_counter == 1'b1);
  assign when_LsuL1Plugin_l509 = (LsuL1Plugin_logic_writeback_slots_0_timer_done && (LsuL1Plugin_logic_writeback_slots_0_fire || (! LsuL1Plugin_logic_writeback_slots_0_busy)));
  assign LsuL1Plugin_logic_writeback_slots_0_free = (! LsuL1Plugin_logic_writeback_slots_0_valid);
  assign LsuL1_WRITEBACK_BUSY = (LsuL1Plugin_logic_writeback_slots_0_valid || LsuL1Plugin_logic_writeback_slots_0_fire);
  assign LsuL1Plugin_logic_writebackBusy = (|LsuL1Plugin_logic_writeback_slots_0_valid);
  assign LsuL1Plugin_logic_writeback_free = LsuL1Plugin_logic_writeback_slots_0_free;
  assign LsuL1Plugin_logic_writeback_full = (&(! LsuL1Plugin_logic_writeback_slots_0_free));
  always @(*) begin
    LsuL1Plugin_logic_writeback_push_valid = 1'b0;
    if(LsuL1Plugin_logic_ls_ctrl_doFlush) begin
      LsuL1Plugin_logic_writeback_push_valid = 1'b1;
    end
    if(LsuL1Plugin_logic_ls_ctrl_doRefill) begin
      LsuL1Plugin_logic_writeback_push_valid = LsuL1Plugin_logic_ls_ctrl_refillWayNeedWriteback;
    end
    if(LsuL1Plugin_logic_ls_ctrl_preventSideEffects) begin
      LsuL1Plugin_logic_writeback_push_valid = 1'b0;
    end
  end

  always @(*) begin
    LsuL1Plugin_logic_writeback_push_payload_address = 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
    if(LsuL1Plugin_logic_ls_ctrl_doFlush) begin
      LsuL1Plugin_logic_writeback_push_payload_address = ({6'd0,{_zz_LsuL1Plugin_logic_waysWrite_tag_address,toplevel_execute_ctrl4_down_LsuL1_MIXED_ADDRESS_lane0[11 : 6]}} <<< 3'd6);
    end
    if(LsuL1Plugin_logic_ls_ctrl_doRefill) begin
      LsuL1Plugin_logic_writeback_push_payload_address = ({6'd0,{_zz_LsuL1Plugin_logic_writeback_push_payload_address,toplevel_execute_ctrl4_down_LsuL1_MIXED_ADDRESS_lane0[11 : 6]}} <<< 3'd6);
    end
  end

  always @(*) begin
    LsuL1Plugin_logic_writeback_push_payload_way = 1'bx;
    if(LsuL1Plugin_logic_ls_ctrl_doFlush) begin
      LsuL1Plugin_logic_writeback_push_payload_way = LsuL1Plugin_logic_ls_ctrl_needFlushSel;
    end
    if(LsuL1Plugin_logic_ls_ctrl_doRefill) begin
      LsuL1Plugin_logic_writeback_push_payload_way = LsuL1Plugin_logic_ls_ctrl_targetWay;
    end
  end

  assign when_LsuL1Plugin_l532 = LsuL1Plugin_logic_writeback_free[0];
  assign LsuL1Plugin_logic_writeback_read_arbiter_slotsWithId_0_0 = (LsuL1Plugin_logic_writeback_slots_0_valid && (! LsuL1Plugin_logic_writeback_slots_0_readCmdDone));
  assign LsuL1Plugin_logic_writeback_read_arbiter_hits = LsuL1Plugin_logic_writeback_read_arbiter_slotsWithId_0_0;
  assign LsuL1Plugin_logic_writeback_read_arbiter_hit = (|LsuL1Plugin_logic_writeback_read_arbiter_hits);
  always @(*) begin
    LsuL1Plugin_logic_writeback_read_arbiter_oh = (LsuL1Plugin_logic_writeback_read_arbiter_hits & 1'b1);
    if(when_LsuL1Plugin_l288_1) begin
      LsuL1Plugin_logic_writeback_read_arbiter_oh = LsuL1Plugin_logic_writeback_read_arbiter_lock;
    end
  end

  assign when_LsuL1Plugin_l288_1 = (|LsuL1Plugin_logic_writeback_read_arbiter_lock);
  assign LsuL1Plugin_logic_writeback_read_address = LsuL1Plugin_logic_writeback_slots_0_address;
  assign LsuL1Plugin_logic_writeback_read_way = LsuL1Plugin_logic_writeback_slots_0_way;
  assign LsuL1Plugin_logic_writeback_read_slotRead_valid = LsuL1Plugin_logic_writeback_read_arbiter_hit;
  assign LsuL1Plugin_logic_writeback_read_slotRead_payload_wordIndex = LsuL1Plugin_logic_writeback_read_wordIndex;
  assign LsuL1Plugin_logic_writeback_read_slotRead_payload_way = LsuL1Plugin_logic_writeback_read_way;
  assign LsuL1Plugin_logic_writeback_read_slotRead_payload_last = (LsuL1Plugin_logic_writeback_read_wordIndex == 3'b111);
  assign when_LsuL1Plugin_l577 = (LsuL1Plugin_logic_writeback_read_slotRead_valid && LsuL1Plugin_logic_writeback_read_slotRead_payload_last);
  always @(*) begin
    LsuL1Plugin_logic_banks_0_read_cmd_valid = LsuL1Plugin_logic_banks_0_usedByWriteback;
    if(when_LsuL1Plugin_l690) begin
      LsuL1Plugin_logic_banks_0_read_cmd_valid = 1'b1;
    end
  end

  assign LsuL1Plugin_logic_banks_0_usedByWriteback = (LsuL1Plugin_logic_writeback_read_slotRead_valid && (LsuL1Plugin_logic_writeback_read_way == 1'b0));
  always @(*) begin
    LsuL1Plugin_logic_banks_0_read_cmd_payload = {LsuL1Plugin_logic_writeback_read_address[11 : 6],LsuL1Plugin_logic_writeback_read_wordIndex};
    if(when_LsuL1Plugin_l691) begin
      LsuL1Plugin_logic_banks_0_read_cmd_payload = LsuL1Plugin_logic_ls_rb0_readAddress;
    end
  end

  always @(*) begin
    LsuL1Plugin_logic_banks_1_read_cmd_valid = LsuL1Plugin_logic_banks_1_usedByWriteback;
    if(when_LsuL1Plugin_l690_1) begin
      LsuL1Plugin_logic_banks_1_read_cmd_valid = 1'b1;
    end
  end

  assign LsuL1Plugin_logic_banks_1_usedByWriteback = (LsuL1Plugin_logic_writeback_read_slotRead_valid && (LsuL1Plugin_logic_writeback_read_way == 1'b1));
  always @(*) begin
    LsuL1Plugin_logic_banks_1_read_cmd_payload = {LsuL1Plugin_logic_writeback_read_address[11 : 6],LsuL1Plugin_logic_writeback_read_wordIndex};
    if(when_LsuL1Plugin_l691_1) begin
      LsuL1Plugin_logic_banks_1_read_cmd_payload = LsuL1Plugin_logic_ls_rb0_readAddress;
    end
  end

  assign LsuL1Plugin_logic_writeback_read_readedData = _zz_LsuL1Plugin_logic_writeback_read_readedData;
  assign LsuL1Plugin_logic_writeback_write_arbiter_slotsWithId_0_0 = ((LsuL1Plugin_logic_writeback_slots_0_valid && LsuL1Plugin_logic_writeback_slots_0_victimBufferReady) && (! LsuL1Plugin_logic_writeback_slots_0_writeCmdDone));
  assign LsuL1Plugin_logic_writeback_write_arbiter_hits = LsuL1Plugin_logic_writeback_write_arbiter_slotsWithId_0_0;
  assign LsuL1Plugin_logic_writeback_write_arbiter_hit = (|LsuL1Plugin_logic_writeback_write_arbiter_hits);
  always @(*) begin
    LsuL1Plugin_logic_writeback_write_arbiter_oh = (LsuL1Plugin_logic_writeback_write_arbiter_hits & 1'b1);
    if(when_LsuL1Plugin_l288_2) begin
      LsuL1Plugin_logic_writeback_write_arbiter_oh = LsuL1Plugin_logic_writeback_write_arbiter_lock;
    end
  end

  assign when_LsuL1Plugin_l288_2 = (|LsuL1Plugin_logic_writeback_write_arbiter_lock);
  assign LsuL1Plugin_logic_writeback_write_last = (LsuL1Plugin_logic_writeback_write_wordIndex == 3'b111);
  assign LsuL1Plugin_logic_writeback_write_bufferRead_valid = LsuL1Plugin_logic_writeback_write_arbiter_hit;
  assign LsuL1Plugin_logic_writeback_write_bufferRead_payload_last = LsuL1Plugin_logic_writeback_write_last;
  assign LsuL1Plugin_logic_writeback_write_bufferRead_payload_address = LsuL1Plugin_logic_writeback_slots_0_address;
  assign LsuL1Plugin_logic_writeback_write_bufferRead_fire = (LsuL1Plugin_logic_writeback_write_bufferRead_valid && LsuL1Plugin_logic_writeback_write_bufferRead_ready);
  assign when_LsuL1Plugin_l651 = (LsuL1Plugin_logic_writeback_write_bufferRead_fire && LsuL1Plugin_logic_writeback_write_last);
  always @(*) begin
    LsuL1Plugin_logic_writeback_write_bufferRead_ready = LsuL1Plugin_logic_writeback_write_cmd_ready;
    if(when_Stream_l393_2) begin
      LsuL1Plugin_logic_writeback_write_bufferRead_ready = 1'b1;
    end
  end

  assign when_Stream_l393_2 = (! LsuL1Plugin_logic_writeback_write_cmd_valid);
  assign LsuL1Plugin_logic_writeback_write_cmd_valid = LsuL1Plugin_logic_writeback_write_bufferRead_rValid;
  assign LsuL1Plugin_logic_writeback_write_cmd_payload_address = LsuL1Plugin_logic_writeback_write_bufferRead_rData_address;
  assign LsuL1Plugin_logic_writeback_write_cmd_payload_last = LsuL1Plugin_logic_writeback_write_bufferRead_rData_last;
  assign _zz_LsuL1Plugin_logic_writeback_write_word = LsuL1Plugin_logic_writeback_write_wordIndex;
  assign LsuL1Plugin_logic_writeback_write_word = LsuL1Plugin_logic_writeback_victimBuffer_spinal_port1;
  assign LsuL1Plugin_logic_bus_write_cmd_valid = LsuL1Plugin_logic_writeback_write_cmd_valid;
  assign LsuL1Plugin_logic_writeback_write_cmd_ready = LsuL1Plugin_logic_bus_write_cmd_ready;
  assign LsuL1Plugin_logic_bus_write_cmd_payload_fragment_address = LsuL1Plugin_logic_writeback_write_cmd_payload_address;
  assign LsuL1Plugin_logic_bus_write_cmd_payload_fragment_data = LsuL1Plugin_logic_writeback_write_word;
  assign LsuL1Plugin_logic_bus_write_cmd_payload_last = LsuL1Plugin_logic_writeback_write_cmd_payload_last;
  assign LsuL1Plugin_logic_ls_rb0_readAddress = toplevel_execute_ctrl2_down_LsuL1_MIXED_ADDRESS_lane0[11 : 3];
  always @(*) begin
    toplevel_execute_ctrl2_down_LsuL1Plugin_logic_BANK_BUSY_lane0[0] = LsuL1Plugin_logic_banks_0_usedByWriteback;
    toplevel_execute_ctrl2_down_LsuL1Plugin_logic_BANK_BUSY_lane0[1] = LsuL1Plugin_logic_banks_1_usedByWriteback;
  end

  assign when_LsuL1Plugin_l690 = (! execute_freeze_valid);
  assign when_LsuL1Plugin_l691 = (! LsuL1Plugin_logic_banks_0_usedByWriteback);
  assign when_LsuL1Plugin_l690_1 = (! execute_freeze_valid);
  assign when_LsuL1Plugin_l691_1 = (! LsuL1Plugin_logic_banks_1_usedByWriteback);
  assign when_LsuL1Plugin_l706 = (! execute_freeze_valid);
  assign toplevel_execute_ctrl3_down_LsuL1Plugin_logic_BANKS_WORDS_lane0_0 = LsuL1Plugin_logic_banks_0_read_rsp;
  always @(*) begin
    toplevel_execute_ctrl3_down_LsuL1Plugin_logic_BANK_BUSY_REMAPPED_lane0[0] = (toplevel_execute_ctrl3_down_LsuL1Plugin_logic_BANK_BUSY_lane0[1'b0] || LsuL1Plugin_logic_ls_rb1_onBanks_0_busyReg);
    toplevel_execute_ctrl3_down_LsuL1Plugin_logic_BANK_BUSY_REMAPPED_lane0[1] = (toplevel_execute_ctrl3_down_LsuL1Plugin_logic_BANK_BUSY_lane0[1'b1] || LsuL1Plugin_logic_ls_rb1_onBanks_1_busyReg);
  end

  assign when_LsuL1Plugin_l706_1 = (! execute_freeze_valid);
  assign toplevel_execute_ctrl3_down_LsuL1Plugin_logic_BANKS_WORDS_lane0_1 = LsuL1Plugin_logic_banks_1_read_rsp;
  assign toplevel_execute_ctrl3_down_LsuL1Plugin_logic_BANKS_MUXES_lane0_0 = _zz_toplevel_execute_ctrl3_down_LsuL1Plugin_logic_BANKS_MUXES_lane0_0;
  assign toplevel_execute_ctrl3_down_LsuL1Plugin_logic_BANKS_MUXES_lane0_1 = _zz_toplevel_execute_ctrl3_down_LsuL1Plugin_logic_BANKS_MUXES_lane0_1;
  assign _zz_toplevel_execute_ctrl4_down_LsuL1Plugin_logic_MUXED_DATA_lane0 = toplevel_execute_ctrl4_down_LsuL1Plugin_logic_WAYS_HITS_lane0[0];
  assign _zz_toplevel_execute_ctrl4_down_LsuL1Plugin_logic_MUXED_DATA_lane0_1 = toplevel_execute_ctrl4_down_LsuL1Plugin_logic_WAYS_HITS_lane0[1];
  assign toplevel_execute_ctrl4_down_LsuL1Plugin_logic_MUXED_DATA_lane0 = ((_zz_toplevel_execute_ctrl4_down_LsuL1Plugin_logic_MUXED_DATA_lane0 ? toplevel_execute_ctrl4_down_LsuL1Plugin_logic_BANKS_MUXES_lane0_0 : 32'h0) | (_zz_toplevel_execute_ctrl4_down_LsuL1Plugin_logic_MUXED_DATA_lane0_1 ? toplevel_execute_ctrl4_down_LsuL1Plugin_logic_BANKS_MUXES_lane0_1 : 32'h0));
  always @(*) begin
    toplevel_execute_ctrl3_down_LsuL1Plugin_logic_WRITE_TO_READ_HAZARDS_lane0[0] = ((toplevel_execute_ctrl2_down_LsuL1Plugin_logic_EVENT_WRITE_VALID_lane0 && (toplevel_execute_ctrl2_down_LsuL1Plugin_logic_EVENT_WRITE_ADDRESS_lane0[31 : 2] == toplevel_execute_ctrl3_down_LsuL1_PHYSICAL_ADDRESS_lane0[31 : 2])) && 1'b1);
    toplevel_execute_ctrl3_down_LsuL1Plugin_logic_WRITE_TO_READ_HAZARDS_lane0[1] = ((toplevel_execute_ctrl3_down_LsuL1Plugin_logic_EVENT_WRITE_VALID_lane0 && (toplevel_execute_ctrl3_down_LsuL1Plugin_logic_EVENT_WRITE_ADDRESS_lane0[31 : 2] == toplevel_execute_ctrl3_down_LsuL1_PHYSICAL_ADDRESS_lane0[31 : 2])) && 1'b1);
  end

  assign LsuL1Plugin_logic_shared_lsuRead_cmd_valid = (! execute_freeze_valid);
  assign LsuL1Plugin_logic_shared_lsuRead_cmd_payload = toplevel_execute_ctrl2_down_LsuL1_MIXED_ADDRESS_lane0[11 : 6];
  assign toplevel_execute_ctrl2_down_LsuL1Plugin_logic_ls_rt0_SHARED_BYPASS_VALID_lane0 = (LsuL1Plugin_logic_shared_write_valid && (LsuL1Plugin_logic_shared_write_payload_address == toplevel_execute_ctrl2_down_LsuL1_MIXED_ADDRESS_lane0[11 : 6]));
  assign toplevel_execute_ctrl2_down_LsuL1Plugin_logic_ls_rt0_SHARED_BYPASS_VALUE_lane0_plru_0 = LsuL1Plugin_logic_shared_write_payload_data_plru_0;
  assign toplevel_execute_ctrl2_down_LsuL1Plugin_logic_ls_rt0_SHARED_BYPASS_VALUE_lane0_dirty = LsuL1Plugin_logic_shared_write_payload_data_dirty;
  assign LsuL1Plugin_logic_ways_0_lsuRead_cmd_valid = (! execute_freeze_valid);
  assign LsuL1Plugin_logic_ways_0_lsuRead_cmd_payload = toplevel_execute_ctrl2_down_LsuL1_MIXED_ADDRESS_lane0[11 : 6];
  assign LsuL1Plugin_logic_ways_1_lsuRead_cmd_valid = (! execute_freeze_valid);
  assign LsuL1Plugin_logic_ways_1_lsuRead_cmd_payload = toplevel_execute_ctrl2_down_LsuL1_MIXED_ADDRESS_lane0[11 : 6];
  always @(*) begin
    toplevel_execute_ctrl3_up_LsuL1Plugin_logic_SHARED_lane0_plru_0 = LsuL1Plugin_logic_shared_lsuRead_rsp_plru_0;
    if(toplevel_execute_ctrl3_down_LsuL1Plugin_logic_ls_rt0_SHARED_BYPASS_VALID_lane0) begin
      toplevel_execute_ctrl3_up_LsuL1Plugin_logic_SHARED_lane0_plru_0 = toplevel_execute_ctrl3_down_LsuL1Plugin_logic_ls_rt0_SHARED_BYPASS_VALUE_lane0_plru_0;
    end
  end

  always @(*) begin
    toplevel_execute_ctrl3_up_LsuL1Plugin_logic_SHARED_lane0_dirty = LsuL1Plugin_logic_shared_lsuRead_rsp_dirty;
    if(toplevel_execute_ctrl3_down_LsuL1Plugin_logic_ls_rt0_SHARED_BYPASS_VALID_lane0) begin
      toplevel_execute_ctrl3_up_LsuL1Plugin_logic_SHARED_lane0_dirty = toplevel_execute_ctrl3_down_LsuL1Plugin_logic_ls_rt0_SHARED_BYPASS_VALUE_lane0_dirty;
    end
  end

  assign toplevel_execute_ctrl3_down_LsuL1Plugin_logic_WAYS_TAGS_lane0_0_loaded = LsuL1Plugin_logic_ways_0_lsuRead_rsp_loaded;
  assign toplevel_execute_ctrl3_down_LsuL1Plugin_logic_WAYS_TAGS_lane0_0_address = LsuL1Plugin_logic_ways_0_lsuRead_rsp_address;
  assign toplevel_execute_ctrl3_down_LsuL1Plugin_logic_WAYS_TAGS_lane0_0_fault = LsuL1Plugin_logic_ways_0_lsuRead_rsp_fault;
  assign toplevel_execute_ctrl3_down_LsuL1Plugin_logic_WAYS_TAGS_lane0_1_loaded = LsuL1Plugin_logic_ways_1_lsuRead_rsp_loaded;
  assign toplevel_execute_ctrl3_down_LsuL1Plugin_logic_WAYS_TAGS_lane0_1_address = LsuL1Plugin_logic_ways_1_lsuRead_rsp_address;
  assign toplevel_execute_ctrl3_down_LsuL1Plugin_logic_WAYS_TAGS_lane0_1_fault = LsuL1Plugin_logic_ways_1_lsuRead_rsp_fault;
  assign LsuL1Plugin_logic_ls_sharedBypassers_0_hit = (LsuL1Plugin_logic_shared_write_valid && (LsuL1Plugin_logic_shared_write_payload_address == toplevel_execute_ctrl3_down_LsuL1_MIXED_ADDRESS_lane0[11 : 6]));
  assign toplevel_execute_ctrl3_LsuL1Plugin_logic_SHARED_lane0_bypass_plru_0 = (LsuL1Plugin_logic_ls_sharedBypassers_0_hit ? LsuL1Plugin_logic_shared_write_payload_data_plru_0 : toplevel_execute_ctrl3_up_LsuL1Plugin_logic_SHARED_lane0_plru_0);
  assign toplevel_execute_ctrl3_LsuL1Plugin_logic_SHARED_lane0_bypass_dirty = (LsuL1Plugin_logic_ls_sharedBypassers_0_hit ? LsuL1Plugin_logic_shared_write_payload_data_dirty : toplevel_execute_ctrl3_up_LsuL1Plugin_logic_SHARED_lane0_dirty);
  always @(*) begin
    toplevel_execute_ctrl3_down_LsuL1Plugin_logic_WAYS_HITS_lane0[0] = (toplevel_execute_ctrl3_down_LsuL1Plugin_logic_WAYS_TAGS_lane0_0_loaded && (toplevel_execute_ctrl3_down_LsuL1Plugin_logic_WAYS_TAGS_lane0_0_address == toplevel_execute_ctrl3_down_LsuL1_PHYSICAL_ADDRESS_lane0[31 : 12]));
    toplevel_execute_ctrl3_down_LsuL1Plugin_logic_WAYS_HITS_lane0[1] = (toplevel_execute_ctrl3_down_LsuL1Plugin_logic_WAYS_TAGS_lane0_1_loaded && (toplevel_execute_ctrl3_down_LsuL1Plugin_logic_WAYS_TAGS_lane0_1_address == toplevel_execute_ctrl3_down_LsuL1_PHYSICAL_ADDRESS_lane0[31 : 12]));
  end

  assign toplevel_execute_ctrl4_down_LsuL1Plugin_logic_WAYS_HIT_lane0 = (|toplevel_execute_ctrl4_down_LsuL1Plugin_logic_WAYS_HITS_lane0);
  assign toplevel_execute_ctrl4_down_LsuL1Plugin_logic_NEED_UNIQUE_lane0 = (toplevel_execute_ctrl4_down_LsuL1_STORE_lane0 || toplevel_execute_ctrl4_down_LsuL1_ATOMIC_lane0);
  assign LsuL1Plugin_logic_ls_ctrl_plruLogic_core_evict_logic_0_state = LsuL1Plugin_logic_ls_ctrl_plruLogic_core_io_context_state_0[0];
  assign LsuL1Plugin_logic_ls_ctrl_plruLogic_core_evict_sel_0 = (! LsuL1Plugin_logic_ls_ctrl_plruLogic_core_evict_logic_0_state);
  assign LsuL1Plugin_logic_ls_ctrl_plruLogic_core_io_evict_id = LsuL1Plugin_logic_ls_ctrl_plruLogic_core_evict_sel_0;
  assign LsuL1Plugin_logic_ls_ctrl_plruLogic_core_io_update_state_0[0] = LsuL1Plugin_logic_ls_ctrl_plruLogic_core_io_update_id[0];
  assign LsuL1Plugin_logic_ls_ctrl_plruLogic_core_io_context_state_0 = toplevel_execute_ctrl4_down_LsuL1Plugin_logic_SHARED_lane0_plru_0;
  always @(*) begin
    LsuL1Plugin_logic_ls_ctrl_wayWriteReservation_take = 1'b0;
    if(LsuL1Plugin_logic_ls_ctrl_doFlush) begin
      LsuL1Plugin_logic_ls_ctrl_wayWriteReservation_take = 1'b1;
    end
  end

  assign LsuL1Plugin_logic_ls_ctrl_bankWriteReservation_take = 1'b0;
  assign LsuL1Plugin_logic_ls_ctrl_refillWayWithoutUpdate = LsuL1Plugin_logic_ls_ctrl_plruLogic_core_io_evict_id;
  assign LsuL1Plugin_logic_ls_ctrl_refillWayNeedWriteback = _zz_LsuL1Plugin_logic_ls_ctrl_refillWayNeedWriteback[LsuL1Plugin_logic_ls_ctrl_refillWayWithoutUpdate];
  assign LsuL1Plugin_logic_ls_ctrl_refillHazards = (LsuL1Plugin_logic_refill_slots_0_valid && (LsuL1Plugin_logic_refill_slots_0_address[11 : 6] == toplevel_execute_ctrl4_down_LsuL1_PHYSICAL_ADDRESS_lane0[11 : 6]));
  assign LsuL1Plugin_logic_ls_ctrl_writebackHazards = (LsuL1Plugin_logic_writeback_slots_0_valid && (LsuL1Plugin_logic_writeback_slots_0_address[11 : 6] == toplevel_execute_ctrl4_down_LsuL1_PHYSICAL_ADDRESS_lane0[11 : 6]));
  assign LsuL1Plugin_logic_ls_ctrl_refillHazard = (|LsuL1Plugin_logic_ls_ctrl_refillHazards);
  assign LsuL1Plugin_logic_ls_ctrl_writebackHazard = (|LsuL1Plugin_logic_ls_ctrl_writebackHazards);
  assign LsuL1Plugin_logic_ls_ctrl_wasDirty = (|(toplevel_execute_ctrl4_down_LsuL1Plugin_logic_SHARED_lane0_dirty & toplevel_execute_ctrl4_down_LsuL1Plugin_logic_WAYS_HITS_lane0));
  assign LsuL1Plugin_logic_ls_ctrl_loadedDirties = ({toplevel_execute_ctrl4_down_LsuL1Plugin_logic_WAYS_TAGS_lane0_1_loaded,toplevel_execute_ctrl4_down_LsuL1Plugin_logic_WAYS_TAGS_lane0_0_loaded} & toplevel_execute_ctrl4_down_LsuL1Plugin_logic_SHARED_lane0_dirty);
  assign LsuL1Plugin_logic_ls_ctrl_refillWayWasDirty = LsuL1Plugin_logic_ls_ctrl_loadedDirties[LsuL1Plugin_logic_ls_ctrl_refillWayWithoutUpdate];
  assign LsuL1Plugin_logic_ls_ctrl_writeToReadHazard = 1'b0;
  assign LsuL1Plugin_logic_ls_ctrl_bankNotRead = (|(toplevel_execute_ctrl4_down_LsuL1Plugin_logic_BANK_BUSY_REMAPPED_lane0 & toplevel_execute_ctrl4_down_LsuL1Plugin_logic_WAYS_HITS_lane0));
  assign LsuL1Plugin_logic_ls_ctrl_loadHazard = ((toplevel_execute_ctrl4_down_LsuL1_LOAD_lane0 && (! toplevel_execute_ctrl4_down_LsuL1_PREFETCH_lane0)) && (LsuL1Plugin_logic_ls_ctrl_bankNotRead || LsuL1Plugin_logic_ls_ctrl_writeToReadHazard));
  assign LsuL1Plugin_logic_ls_ctrl_storeHazard = ((toplevel_execute_ctrl4_down_LsuL1_STORE_lane0 && (! toplevel_execute_ctrl4_down_LsuL1_PREFETCH_lane0)) && (! LsuL1Plugin_logic_ls_ctrl_bankWriteReservation_win));
  assign LsuL1Plugin_logic_ls_ctrl_flushHazard = (toplevel_execute_ctrl4_down_LsuL1_FLUSH_lane0 && (! LsuL1Plugin_logic_ls_ctrl_wayWriteReservation_win));
  assign LsuL1Plugin_logic_ls_ctrl_coherencyHazard = 1'b0;
  assign toplevel_execute_ctrl4_down_LsuL1Plugin_logic_HAZARD_FORCED_lane0 = 1'b0;
  assign toplevel_execute_ctrl4_down_LsuL1_HAZARD_lane0 = (((((LsuL1Plugin_logic_ls_ctrl_hazardReg || LsuL1Plugin_logic_ls_ctrl_loadHazard) || LsuL1Plugin_logic_ls_ctrl_refillHazard) || LsuL1Plugin_logic_ls_ctrl_storeHazard) || LsuL1Plugin_logic_ls_ctrl_coherencyHazard) || toplevel_execute_ctrl4_down_LsuL1Plugin_logic_HAZARD_FORCED_lane0);
  assign toplevel_execute_ctrl4_down_LsuL1_FLUSH_HAZARD_lane0 = (LsuL1Plugin_logic_ls_ctrl_flushHazardReg || LsuL1Plugin_logic_ls_ctrl_flushHazard);
  assign toplevel_execute_ctrl4_down_LsuL1_MISS_lane0 = (! toplevel_execute_ctrl4_down_LsuL1Plugin_logic_WAYS_HIT_lane0);
  assign toplevel_execute_ctrl4_down_LsuL1_FAULT_lane0 = ((toplevel_execute_ctrl4_down_LsuL1Plugin_logic_WAYS_HIT_lane0 && (|(toplevel_execute_ctrl4_down_LsuL1Plugin_logic_WAYS_HITS_lane0 & {toplevel_execute_ctrl4_down_LsuL1Plugin_logic_WAYS_TAGS_lane0_1_fault,toplevel_execute_ctrl4_down_LsuL1Plugin_logic_WAYS_TAGS_lane0_0_fault}))) && (! toplevel_execute_ctrl4_down_LsuL1_FLUSH_lane0));
  assign toplevel_execute_ctrl4_down_LsuL1_MISS_UNIQUE_lane0 = ((toplevel_execute_ctrl4_down_LsuL1Plugin_logic_WAYS_HIT_lane0 && toplevel_execute_ctrl4_down_LsuL1Plugin_logic_NEED_UNIQUE_lane0) && 1'b0);
  assign toplevel_execute_ctrl4_down_LsuL1_REFILL_HIT_lane0 = LsuL1Plugin_logic_ls_ctrl_refillHazard;
  assign LsuL1Plugin_logic_ls_ctrl_canRefill = (((LsuL1Plugin_logic_ls_ctrl_wayWriteReservation_win && (! (LsuL1Plugin_logic_ls_ctrl_refillWayNeedWriteback && LsuL1Plugin_logic_writeback_full))) && (! LsuL1Plugin_logic_refill_full)) && (! LsuL1Plugin_logic_ls_ctrl_writebackHazard));
  assign LsuL1Plugin_logic_ls_ctrl_canFlush = (((LsuL1Plugin_logic_ls_ctrl_wayWriteReservation_win && (! LsuL1Plugin_logic_writeback_full)) && (! (|LsuL1Plugin_logic_refill_slots_0_valid))) && (! LsuL1Plugin_logic_ls_ctrl_writebackHazard));
  assign LsuL1Plugin_logic_ls_ctrl_needFlushs = LsuL1Plugin_logic_ls_ctrl_loadedDirties;
  assign _zz_LsuL1Plugin_logic_ls_ctrl_needFlushs_bools_0 = LsuL1Plugin_logic_ls_ctrl_needFlushs;
  assign LsuL1Plugin_logic_ls_ctrl_needFlushs_bools_0 = _zz_LsuL1Plugin_logic_ls_ctrl_needFlushs_bools_0[0];
  assign LsuL1Plugin_logic_ls_ctrl_needFlushs_bools_1 = _zz_LsuL1Plugin_logic_ls_ctrl_needFlushs_bools_0[1];
  always @(*) begin
    _zz_LsuL1Plugin_logic_ls_ctrl_needFlushOh[0] = (LsuL1Plugin_logic_ls_ctrl_needFlushs_bools_0 && (! 1'b0));
    _zz_LsuL1Plugin_logic_ls_ctrl_needFlushOh[1] = (LsuL1Plugin_logic_ls_ctrl_needFlushs_bools_1 && (! LsuL1Plugin_logic_ls_ctrl_needFlushs_bools_0));
  end

  assign LsuL1Plugin_logic_ls_ctrl_needFlushOh = _zz_LsuL1Plugin_logic_ls_ctrl_needFlushOh;
  assign _zz_LsuL1Plugin_logic_ls_ctrl_needFlushSel = LsuL1Plugin_logic_ls_ctrl_needFlushOh[1];
  assign LsuL1Plugin_logic_ls_ctrl_needFlushSel = _zz_LsuL1Plugin_logic_ls_ctrl_needFlushSel;
  assign LsuL1Plugin_logic_ls_ctrl_isAccess = (! toplevel_execute_ctrl4_down_LsuL1_FLUSH_lane0);
  assign LsuL1Plugin_logic_ls_ctrl_askRefill = ((LsuL1Plugin_logic_ls_ctrl_isAccess && toplevel_execute_ctrl4_down_LsuL1_MISS_lane0) && LsuL1Plugin_logic_ls_ctrl_canRefill);
  assign LsuL1Plugin_logic_ls_ctrl_askUpgrade = ((LsuL1Plugin_logic_ls_ctrl_isAccess && toplevel_execute_ctrl4_down_LsuL1_MISS_UNIQUE_lane0) && LsuL1Plugin_logic_ls_ctrl_canRefill);
  assign LsuL1Plugin_logic_ls_ctrl_askFlush = ((toplevel_execute_ctrl4_down_LsuL1_FLUSH_lane0 && LsuL1Plugin_logic_ls_ctrl_canFlush) && (|LsuL1Plugin_logic_ls_ctrl_needFlushs));
  assign LsuL1Plugin_logic_ls_ctrl_doRefill = (toplevel_execute_ctrl4_down_LsuL1_SEL_lane0 && LsuL1Plugin_logic_ls_ctrl_askRefill);
  assign LsuL1Plugin_logic_ls_ctrl_doUpgrade = (toplevel_execute_ctrl4_down_LsuL1_SEL_lane0 && LsuL1Plugin_logic_ls_ctrl_askUpgrade);
  assign LsuL1Plugin_logic_ls_ctrl_doFlush = (toplevel_execute_ctrl4_down_LsuL1_SEL_lane0 && LsuL1Plugin_logic_ls_ctrl_askFlush);
  assign LsuL1Plugin_logic_ls_ctrl_doWrite = ((((toplevel_execute_ctrl4_down_LsuL1_SEL_lane0 && toplevel_execute_ctrl4_down_LsuL1_STORE_lane0) && toplevel_execute_ctrl4_down_LsuL1Plugin_logic_WAYS_HIT_lane0) && _zz_LsuL1Plugin_logic_ls_ctrl_doWrite[0]) && (! toplevel_execute_ctrl4_down_LsuL1_SKIP_WRITE_lane0));
  assign LsuL1Plugin_logic_ls_ctrl_wayId = _zz_toplevel_execute_ctrl4_down_LsuL1Plugin_logic_MUXED_DATA_lane0_1;
  assign LsuL1Plugin_logic_ls_ctrl_targetWay = (LsuL1Plugin_logic_ls_ctrl_askUpgrade ? LsuL1Plugin_logic_ls_ctrl_wayId : LsuL1Plugin_logic_ls_ctrl_refillWayWithoutUpdate);
  always @(*) begin
    LsuL1Plugin_logic_ls_ctrl_plruLogic_core_io_update_id = LsuL1Plugin_logic_ls_ctrl_wayId;
    if(LsuL1Plugin_logic_ls_ctrl_doRefill) begin
      LsuL1Plugin_logic_ls_ctrl_plruLogic_core_io_update_id = LsuL1Plugin_logic_ls_ctrl_targetWay;
    end
  end

  assign LsuL1Plugin_logic_ls_ctrl_doRefillPush = (LsuL1Plugin_logic_ls_ctrl_doRefill || LsuL1Plugin_logic_ls_ctrl_doUpgrade);
  always @(*) begin
    LsuL1Plugin_logic_refill_push_valid = LsuL1Plugin_logic_ls_ctrl_doRefillPush;
    if(LsuL1Plugin_logic_ls_ctrl_preventSideEffects) begin
      LsuL1Plugin_logic_refill_push_valid = 1'b0;
    end
  end

  assign LsuL1Plugin_logic_refill_push_payload_address = toplevel_execute_ctrl4_down_LsuL1_PHYSICAL_ADDRESS_lane0;
  assign LsuL1Plugin_logic_refill_push_payload_unique = toplevel_execute_ctrl4_down_LsuL1Plugin_logic_NEED_UNIQUE_lane0;
  assign LsuL1Plugin_logic_refill_push_payload_data = LsuL1Plugin_logic_ls_ctrl_askRefill;
  always @(*) begin
    LsuL1Plugin_logic_refill_push_payload_way = LsuL1Plugin_logic_ls_ctrl_targetWay;
    if(LsuL1Plugin_logic_ls_ctrl_askUpgrade) begin
      LsuL1Plugin_logic_refill_push_payload_way = LsuL1Plugin_logic_ls_ctrl_wayId;
    end
  end

  always @(*) begin
    LsuL1Plugin_logic_refill_push_payload_victim = ((LsuL1Plugin_logic_ls_ctrl_refillWayNeedWriteback && LsuL1Plugin_logic_ls_ctrl_refillWayWasDirty) ? LsuL1Plugin_logic_writeback_free : 1'b0);
    if(LsuL1Plugin_logic_ls_ctrl_askUpgrade) begin
      LsuL1Plugin_logic_refill_push_payload_victim = 1'b0;
    end
  end

  assign LsuL1Plugin_logic_refill_push_payload_dirty = toplevel_execute_ctrl4_down_LsuL1_STORE_lane0;
  assign toplevel_execute_ctrl4_down_LsuL1_WAIT_REFILL_lane0 = (LsuL1Plugin_logic_ls_ctrl_refillHazards | (((! toplevel_execute_ctrl4_down_LsuL1_HAZARD_lane0) && (LsuL1Plugin_logic_ls_ctrl_askRefill || LsuL1Plugin_logic_ls_ctrl_askUpgrade)) ? (LsuL1Plugin_logic_refill_full ? 1'b1 : LsuL1Plugin_logic_refill_free) : 1'b0));
  assign toplevel_execute_ctrl4_down_LsuL1_WAIT_WRITEBACK_lane0 = 1'b0;
  assign when_LsuL1Plugin_l876 = (toplevel_execute_ctrl4_down_LsuL1_SEL_lane0 && (! toplevel_execute_ctrl4_down_LsuL1_ABORD_lane0));
  assign _zz_38 = {LsuL1Plugin_logic_ls_ctrl_askRefill,{LsuL1Plugin_logic_ls_ctrl_doUpgrade,LsuL1Plugin_logic_ls_ctrl_doFlush}};
  always @(*) begin
    LsuL1Plugin_logic_shared_write_valid = 1'b0;
    if(LsuL1Plugin_logic_ls_ctrl_doFlush) begin
      LsuL1Plugin_logic_shared_write_valid = 1'b1;
    end
    if(LsuL1Plugin_logic_ls_ctrl_doRefill) begin
      LsuL1Plugin_logic_shared_write_valid = 1'b1;
    end
    if(when_LsuL1Plugin_l956) begin
      LsuL1Plugin_logic_shared_write_valid = 1'b1;
    end
    if(LsuL1Plugin_logic_ls_ctrl_preventSideEffects) begin
      LsuL1Plugin_logic_shared_write_valid = 1'b0;
    end
    if(when_LsuL1Plugin_l1160) begin
      LsuL1Plugin_logic_shared_write_valid = 1'b1;
    end
  end

  always @(*) begin
    LsuL1Plugin_logic_shared_write_payload_address = toplevel_execute_ctrl4_down_LsuL1_MIXED_ADDRESS_lane0[11 : 6];
    if(when_LsuL1Plugin_l1160) begin
      LsuL1Plugin_logic_shared_write_payload_address = LsuL1Plugin_logic_initializer_counter[5:0];
    end
  end

  always @(*) begin
    LsuL1Plugin_logic_shared_write_payload_data_plru_0 = LsuL1Plugin_logic_ls_ctrl_plruLogic_core_io_update_state_0;
    if(when_LsuL1Plugin_l1160) begin
      LsuL1Plugin_logic_shared_write_payload_data_plru_0 = _zz_LsuL1Plugin_logic_shared_write_payload_data_plru_0_1[0 : 0];
    end
  end

  always @(*) begin
    LsuL1Plugin_logic_shared_write_payload_data_dirty = ((toplevel_execute_ctrl4_down_LsuL1Plugin_logic_SHARED_lane0_dirty | (LsuL1Plugin_logic_ls_ctrl_doWrite ? toplevel_execute_ctrl4_down_LsuL1Plugin_logic_WAYS_HITS_lane0 : 2'b00)) & (~ ((LsuL1Plugin_logic_ls_ctrl_doRefill ? _zz_LsuL1Plugin_logic_shared_write_payload_data_dirty : 2'b00) | (LsuL1Plugin_logic_ls_ctrl_doFlush ? LsuL1Plugin_logic_ls_ctrl_needFlushOh : 2'b00))));
    if(when_LsuL1Plugin_l1160) begin
      LsuL1Plugin_logic_shared_write_payload_data_dirty = _zz_LsuL1Plugin_logic_shared_write_payload_data_plru_0[2 : 1];
    end
  end

  assign _zz_39 = ({1'd0,1'b1} <<< toplevel_execute_ctrl4_down_LsuL1_PHYSICAL_ADDRESS_lane0[2 : 2]);
  assign when_LsuL1Plugin_l890 = toplevel_execute_ctrl4_down_LsuL1Plugin_logic_WAYS_HITS_lane0[0];
  assign when_LsuL1Plugin_l890_1 = toplevel_execute_ctrl4_down_LsuL1Plugin_logic_WAYS_HITS_lane0[1];
  assign toplevel_execute_ctrl4_down_LsuL1_FLUSH_HIT_lane0 = (|LsuL1Plugin_logic_ls_ctrl_needFlushs);
  assign _zz_LsuL1Plugin_logic_waysWrite_tag_address = _zz__zz_LsuL1Plugin_logic_waysWrite_tag_address;
  assign toplevel_execute_ctrl2_down_LsuL1Plugin_logic_EVENT_WRITE_VALID_lane0 = LsuL1Plugin_logic_ls_ctrl_doWrite;
  assign toplevel_execute_ctrl2_down_LsuL1Plugin_logic_EVENT_WRITE_ADDRESS_lane0 = toplevel_execute_ctrl4_down_LsuL1_PHYSICAL_ADDRESS_lane0;
  assign toplevel_execute_ctrl2_down_LsuL1Plugin_logic_EVENT_WRITE_DATA_lane0 = toplevel_execute_ctrl4_down_LsuL1_WRITE_DATA_lane0;
  assign toplevel_execute_ctrl2_down_LsuL1Plugin_logic_EVENT_WRITE_MASK_lane0 = toplevel_execute_ctrl4_down_LsuL1_MASK_lane0;
  assign when_LsuL1Plugin_l956 = ((toplevel_execute_ctrl4_down_LsuL1_SEL_lane0 && (! toplevel_execute_ctrl4_down_LsuL1_HAZARD_lane0)) && (! toplevel_execute_ctrl4_down_LsuL1_MISS_lane0));
  always @(*) begin
    toplevel_execute_ctrl4_down_LsuL1Plugin_logic_BYPASSED_DATA_lane0 = toplevel_execute_ctrl4_down_LsuL1Plugin_logic_MUXED_DATA_lane0;
    if(when_LsuL1Plugin_l963) begin
      if(when_LsuL1Plugin_l967) begin
        toplevel_execute_ctrl4_down_LsuL1Plugin_logic_BYPASSED_DATA_lane0[7 : 0] = toplevel_execute_ctrl4_down_LsuL1Plugin_logic_EVENT_WRITE_DATA_lane0[7 : 0];
      end
      if(when_LsuL1Plugin_l967_1) begin
        toplevel_execute_ctrl4_down_LsuL1Plugin_logic_BYPASSED_DATA_lane0[15 : 8] = toplevel_execute_ctrl4_down_LsuL1Plugin_logic_EVENT_WRITE_DATA_lane0[15 : 8];
      end
      if(when_LsuL1Plugin_l967_2) begin
        toplevel_execute_ctrl4_down_LsuL1Plugin_logic_BYPASSED_DATA_lane0[23 : 16] = toplevel_execute_ctrl4_down_LsuL1Plugin_logic_EVENT_WRITE_DATA_lane0[23 : 16];
      end
      if(when_LsuL1Plugin_l967_3) begin
        toplevel_execute_ctrl4_down_LsuL1Plugin_logic_BYPASSED_DATA_lane0[31 : 24] = toplevel_execute_ctrl4_down_LsuL1Plugin_logic_EVENT_WRITE_DATA_lane0[31 : 24];
      end
    end
    if(when_LsuL1Plugin_l963_1) begin
      if(when_LsuL1Plugin_l967_4) begin
        toplevel_execute_ctrl4_down_LsuL1Plugin_logic_BYPASSED_DATA_lane0[7 : 0] = toplevel_execute_ctrl3_down_LsuL1Plugin_logic_EVENT_WRITE_DATA_lane0[7 : 0];
      end
      if(when_LsuL1Plugin_l967_5) begin
        toplevel_execute_ctrl4_down_LsuL1Plugin_logic_BYPASSED_DATA_lane0[15 : 8] = toplevel_execute_ctrl3_down_LsuL1Plugin_logic_EVENT_WRITE_DATA_lane0[15 : 8];
      end
      if(when_LsuL1Plugin_l967_6) begin
        toplevel_execute_ctrl4_down_LsuL1Plugin_logic_BYPASSED_DATA_lane0[23 : 16] = toplevel_execute_ctrl3_down_LsuL1Plugin_logic_EVENT_WRITE_DATA_lane0[23 : 16];
      end
      if(when_LsuL1Plugin_l967_7) begin
        toplevel_execute_ctrl4_down_LsuL1Plugin_logic_BYPASSED_DATA_lane0[31 : 24] = toplevel_execute_ctrl3_down_LsuL1Plugin_logic_EVENT_WRITE_DATA_lane0[31 : 24];
      end
    end
  end

  assign when_LsuL1Plugin_l963 = toplevel_execute_ctrl4_down_LsuL1Plugin_logic_WRITE_TO_READ_HAZARDS_lane0[1];
  assign when_LsuL1Plugin_l967 = toplevel_execute_ctrl4_down_LsuL1Plugin_logic_EVENT_WRITE_MASK_lane0[0];
  assign when_LsuL1Plugin_l967_1 = toplevel_execute_ctrl4_down_LsuL1Plugin_logic_EVENT_WRITE_MASK_lane0[1];
  assign when_LsuL1Plugin_l967_2 = toplevel_execute_ctrl4_down_LsuL1Plugin_logic_EVENT_WRITE_MASK_lane0[2];
  assign when_LsuL1Plugin_l967_3 = toplevel_execute_ctrl4_down_LsuL1Plugin_logic_EVENT_WRITE_MASK_lane0[3];
  assign when_LsuL1Plugin_l963_1 = toplevel_execute_ctrl4_down_LsuL1Plugin_logic_WRITE_TO_READ_HAZARDS_lane0[0];
  assign when_LsuL1Plugin_l967_4 = toplevel_execute_ctrl3_down_LsuL1Plugin_logic_EVENT_WRITE_MASK_lane0[0];
  assign when_LsuL1Plugin_l967_5 = toplevel_execute_ctrl3_down_LsuL1Plugin_logic_EVENT_WRITE_MASK_lane0[1];
  assign when_LsuL1Plugin_l967_6 = toplevel_execute_ctrl3_down_LsuL1Plugin_logic_EVENT_WRITE_MASK_lane0[2];
  assign when_LsuL1Plugin_l967_7 = toplevel_execute_ctrl3_down_LsuL1Plugin_logic_EVENT_WRITE_MASK_lane0[3];
  assign toplevel_execute_ctrl4_down_LsuL1_READ_DATA_lane0 = toplevel_execute_ctrl4_down_LsuL1Plugin_logic_BYPASSED_DATA_lane0;
  assign LsuL1Plugin_logic_ls_ctrl_preventSideEffects = (toplevel_execute_ctrl4_down_LsuL1_ABORD_lane0 || execute_freeze_valid);
  assign LsuL1Plugin_logic_initializer_done = LsuL1Plugin_logic_initializer_counter[6];
  assign when_LsuL1Plugin_l1160 = (! LsuL1Plugin_logic_initializer_done);
  assign _zz_LsuL1Plugin_logic_shared_write_payload_data_plru_0 = 3'b000;
  assign LsuL1Plugin_logic_initializerMem_busy = (! LsuL1Plugin_logic_initializerMem_counter[9]);
  assign LsuL1Plugin_logic_refill_read_reservation_win = (! 1'b0);
  assign LsuL1Plugin_logic_ls_ctrl_wayWriteReservation_win = (! (|LsuL1Plugin_logic_refill_read_reservation_take));
  assign LsuL1Plugin_logic_refill_read_writeReservation_win = (! 1'b0);
  assign LsuL1Plugin_logic_ls_ctrl_bankWriteReservation_win = (! (|LsuL1Plugin_logic_refill_read_writeReservation_take));
  always @(*) begin
    LsuPlugin_logic_flusher_arbiter_io_output_ready = 1'b0;
    case(LsuPlugin_logic_flusher_stateReg)
      LsuPlugin_logic_flusher_enumDef_CMD : begin
      end
      LsuPlugin_logic_flusher_enumDef_COMPLETION : begin
        if(when_LsuPlugin_l305) begin
          LsuPlugin_logic_flusher_arbiter_io_output_ready = 1'b1;
        end
      end
      default : begin
      end
    endcase
  end

  assign PrivilegedPlugin_api_lsuTriggerBus_load = toplevel_execute_ctrl3_down_LsuL1_LOAD_lane0;
  assign PrivilegedPlugin_api_lsuTriggerBus_store = toplevel_execute_ctrl3_down_LsuL1_STORE_lane0;
  assign PrivilegedPlugin_api_lsuTriggerBus_virtual = toplevel_execute_ctrl3_down_LsuL1_MIXED_ADDRESS_lane0;
  assign PrivilegedPlugin_api_lsuTriggerBus_size = toplevel_execute_ctrl3_down_LsuL1_SIZE_lane0;
  assign toplevel_execute_ctrl3_down_LsuPlugin_logic_onTrigger_HIT_lane0 = 1'b0;
  assign toplevel_execute_ctrl2_down_LsuPlugin_logic_FORCE_PHYSICAL_lane0 = (toplevel_execute_ctrl2_down_LsuPlugin_logic_FROM_ACCESS_lane0 || toplevel_execute_ctrl2_down_LsuPlugin_logic_FROM_WB_lane0);
  assign LsuPlugin_logic_onAddress0_ls_prefetchOp = toplevel_execute_ctrl2_down_Decode_UOP_lane0[24 : 20];
  assign LsuPlugin_logic_onAddress0_ls_port_valid = (toplevel_execute_ctrl2_up_LANE_SEL_lane0 && toplevel_execute_ctrl2_down_AguPlugin_SEL_lane0);
  assign LsuPlugin_logic_onAddress0_ls_port_payload_address = toplevel_execute_ctrl2_down_early0_SrcPlugin_ADD_SUB_lane0;
  assign LsuPlugin_logic_onAddress0_ls_port_payload_size = toplevel_execute_ctrl2_down_AguPlugin_SIZE_lane0;
  assign LsuPlugin_logic_onAddress0_ls_port_payload_load = toplevel_execute_ctrl2_down_AguPlugin_LOAD_lane0;
  assign LsuPlugin_logic_onAddress0_ls_port_payload_store = toplevel_execute_ctrl2_down_AguPlugin_STORE_lane0;
  assign LsuPlugin_logic_onAddress0_ls_port_payload_atomic = toplevel_execute_ctrl2_down_AguPlugin_ATOMIC_lane0;
  assign LsuPlugin_logic_onAddress0_ls_port_payload_op = LsuL1CmdOpcode_LSU;
  assign LsuPlugin_logic_onAddress0_ls_port_fire = (LsuPlugin_logic_onAddress0_ls_port_valid && LsuPlugin_logic_onAddress0_ls_port_ready);
  assign LsuPlugin_logic_onAddress0_ls_port_payload_storeId = LsuPlugin_logic_onAddress0_ls_storeId;
  assign when_LsuPlugin_l200 = (|(LsuPlugin_logic_onAddress0_access_waiter_refill & (~ LsuL1_REFILL_BUSY)));
  assign LsuPlugin_logic_onAddress0_access_sbWaiter = 1'b0;
  assign _zz_MmuPlugin_logic_accessBus_cmd_ready = (! (LsuPlugin_logic_onAddress0_access_waiter_valid || LsuPlugin_logic_onAddress0_access_sbWaiter));
  assign MmuPlugin_logic_accessBus_cmd_ready = (LsuPlugin_logic_onAddress0_access_port_ready && _zz_MmuPlugin_logic_accessBus_cmd_ready);
  assign LsuPlugin_logic_onAddress0_access_port_valid = (MmuPlugin_logic_accessBus_cmd_valid && _zz_MmuPlugin_logic_accessBus_cmd_ready);
  assign LsuPlugin_logic_onAddress0_access_port_payload_address = MmuPlugin_logic_accessBus_cmd_payload_address;
  assign LsuPlugin_logic_onAddress0_access_port_payload_size = MmuPlugin_logic_accessBus_cmd_payload_size;
  assign LsuPlugin_logic_onAddress0_access_port_payload_load = 1'b1;
  assign LsuPlugin_logic_onAddress0_access_port_payload_store = 1'b0;
  assign LsuPlugin_logic_onAddress0_access_port_payload_atomic = 1'b0;
  assign LsuPlugin_logic_onAddress0_access_port_payload_op = LsuL1CmdOpcode_ACCESS_1;
  assign LsuPlugin_logic_onAddress0_access_port_payload_storeId = 12'h0;
  assign LsuPlugin_logic_onAddress0_flush_port_valid = ((LsuPlugin_logic_flusher_stateReg == LsuPlugin_logic_flusher_enumDef_CMD) && (! LsuPlugin_logic_flusher_cmdCounter[6]));
  assign LsuPlugin_logic_onAddress0_flush_port_payload_address = {19'd0, _zz_LsuPlugin_logic_onAddress0_flush_port_payload_address};
  assign LsuPlugin_logic_onAddress0_flush_port_payload_size = 2'b00;
  assign LsuPlugin_logic_onAddress0_flush_port_payload_load = 1'b0;
  assign LsuPlugin_logic_onAddress0_flush_port_payload_store = 1'b0;
  assign LsuPlugin_logic_onAddress0_flush_port_payload_atomic = 1'b0;
  assign LsuPlugin_logic_onAddress0_flush_port_payload_op = LsuL1CmdOpcode_FLUSH;
  assign LsuPlugin_logic_onAddress0_flush_port_payload_storeId = 12'h0;
  assign LsuPlugin_logic_onAddress0_flush_port_fire = (LsuPlugin_logic_onAddress0_flush_port_valid && LsuPlugin_logic_onAddress0_flush_port_ready);
  assign LsuPlugin_logic_onAddress0_ls_port_ready = LsuPlugin_logic_onAddress0_arbiter_io_inputs_0_ready;
  assign LsuPlugin_logic_onAddress0_access_port_ready = LsuPlugin_logic_onAddress0_arbiter_io_inputs_1_ready;
  assign LsuPlugin_logic_onAddress0_flush_port_ready = LsuPlugin_logic_onAddress0_arbiter_io_inputs_2_ready;
  assign LsuPlugin_logic_onAddress0_arbiter_io_output_ready = (! execute_freeze_valid);
  assign toplevel_execute_ctrl2_down_LsuL1_SEL_lane0 = LsuPlugin_logic_onAddress0_arbiter_io_output_valid;
  assign toplevel_execute_ctrl2_down_LsuL1_MIXED_ADDRESS_lane0 = LsuPlugin_logic_onAddress0_arbiter_io_output_payload_address;
  always @(*) begin
    _zz_toplevel_execute_ctrl2_down_LsuL1_MASK_lane0 = 4'bxxxx;
    case(LsuPlugin_logic_onAddress0_arbiter_io_output_payload_size)
      2'b00 : begin
        _zz_toplevel_execute_ctrl2_down_LsuL1_MASK_lane0 = 4'b0001;
      end
      2'b01 : begin
        _zz_toplevel_execute_ctrl2_down_LsuL1_MASK_lane0 = 4'b0011;
      end
      2'b10 : begin
        _zz_toplevel_execute_ctrl2_down_LsuL1_MASK_lane0 = 4'b1111;
      end
      default : begin
      end
    endcase
  end

  assign toplevel_execute_ctrl2_down_LsuL1_MASK_lane0 = (_zz_toplevel_execute_ctrl2_down_LsuL1_MASK_lane0 <<< LsuPlugin_logic_onAddress0_arbiter_io_output_payload_address[1 : 0]);
  assign toplevel_execute_ctrl2_down_LsuL1_SIZE_lane0 = LsuPlugin_logic_onAddress0_arbiter_io_output_payload_size;
  assign toplevel_execute_ctrl2_down_LsuL1_LOAD_lane0 = LsuPlugin_logic_onAddress0_arbiter_io_output_payload_load;
  assign toplevel_execute_ctrl2_down_LsuL1_ATOMIC_lane0 = LsuPlugin_logic_onAddress0_arbiter_io_output_payload_atomic;
  assign toplevel_execute_ctrl2_down_LsuL1_STORE_lane0 = LsuPlugin_logic_onAddress0_arbiter_io_output_payload_store;
  assign toplevel_execute_ctrl2_down_LsuL1_PREFETCH_lane0 = (LsuPlugin_logic_onAddress0_arbiter_io_output_payload_op == LsuL1CmdOpcode_PREFETCH);
  assign toplevel_execute_ctrl2_down_LsuL1_FLUSH_lane0 = (LsuPlugin_logic_onAddress0_arbiter_io_output_payload_op == LsuL1CmdOpcode_FLUSH);
  assign toplevel_execute_ctrl2_down_Decode_STORE_ID_lane0 = LsuPlugin_logic_onAddress0_arbiter_io_output_payload_storeId;
  assign toplevel_execute_ctrl2_down_LsuPlugin_logic_FROM_ACCESS_lane0 = (LsuPlugin_logic_onAddress0_arbiter_io_output_payload_op == LsuL1CmdOpcode_ACCESS_1);
  assign toplevel_execute_ctrl2_down_LsuPlugin_logic_FROM_WB_lane0 = (LsuPlugin_logic_onAddress0_arbiter_io_output_payload_op == LsuL1CmdOpcode_STORE_BUFFER);
  assign toplevel_execute_ctrl2_down_LsuPlugin_logic_FROM_LSU_lane0 = (LsuPlugin_logic_onAddress0_arbiter_io_output_payload_op == LsuL1CmdOpcode_LSU);
  assign toplevel_execute_ctrl2_down_LsuPlugin_logic_FROM_PREFETCH_lane0 = (LsuPlugin_logic_onAddress0_arbiter_io_output_payload_op == LsuL1CmdOpcode_PREFETCH);
  assign toplevel_execute_ctrl3_down_LsuL1_PHYSICAL_ADDRESS_lane0 = toplevel_execute_ctrl3_down_MMU_TRANSLATED_lane0;
  assign when_LsuPlugin_l449 = (toplevel_execute_ctrl3_down_LsuPlugin_logic_FROM_LSU_lane0 && (! toplevel_execute_ctrl3_up_LANE_SEL_lane0));
  assign when_LsuPlugin_l449_1 = (toplevel_execute_ctrl4_down_LsuPlugin_logic_FROM_LSU_lane0 && (! toplevel_execute_ctrl4_up_LANE_SEL_lane0));
  assign toplevel_execute_ctrl3_down_LsuPlugin_logic_preCtrl_MISS_ALIGNED_lane0 = (|{((toplevel_execute_ctrl3_down_LsuL1_SIZE_lane0 == 2'b10) && (toplevel_execute_ctrl3_down_LsuL1_MIXED_ADDRESS_lane0[1 : 0] != 2'b00)),((toplevel_execute_ctrl3_down_LsuL1_SIZE_lane0 == 2'b01) && (toplevel_execute_ctrl3_down_LsuL1_MIXED_ADDRESS_lane0[0 : 0] != 1'b0))});
  assign toplevel_execute_ctrl3_down_LsuPlugin_logic_preCtrl_IS_AMO_lane0 = (((toplevel_execute_ctrl3_down_AguPlugin_SEL_lane0 && toplevel_execute_ctrl3_down_LsuL1_ATOMIC_lane0) && toplevel_execute_ctrl3_down_LsuL1_STORE_lane0) && toplevel_execute_ctrl3_down_LsuL1_LOAD_lane0);
  assign LsuPlugin_logic_onPma_cached_cmd_address = toplevel_execute_ctrl3_down_MMU_TRANSLATED_lane0;
  assign LsuPlugin_logic_onPma_cached_cmd_op[0] = toplevel_execute_ctrl3_down_LsuL1_STORE_lane0;
  assign LsuPlugin_logic_onPma_io_cmd_address = toplevel_execute_ctrl3_down_MMU_TRANSLATED_lane0;
  assign LsuPlugin_logic_onPma_io_cmd_size = toplevel_execute_ctrl3_down_LsuL1_SIZE_lane0;
  assign LsuPlugin_logic_onPma_io_cmd_op[0] = toplevel_execute_ctrl3_down_LsuL1_STORE_lane0;
  assign toplevel_execute_ctrl3_down_LsuPlugin_logic_onPma_CACHED_RSP_lane0_fault = LsuPlugin_logic_onPma_cached_rsp_fault;
  assign toplevel_execute_ctrl3_down_LsuPlugin_logic_onPma_CACHED_RSP_lane0_io = LsuPlugin_logic_onPma_cached_rsp_io;
  assign toplevel_execute_ctrl3_down_LsuPlugin_logic_onPma_IO_RSP_lane0_fault = LsuPlugin_logic_onPma_io_rsp_fault;
  assign toplevel_execute_ctrl3_down_LsuPlugin_logic_onPma_IO_RSP_lane0_io = LsuPlugin_logic_onPma_io_rsp_io;
  assign toplevel_execute_ctrl3_down_LsuPlugin_logic_onPma_IO_lane0 = (((toplevel_execute_ctrl3_down_LsuPlugin_logic_onPma_CACHED_RSP_lane0_fault && (! toplevel_execute_ctrl3_down_LsuPlugin_logic_onPma_IO_RSP_lane0_fault)) && (! toplevel_execute_ctrl3_down_LsuPlugin_logic_FENCE_lane0)) && (! toplevel_execute_ctrl3_down_LsuPlugin_logic_FROM_PREFETCH_lane0));
  assign LsuPlugin_logic_onPma_addressExtension = (MmuPlugin_api_lsuTranslationEnable ? _zz_LsuPlugin_logic_onPma_addressExtension[31] : 1'b0);
  assign toplevel_execute_ctrl3_down_LsuPlugin_logic_onPma_FROM_LSU_MSB_FAILED_lane0 = (toplevel_execute_ctrl3_down_LsuPlugin_logic_FROM_LSU_lane0 && 1'b0);
  assign toplevel_execute_ctrl3_down_LsuPlugin_logic_MMU_PAGE_FAULT_lane0 = (toplevel_execute_ctrl3_down_MMU_PAGE_FAULT_lane0 || (toplevel_execute_ctrl3_down_AguPlugin_STORE_lane0 ? (! toplevel_execute_ctrl3_down_MMU_ALLOW_WRITE_lane0) : (! toplevel_execute_ctrl3_down_MMU_ALLOW_READ_lane0)));
  assign toplevel_execute_ctrl3_down_LsuPlugin_logic_MMU_FAILURE_lane0 = ((((toplevel_execute_ctrl3_down_LsuPlugin_logic_MMU_PAGE_FAULT_lane0 || toplevel_execute_ctrl3_down_MMU_ACCESS_FAULT_lane0) || toplevel_execute_ctrl3_down_MMU_REFILL_lane0) || toplevel_execute_ctrl3_down_MMU_HAZARD_lane0) || toplevel_execute_ctrl3_down_LsuPlugin_logic_onPma_FROM_LSU_MSB_FAILED_lane0);
  always @(*) begin
    LsuPlugin_logic_onCtrl_lsuTrap = 1'b0;
    if(LsuPlugin_logic_onCtrl_traps_accessFault) begin
      LsuPlugin_logic_onCtrl_lsuTrap = 1'b1;
    end
    if(LsuPlugin_logic_onCtrl_traps_l1Failed) begin
      LsuPlugin_logic_onCtrl_lsuTrap = 1'b1;
    end
    if(LsuPlugin_logic_onCtrl_traps_pmaFault) begin
      LsuPlugin_logic_onCtrl_lsuTrap = 1'b1;
    end
    if(toplevel_execute_ctrl4_down_LsuPlugin_logic_MMU_PAGE_FAULT_lane0) begin
      LsuPlugin_logic_onCtrl_lsuTrap = 1'b1;
    end
    if(toplevel_execute_ctrl4_down_MMU_ACCESS_FAULT_lane0) begin
      LsuPlugin_logic_onCtrl_lsuTrap = 1'b1;
    end
    if(toplevel_execute_ctrl4_down_MMU_REFILL_lane0) begin
      LsuPlugin_logic_onCtrl_lsuTrap = 1'b1;
    end
    if(toplevel_execute_ctrl4_down_MMU_HAZARD_lane0) begin
      LsuPlugin_logic_onCtrl_lsuTrap = 1'b1;
    end
    if(toplevel_execute_ctrl4_down_LsuPlugin_logic_onPma_FROM_LSU_MSB_FAILED_lane0) begin
      LsuPlugin_logic_onCtrl_lsuTrap = 1'b1;
    end
    if(toplevel_execute_ctrl4_down_LsuPlugin_logic_preCtrl_MISS_ALIGNED_lane0) begin
      LsuPlugin_logic_onCtrl_lsuTrap = 1'b1;
    end
    if(toplevel_execute_ctrl4_down_LsuPlugin_logic_onTrigger_HIT_lane0) begin
      LsuPlugin_logic_onCtrl_lsuTrap = 1'b1;
    end
    if(when_LsuPlugin_l710) begin
      LsuPlugin_logic_onCtrl_lsuTrap = 1'b0;
    end
  end

  always @(*) begin
    LsuPlugin_logic_onCtrl_writeData = 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
    LsuPlugin_logic_onCtrl_writeData[31 : 0] = toplevel_execute_ctrl4_up_integer_RS2_lane0;
    if(toplevel_execute_ctrl4_down_LsuPlugin_logic_preCtrl_IS_AMO_lane0) begin
      LsuPlugin_logic_onCtrl_writeData[31 : 0] = LsuPlugin_logic_onCtrl_rva_aluBuffer;
    end
  end

  assign when_LsuPlugin_l491 = ((! LsuPlugin_logic_onCtrl_lsuTrap) && (! toplevel_execute_lane0_ctrls_4_upIsCancel));
  assign LsuPlugin_logic_onCtrl_io_doIt = ((toplevel_execute_ctrl4_up_LANE_SEL_lane0 && toplevel_execute_ctrl4_down_LsuL1_SEL_lane0) && toplevel_execute_ctrl4_down_LsuPlugin_logic_onPma_IO_lane0);
  assign LsuPlugin_logic_bus_cmd_fire = (LsuPlugin_logic_bus_cmd_valid && LsuPlugin_logic_bus_cmd_ready);
  assign when_LsuPlugin_l495 = (! execute_freeze_valid);
  assign LsuPlugin_logic_bus_cmd_valid = (((LsuPlugin_logic_onCtrl_io_doItReg && (! LsuPlugin_logic_onCtrl_io_cmdSent)) && LsuPlugin_logic_onCtrl_io_allowIt) && (! LsuPlugin_logic_onCtrl_io_tooEarly));
  assign LsuPlugin_logic_bus_cmd_payload_write = toplevel_execute_ctrl4_down_LsuL1_STORE_lane0;
  assign LsuPlugin_logic_bus_cmd_payload_address = toplevel_execute_ctrl4_down_LsuL1_PHYSICAL_ADDRESS_lane0;
  assign LsuPlugin_logic_bus_cmd_payload_data = toplevel_execute_ctrl4_down_LsuL1_WRITE_DATA_lane0;
  assign LsuPlugin_logic_bus_cmd_payload_size = toplevel_execute_ctrl4_down_LsuL1_SIZE_lane0;
  assign LsuPlugin_logic_bus_cmd_payload_mask = toplevel_execute_ctrl4_down_LsuL1_MASK_lane0;
  assign LsuPlugin_logic_bus_cmd_payload_io = 1'b1;
  assign LsuPlugin_logic_bus_cmd_payload_fromHart = 1'b1;
  assign LsuPlugin_logic_bus_cmd_payload_uopId = toplevel_execute_ctrl4_down_Decode_UOP_ID_lane0;
  assign LsuPlugin_logic_bus_rsp_toStream_valid = LsuPlugin_logic_bus_rsp_valid;
  assign LsuPlugin_logic_bus_rsp_toStream_payload_error = LsuPlugin_logic_bus_rsp_payload_error;
  assign LsuPlugin_logic_bus_rsp_toStream_payload_data = LsuPlugin_logic_bus_rsp_payload_data;
  assign LsuPlugin_logic_onCtrl_io_rsp_fire = (LsuPlugin_logic_onCtrl_io_rsp_valid && LsuPlugin_logic_onCtrl_io_rsp_ready);
  assign LsuPlugin_logic_bus_rsp_toStream_ready = (! LsuPlugin_logic_bus_rsp_toStream_rValid);
  assign LsuPlugin_logic_onCtrl_io_rsp_valid = LsuPlugin_logic_bus_rsp_toStream_rValid;
  assign LsuPlugin_logic_onCtrl_io_rsp_payload_error = LsuPlugin_logic_bus_rsp_toStream_rData_error;
  assign LsuPlugin_logic_onCtrl_io_rsp_payload_data = LsuPlugin_logic_bus_rsp_toStream_rData_data;
  assign LsuPlugin_logic_onCtrl_io_rsp_ready = (! execute_freeze_valid);
  assign LsuPlugin_logic_onCtrl_io_freezeIt = (LsuPlugin_logic_onCtrl_io_doIt && (LsuPlugin_logic_onCtrl_io_tooEarly || ((! LsuPlugin_logic_onCtrl_io_rsp_valid) && LsuPlugin_logic_onCtrl_io_allowIt)));
  assign LsuPlugin_logic_onCtrl_loadData_input = (LsuPlugin_logic_onCtrl_io_cmdSent ? LsuPlugin_logic_onCtrl_io_rsp_payload_data : toplevel_execute_ctrl4_down_LsuL1_READ_DATA_lane0);
  assign LsuPlugin_logic_onCtrl_loadData_splited_0 = LsuPlugin_logic_onCtrl_loadData_input[7 : 0];
  assign LsuPlugin_logic_onCtrl_loadData_splited_1 = LsuPlugin_logic_onCtrl_loadData_input[15 : 8];
  assign LsuPlugin_logic_onCtrl_loadData_splited_2 = LsuPlugin_logic_onCtrl_loadData_input[23 : 16];
  assign LsuPlugin_logic_onCtrl_loadData_splited_3 = LsuPlugin_logic_onCtrl_loadData_input[31 : 24];
  always @(*) begin
    LsuPlugin_logic_onCtrl_loadData_shited[7 : 0] = _zz_LsuPlugin_logic_onCtrl_loadData_shited;
    LsuPlugin_logic_onCtrl_loadData_shited[15 : 8] = _zz_LsuPlugin_logic_onCtrl_loadData_shited_2;
    LsuPlugin_logic_onCtrl_loadData_shited[23 : 16] = LsuPlugin_logic_onCtrl_loadData_splited_2;
    LsuPlugin_logic_onCtrl_loadData_shited[31 : 24] = LsuPlugin_logic_onCtrl_loadData_splited_3;
  end

  assign toplevel_execute_ctrl4_down_LsuPlugin_logic_onCtrl_loadData_RESULT_lane0 = LsuPlugin_logic_onCtrl_loadData_shited;
  assign LsuPlugin_logic_onCtrl_storeData_mapping_0_1 = {4{LsuPlugin_logic_onCtrl_writeData[7 : 0]}};
  assign LsuPlugin_logic_onCtrl_storeData_mapping_1_1 = {2{LsuPlugin_logic_onCtrl_writeData[15 : 0]}};
  assign LsuPlugin_logic_onCtrl_storeData_mapping_2_1 = {1{LsuPlugin_logic_onCtrl_writeData[31 : 0]}};
  always @(*) begin
    _zz_toplevel_execute_ctrl4_down_LsuL1_WRITE_DATA_lane0 = 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
    case(toplevel_execute_ctrl4_down_LsuL1_SIZE_lane0)
      2'b00 : begin
        _zz_toplevel_execute_ctrl4_down_LsuL1_WRITE_DATA_lane0 = LsuPlugin_logic_onCtrl_storeData_mapping_0_1;
      end
      2'b01 : begin
        _zz_toplevel_execute_ctrl4_down_LsuL1_WRITE_DATA_lane0 = LsuPlugin_logic_onCtrl_storeData_mapping_1_1;
      end
      2'b10 : begin
        _zz_toplevel_execute_ctrl4_down_LsuL1_WRITE_DATA_lane0 = LsuPlugin_logic_onCtrl_storeData_mapping_2_1;
      end
      default : begin
      end
    endcase
  end

  assign toplevel_execute_ctrl4_down_LsuL1_WRITE_DATA_lane0 = _zz_toplevel_execute_ctrl4_down_LsuL1_WRITE_DATA_lane0;
  assign toplevel_execute_ctrl4_down_LsuPlugin_logic_onCtrl_SC_MISS_lane0 = LsuPlugin_logic_onCtrl_scMiss;
  assign _zz_LsuPlugin_logic_onCtrl_rva_alu_compare = toplevel_execute_ctrl4_down_Decode_UOP_lane0[31 : 29];
  assign _zz_LsuPlugin_logic_onCtrl_rva_alu_selectRf = toplevel_execute_ctrl4_down_Decode_UOP_lane0[27];
  assign LsuPlugin_logic_onCtrl_rva_alu_compare = _zz_LsuPlugin_logic_onCtrl_rva_alu_compare[2];
  assign LsuPlugin_logic_onCtrl_rva_alu_unsigned = _zz_LsuPlugin_logic_onCtrl_rva_alu_compare[1];
  assign LsuPlugin_logic_onCtrl_rva_alu_addSub = _zz_LsuPlugin_logic_onCtrl_rva_alu_addSub;
  assign LsuPlugin_logic_onCtrl_rva_alu_less = ((toplevel_execute_ctrl4_down_integer_RS2_lane0[31] == LsuPlugin_logic_onCtrl_rva_srcBuffer[31]) ? LsuPlugin_logic_onCtrl_rva_alu_addSub[31] : (LsuPlugin_logic_onCtrl_rva_alu_unsigned ? LsuPlugin_logic_onCtrl_rva_srcBuffer[31] : toplevel_execute_ctrl4_down_integer_RS2_lane0[31]));
  assign LsuPlugin_logic_onCtrl_rva_alu_selectRf = (_zz_LsuPlugin_logic_onCtrl_rva_alu_selectRf ? 1'b1 : (_zz_LsuPlugin_logic_onCtrl_rva_alu_compare[0] ^ LsuPlugin_logic_onCtrl_rva_alu_less));
  assign switch_Misc_l241_4 = (_zz_LsuPlugin_logic_onCtrl_rva_alu_compare | {_zz_LsuPlugin_logic_onCtrl_rva_alu_selectRf,2'b00});
  always @(*) begin
    case(switch_Misc_l241_4)
      3'b000 : begin
        LsuPlugin_logic_onCtrl_rva_alu_raw = LsuPlugin_logic_onCtrl_rva_alu_addSub;
      end
      3'b001 : begin
        LsuPlugin_logic_onCtrl_rva_alu_raw = (toplevel_execute_ctrl4_down_integer_RS2_lane0 ^ LsuPlugin_logic_onCtrl_rva_srcBuffer);
      end
      3'b010 : begin
        LsuPlugin_logic_onCtrl_rva_alu_raw = (toplevel_execute_ctrl4_down_integer_RS2_lane0 | LsuPlugin_logic_onCtrl_rva_srcBuffer);
      end
      3'b011 : begin
        LsuPlugin_logic_onCtrl_rva_alu_raw = (toplevel_execute_ctrl4_down_integer_RS2_lane0 & LsuPlugin_logic_onCtrl_rva_srcBuffer);
      end
      default : begin
        LsuPlugin_logic_onCtrl_rva_alu_raw = (LsuPlugin_logic_onCtrl_rva_alu_selectRf ? toplevel_execute_ctrl4_down_integer_RS2_lane0 : LsuPlugin_logic_onCtrl_rva_srcBuffer);
      end
    endcase
  end

  assign LsuPlugin_logic_onCtrl_rva_alu_result = LsuPlugin_logic_onCtrl_rva_alu_raw;
  assign LsuPlugin_logic_onCtrl_rva_delay_0 = _zz_LsuPlugin_logic_onCtrl_rva_delay_0;
  assign LsuPlugin_logic_onCtrl_rva_delay_1 = _zz_LsuPlugin_logic_onCtrl_rva_delay_1;
  assign LsuPlugin_logic_onCtrl_rva_freezeIt = ((toplevel_execute_ctrl4_up_LANE_SEL_lane0 && toplevel_execute_ctrl4_down_LsuPlugin_logic_preCtrl_IS_AMO_lane0) && (|{LsuPlugin_logic_onCtrl_rva_delay_1,LsuPlugin_logic_onCtrl_rva_delay_0}));
  always @(*) begin
    LsuPlugin_logic_onCtrl_rva_nc_capture = 1'b0;
    if(when_LsuPlugin_l573) begin
      if(!toplevel_execute_ctrl4_down_LsuL1_STORE_lane0) begin
        if(toplevel_execute_ctrl4_down_LsuL1_ATOMIC_lane0) begin
          LsuPlugin_logic_onCtrl_rva_nc_capture = 1'b1;
        end
      end
    end
  end

  assign when_LsuPlugin_l573 = ((((((! execute_freeze_valid) && toplevel_execute_ctrl4_up_LANE_SEL_lane0) && toplevel_execute_ctrl4_down_LsuPlugin_logic_FROM_LSU_lane0) && toplevel_execute_ctrl4_down_LsuL1_SEL_lane0) && (! LsuPlugin_logic_onCtrl_lsuTrap)) && (! toplevel_execute_ctrl4_down_LsuPlugin_logic_onPma_IO_lane0));
  assign LsuPlugin_logic_onCtrl_scMiss = (! LsuPlugin_logic_onCtrl_rva_nc_reserved);
  assign LsuL1_lockPort_valid = LsuPlugin_logic_onCtrl_rva_nc_reserved;
  assign LsuL1_lockPort_address = LsuPlugin_logic_onCtrl_rva_nc_address;
  assign when_LsuPlugin_l585 = (LsuPlugin_logic_onCtrl_rva_nc_age[5] || LsuPlugin_logic_onCtrl_io_cmdSent);
  always @(*) begin
    LsuPlugin_logic_flushPort_valid = 1'b0;
    if(when_LsuPlugin_l723) begin
      if(LsuPlugin_logic_onCtrl_lsuTrap) begin
        LsuPlugin_logic_flushPort_valid = 1'b1;
      end
    end
  end

  assign LsuPlugin_logic_flushPort_payload_uopId = toplevel_execute_ctrl4_down_Decode_UOP_ID_lane0;
  assign LsuPlugin_logic_flushPort_payload_laneAge = toplevel_execute_ctrl4_down_LANE_AGE_lane0;
  assign LsuPlugin_logic_flushPort_payload_self = 1'b0;
  always @(*) begin
    LsuPlugin_logic_trapPort_valid = 1'b0;
    if(when_LsuPlugin_l723) begin
      if(LsuPlugin_logic_onCtrl_lsuTrap) begin
        LsuPlugin_logic_trapPort_valid = 1'b1;
      end
    end
  end

  assign LsuPlugin_logic_trapPort_payload_laneAge = toplevel_execute_ctrl4_down_LANE_AGE_lane0;
  assign LsuPlugin_logic_trapPort_payload_tval = toplevel_execute_ctrl4_down_LsuL1_MIXED_ADDRESS_lane0;
  always @(*) begin
    LsuPlugin_logic_trapPort_payload_exception = 1'bx;
    if(LsuPlugin_logic_onCtrl_traps_accessFault) begin
      LsuPlugin_logic_trapPort_payload_exception = 1'b1;
    end
    if(LsuPlugin_logic_onCtrl_traps_l1Failed) begin
      LsuPlugin_logic_trapPort_payload_exception = 1'b0;
    end
    if(LsuPlugin_logic_onCtrl_traps_pmaFault) begin
      LsuPlugin_logic_trapPort_payload_exception = 1'b1;
    end
    if(toplevel_execute_ctrl4_down_LsuPlugin_logic_MMU_PAGE_FAULT_lane0) begin
      LsuPlugin_logic_trapPort_payload_exception = 1'b1;
    end
    if(toplevel_execute_ctrl4_down_MMU_ACCESS_FAULT_lane0) begin
      LsuPlugin_logic_trapPort_payload_exception = 1'b1;
    end
    if(toplevel_execute_ctrl4_down_MMU_REFILL_lane0) begin
      LsuPlugin_logic_trapPort_payload_exception = 1'b0;
    end
    if(toplevel_execute_ctrl4_down_MMU_HAZARD_lane0) begin
      LsuPlugin_logic_trapPort_payload_exception = 1'b0;
    end
    if(toplevel_execute_ctrl4_down_LsuPlugin_logic_onPma_FROM_LSU_MSB_FAILED_lane0) begin
      LsuPlugin_logic_trapPort_payload_exception = 1'b1;
    end
    if(toplevel_execute_ctrl4_down_LsuPlugin_logic_preCtrl_MISS_ALIGNED_lane0) begin
      LsuPlugin_logic_trapPort_payload_exception = 1'b1;
    end
    if(toplevel_execute_ctrl4_down_LsuPlugin_logic_onTrigger_HIT_lane0) begin
      LsuPlugin_logic_trapPort_payload_exception = 1'b0;
    end
  end

  always @(*) begin
    LsuPlugin_logic_trapPort_payload_code = 4'bxxxx;
    if(LsuPlugin_logic_onCtrl_traps_accessFault) begin
      LsuPlugin_logic_trapPort_payload_code = 4'b0101;
      if(toplevel_execute_ctrl4_down_AguPlugin_STORE_lane0) begin
        LsuPlugin_logic_trapPort_payload_code[1] = 1'b1;
      end
    end
    if(LsuPlugin_logic_onCtrl_traps_l1Failed) begin
      LsuPlugin_logic_trapPort_payload_code = 4'b0100;
    end
    if(LsuPlugin_logic_onCtrl_traps_pmaFault) begin
      LsuPlugin_logic_trapPort_payload_code = 4'b0101;
      if(toplevel_execute_ctrl4_down_AguPlugin_STORE_lane0) begin
        LsuPlugin_logic_trapPort_payload_code[1] = 1'b1;
      end
    end
    if(toplevel_execute_ctrl4_down_LsuPlugin_logic_MMU_PAGE_FAULT_lane0) begin
      LsuPlugin_logic_trapPort_payload_code = 4'b1101;
      if(toplevel_execute_ctrl4_down_AguPlugin_STORE_lane0) begin
        LsuPlugin_logic_trapPort_payload_code[1] = 1'b1;
      end
    end
    if(toplevel_execute_ctrl4_down_MMU_ACCESS_FAULT_lane0) begin
      LsuPlugin_logic_trapPort_payload_code = 4'b0101;
      if(toplevel_execute_ctrl4_down_AguPlugin_STORE_lane0) begin
        LsuPlugin_logic_trapPort_payload_code[1] = 1'b1;
      end
    end
    if(toplevel_execute_ctrl4_down_MMU_REFILL_lane0) begin
      LsuPlugin_logic_trapPort_payload_code = 4'b0111;
    end
    if(toplevel_execute_ctrl4_down_MMU_HAZARD_lane0) begin
      LsuPlugin_logic_trapPort_payload_code = 4'b0100;
    end
    if(toplevel_execute_ctrl4_down_LsuPlugin_logic_onPma_FROM_LSU_MSB_FAILED_lane0) begin
      LsuPlugin_logic_trapPort_payload_code = 4'b0101;
      if(toplevel_execute_ctrl4_down_AguPlugin_STORE_lane0) begin
        LsuPlugin_logic_trapPort_payload_code[1] = 1'b1;
      end
      if(when_LsuPlugin_l683) begin
        LsuPlugin_logic_trapPort_payload_code[3] = 1'b1;
      end
    end
    if(toplevel_execute_ctrl4_down_LsuPlugin_logic_preCtrl_MISS_ALIGNED_lane0) begin
      LsuPlugin_logic_trapPort_payload_code = {1'd0, _zz_LsuPlugin_logic_trapPort_payload_code};
    end
    if(toplevel_execute_ctrl4_down_LsuPlugin_logic_onTrigger_HIT_lane0) begin
      LsuPlugin_logic_trapPort_payload_code = 4'b0011;
    end
  end

  always @(*) begin
    LsuPlugin_logic_trapPort_payload_arg = 3'b000;
    LsuPlugin_logic_trapPort_payload_arg[1 : 0] = (toplevel_execute_ctrl4_down_AguPlugin_STORE_lane0 ? 2'b01 : 2'b00);
    LsuPlugin_logic_trapPort_payload_arg[2 : 2] = 1'b1;
  end

  assign LsuPlugin_logic_onCtrl_traps_accessFault = (toplevel_execute_ctrl4_down_LsuPlugin_logic_onPma_CACHED_RSP_lane0_fault ? ((LsuPlugin_logic_onCtrl_io_rsp_valid && LsuPlugin_logic_onCtrl_io_rsp_payload_error) || toplevel_execute_ctrl4_down_LsuL1_ATOMIC_lane0) : toplevel_execute_ctrl4_down_LsuL1_FAULT_lane0);
  assign LsuPlugin_logic_onCtrl_traps_l1Failed = ((! toplevel_execute_ctrl4_down_LsuPlugin_logic_onPma_CACHED_RSP_lane0_fault) && ((toplevel_execute_ctrl4_down_LsuL1_HAZARD_lane0 || toplevel_execute_ctrl4_down_LsuL1_MISS_lane0) || toplevel_execute_ctrl4_down_LsuL1_MISS_UNIQUE_lane0));
  assign LsuPlugin_logic_onCtrl_traps_pmaFault = (toplevel_execute_ctrl4_down_LsuPlugin_logic_onPma_CACHED_RSP_lane0_fault && toplevel_execute_ctrl4_down_LsuPlugin_logic_onPma_IO_RSP_lane0_fault);
  assign when_LsuPlugin_l683 = (! toplevel_execute_ctrl4_down_MMU_BYPASS_TRANSLATION_lane0);
  assign when_LsuPlugin_l710 = (toplevel_execute_ctrl4_down_LsuPlugin_logic_FENCE_lane0 || toplevel_execute_ctrl4_down_LsuPlugin_logic_FROM_PREFETCH_lane0);
  assign when_LsuPlugin_l723 = (toplevel_execute_ctrl4_up_LANE_SEL_lane0 && toplevel_execute_ctrl4_down_AguPlugin_SEL_lane0);
  assign LsuPlugin_logic_onCtrl_mmuNeeded = (toplevel_execute_ctrl4_down_LsuPlugin_logic_FROM_LSU_lane0 || toplevel_execute_ctrl4_down_LsuPlugin_logic_FROM_PREFETCH_lane0);
  assign toplevel_execute_ctrl4_down_LsuL1_ABORD_lane0 = (|{(LsuPlugin_logic_onCtrl_mmuNeeded && toplevel_execute_ctrl4_down_LsuPlugin_logic_MMU_FAILURE_lane0),{(toplevel_execute_ctrl4_down_LsuPlugin_logic_FROM_LSU_lane0 && ((! toplevel_execute_ctrl4_up_LANE_SEL_lane0) || toplevel_execute_lane0_ctrls_4_upIsCancel)),{((! toplevel_execute_ctrl4_down_LsuL1_FLUSH_lane0) && toplevel_execute_ctrl4_down_LsuPlugin_logic_onPma_CACHED_RSP_lane0_fault),{toplevel_execute_ctrl4_down_LsuL1_FLUSH_HAZARD_lane0,toplevel_execute_ctrl4_down_LsuL1_HAZARD_lane0}}}});
  assign toplevel_execute_ctrl4_down_LsuL1_SKIP_WRITE_lane0 = (|{((toplevel_execute_ctrl4_down_LsuL1_ATOMIC_lane0 && (! toplevel_execute_ctrl4_down_LsuL1_LOAD_lane0)) && LsuPlugin_logic_onCtrl_scMiss),{toplevel_execute_ctrl4_down_LsuPlugin_logic_FROM_PREFETCH_lane0,{(toplevel_execute_ctrl4_down_LsuPlugin_logic_FROM_LSU_lane0 && toplevel_execute_ctrl4_down_LsuPlugin_logic_onTrigger_HIT_lane0),{toplevel_execute_ctrl4_down_LsuPlugin_logic_preCtrl_MISS_ALIGNED_lane0,{toplevel_execute_ctrl4_down_LsuL1_FAULT_lane0,(toplevel_execute_ctrl4_down_LsuL1_MISS_lane0 || toplevel_execute_ctrl4_down_LsuL1_MISS_UNIQUE_lane0)}}}}});
  assign when_LsuPlugin_l761 = ((toplevel_execute_ctrl4_down_LsuL1_SEL_lane0 && toplevel_execute_ctrl4_down_LsuL1_FLUSH_lane0) && ((toplevel_execute_ctrl4_down_LsuL1_FLUSH_HIT_lane0 || toplevel_execute_ctrl4_down_LsuL1_HAZARD_lane0) || toplevel_execute_ctrl4_down_LsuL1_FLUSH_HAZARD_lane0));
  assign MmuPlugin_logic_accessBus_rsp_valid = ((toplevel_execute_ctrl4_down_LsuL1_SEL_lane0 && toplevel_execute_ctrl4_down_LsuPlugin_logic_FROM_ACCESS_lane0) && (! execute_freeze_valid));
  assign MmuPlugin_logic_accessBus_rsp_payload_data = toplevel_execute_ctrl4_down_LsuPlugin_logic_onCtrl_loadData_RESULT_lane0;
  always @(*) begin
    MmuPlugin_logic_accessBus_rsp_payload_error = toplevel_execute_ctrl4_down_LsuL1_FAULT_lane0;
    if(LsuPlugin_logic_onCtrl_traps_pmaFault) begin
      MmuPlugin_logic_accessBus_rsp_payload_error = 1'b1;
    end
  end

  always @(*) begin
    MmuPlugin_logic_accessBus_rsp_payload_redo = LsuPlugin_logic_onCtrl_traps_l1Failed;
    if(LsuPlugin_logic_onCtrl_traps_pmaFault) begin
      MmuPlugin_logic_accessBus_rsp_payload_redo = 1'b0;
    end
  end

  assign MmuPlugin_logic_accessBus_rsp_payload_waitAny = 1'b0;
  assign when_LsuPlugin_l796 = (MmuPlugin_logic_accessBus_rsp_valid && MmuPlugin_logic_accessBus_rsp_payload_redo);
  assign when_LsuPlugin_l204 = (|toplevel_execute_ctrl4_down_LsuL1_WAIT_REFILL_lane0);
  assign when_LsuPlugin_l200_1 = (|(LsuPlugin_logic_onCtrl_hartRegulation_refill & (~ LsuL1_REFILL_BUSY)));
  assign when_LsuPlugin_l803 = ((((((toplevel_execute_ctrl4_up_LANE_SEL_lane0 && toplevel_execute_ctrl4_down_AguPlugin_SEL_lane0) && (! toplevel_execute_ctrl4_down_LsuPlugin_logic_FROM_PREFETCH_lane0)) && (! toplevel_execute_ctrl4_down_LsuPlugin_logic_onPma_IO_lane0)) && (! toplevel_execute_ctrl4_down_LsuPlugin_logic_FENCE_lane0)) && 1'b1) && ((toplevel_execute_ctrl4_down_LsuL1_HAZARD_lane0 || toplevel_execute_ctrl4_down_LsuL1_MISS_lane0) || toplevel_execute_ctrl4_down_LsuL1_MISS_UNIQUE_lane0));
  assign when_LsuPlugin_l204_1 = (|toplevel_execute_ctrl4_down_LsuL1_WAIT_REFILL_lane0);
  assign LsuPlugin_logic_commitProbe_valid = (((toplevel_execute_ctrl4_down_LANE_SEL_lane0 && toplevel_execute_ctrl4_down_isReady) && (! toplevel_execute_lane0_ctrls_4_downIsCancel)) && (toplevel_execute_ctrl4_down_AguPlugin_SEL_lane0 ? toplevel_execute_ctrl4_down_LsuPlugin_logic_FROM_LSU_lane0 : (toplevel_execute_ctrl4_down_LsuPlugin_logic_FROM_PREFETCH_lane0 && toplevel_execute_ctrl4_down_LsuL1_HAZARD_lane0)));
  assign LsuPlugin_logic_commitProbe_payload_address = toplevel_execute_ctrl4_down_LsuL1_MIXED_ADDRESS_lane0;
  assign LsuPlugin_logic_commitProbe_payload_load = toplevel_execute_ctrl4_down_LsuL1_LOAD_lane0;
  assign LsuPlugin_logic_commitProbe_payload_store = toplevel_execute_ctrl4_down_LsuL1_STORE_lane0;
  assign LsuPlugin_logic_commitProbe_payload_trap = LsuPlugin_logic_onCtrl_lsuTrap;
  assign LsuPlugin_logic_commitProbe_payload_miss = ((toplevel_execute_ctrl4_down_LsuL1_MISS_lane0 && (! toplevel_execute_ctrl4_down_LsuL1_HAZARD_lane0)) && (! toplevel_execute_ctrl4_down_LsuPlugin_logic_MMU_FAILURE_lane0));
  assign LsuPlugin_logic_commitProbe_payload_io = toplevel_execute_ctrl4_down_LsuPlugin_logic_onPma_IO_lane0;
  assign LsuPlugin_logic_commitProbe_payload_prefetchFailed = toplevel_execute_ctrl4_down_LsuPlugin_logic_FROM_PREFETCH_lane0;
  assign LsuPlugin_logic_commitProbe_payload_pc = toplevel_execute_ctrl4_down_PC_lane0;
  assign LsuPlugin_logic_iwb_valid = (toplevel_execute_ctrl4_down_AguPlugin_SEL_lane0 && (! toplevel_execute_ctrl4_down_AguPlugin_FLOAT_lane0));
  always @(*) begin
    LsuPlugin_logic_iwb_payload = toplevel_execute_ctrl4_down_LsuPlugin_logic_onCtrl_loadData_RESULT_lane0;
    if(when_LsuPlugin_l824) begin
      LsuPlugin_logic_iwb_payload[0] = toplevel_execute_ctrl4_down_LsuPlugin_logic_onCtrl_SC_MISS_lane0;
      LsuPlugin_logic_iwb_payload[7 : 1] = 7'h0;
    end
  end

  assign when_LsuPlugin_l824 = (toplevel_execute_ctrl4_down_LsuL1_ATOMIC_lane0 && (! toplevel_execute_ctrl4_down_LsuL1_LOAD_lane0));
  assign LsuPlugin_logic_onWb_storeFire = ((((((toplevel_execute_ctrl4_down_LANE_SEL_lane0 && toplevel_execute_ctrl4_down_isReady) && (! toplevel_execute_lane0_ctrls_4_downIsCancel)) && toplevel_execute_ctrl4_down_AguPlugin_SEL_lane0) && toplevel_execute_ctrl4_down_AguPlugin_STORE_lane0) && (! toplevel_execute_ctrl4_down_LsuPlugin_logic_onPma_IO_lane0)) && (! toplevel_execute_ctrl4_down_LsuPlugin_logic_FROM_PREFETCH_lane0));
  assign LsuPlugin_logic_onWb_storeBroadcast = (((((((toplevel_execute_ctrl4_down_isReady && toplevel_execute_ctrl4_down_LsuL1_SEL_lane0) && toplevel_execute_ctrl4_down_LsuL1_STORE_lane0) && (! toplevel_execute_ctrl4_down_LsuL1_ABORD_lane0)) && (! toplevel_execute_ctrl4_down_LsuL1_SKIP_WRITE_lane0)) && (! toplevel_execute_ctrl4_down_LsuL1_MISS_lane0)) && (! toplevel_execute_ctrl4_down_LsuL1_MISS_UNIQUE_lane0)) && (! toplevel_execute_ctrl4_down_LsuL1_HAZARD_lane0));
  assign LsuL1TileLinkPlugin_logic_down_a_fire = (LsuL1TileLinkPlugin_logic_down_a_valid && LsuL1TileLinkPlugin_logic_down_a_ready);
  assign LsuL1TileLinkPlugin_logic_down_a_tracker_last = ((! ((1'b0 || (A_PUT_FULL_DATA == LsuL1TileLinkPlugin_logic_down_a_payload_opcode)) || (A_PUT_PARTIAL_DATA == LsuL1TileLinkPlugin_logic_down_a_payload_opcode))) || (LsuL1Plugin_logic_bus_toTilelink_nonCoherent_onA_beat == _zz_LsuL1TileLinkPlugin_logic_down_a_tracker_last));
  assign when_LsuL1Bus_l402 = (LsuL1TileLinkPlugin_logic_down_a_fire && LsuL1TileLinkPlugin_logic_down_a_tracker_last);
  assign LsuL1Plugin_logic_bus_toTilelink_nonCoherent_onA_sel = (LsuL1Plugin_logic_bus_toTilelink_nonCoherent_onA_lock ? LsuL1Plugin_logic_bus_toTilelink_nonCoherent_onA_selReg : LsuL1Plugin_logic_bus_read_cmd_valid);
  assign LsuL1TileLinkPlugin_logic_down_a_payload_param = 3'b000;
  assign LsuL1TileLinkPlugin_logic_down_a_payload_size = 3'b110;
  assign LsuL1TileLinkPlugin_logic_down_a_payload_mask = 8'hff;
  assign LsuL1TileLinkPlugin_logic_down_a_payload_data = LsuL1Plugin_logic_bus_write_cmd_payload_fragment_data;
  assign LsuL1TileLinkPlugin_logic_down_a_payload_corrupt = 1'b0;
  always @(*) begin
    if(LsuL1Plugin_logic_bus_toTilelink_nonCoherent_onA_sel) begin
      LsuL1TileLinkPlugin_logic_down_a_valid = LsuL1Plugin_logic_bus_read_cmd_valid;
    end else begin
      LsuL1TileLinkPlugin_logic_down_a_valid = LsuL1Plugin_logic_bus_write_cmd_valid;
    end
  end

  always @(*) begin
    if(LsuL1Plugin_logic_bus_toTilelink_nonCoherent_onA_sel) begin
      LsuL1TileLinkPlugin_logic_down_a_payload_opcode = A_GET;
    end else begin
      LsuL1TileLinkPlugin_logic_down_a_payload_opcode = A_PUT_FULL_DATA;
    end
  end

  always @(*) begin
    if(LsuL1Plugin_logic_bus_toTilelink_nonCoherent_onA_sel) begin
      LsuL1TileLinkPlugin_logic_down_a_payload_source = 1'b0;
    end else begin
      LsuL1TileLinkPlugin_logic_down_a_payload_source = 1'b0;
    end
    LsuL1TileLinkPlugin_logic_down_a_payload_source[0] = LsuL1Plugin_logic_bus_toTilelink_nonCoherent_onA_sel;
  end

  always @(*) begin
    if(LsuL1Plugin_logic_bus_toTilelink_nonCoherent_onA_sel) begin
      LsuL1TileLinkPlugin_logic_down_a_payload_address = LsuL1Plugin_logic_bus_read_cmd_payload_address;
    end else begin
      LsuL1TileLinkPlugin_logic_down_a_payload_address = LsuL1Plugin_logic_bus_write_cmd_payload_fragment_address;
    end
    LsuL1TileLinkPlugin_logic_down_a_payload_address[5 : 3] = LsuL1Plugin_logic_bus_toTilelink_nonCoherent_onA_beat;
  end

  assign LsuL1Plugin_logic_bus_write_cmd_ready = ((! LsuL1Plugin_logic_bus_toTilelink_nonCoherent_onA_sel) && LsuL1TileLinkPlugin_logic_down_a_ready);
  assign LsuL1Plugin_logic_bus_read_cmd_ready = (LsuL1Plugin_logic_bus_toTilelink_nonCoherent_onA_sel && LsuL1TileLinkPlugin_logic_down_a_ready);
  assign LsuL1Plugin_logic_bus_toTilelink_nonCoherent_onD_sel = LsuL1TileLinkPlugin_logic_down_d_payload_source[0];
  assign LsuL1Plugin_logic_bus_read_rsp_valid = (LsuL1TileLinkPlugin_logic_down_d_valid && LsuL1Plugin_logic_bus_toTilelink_nonCoherent_onD_sel);
  assign LsuL1Plugin_logic_bus_read_rsp_payload_data = LsuL1TileLinkPlugin_logic_down_d_payload_data;
  assign LsuL1Plugin_logic_bus_read_rsp_payload_error = (LsuL1TileLinkPlugin_logic_down_d_payload_denied || LsuL1TileLinkPlugin_logic_down_d_payload_corrupt);
  assign LsuL1Plugin_logic_bus_write_rsp_valid = (LsuL1TileLinkPlugin_logic_down_d_valid && (! LsuL1Plugin_logic_bus_toTilelink_nonCoherent_onD_sel));
  assign LsuL1Plugin_logic_bus_write_rsp_payload_error = (LsuL1TileLinkPlugin_logic_down_d_payload_denied || LsuL1TileLinkPlugin_logic_down_d_payload_corrupt);
  assign LsuL1TileLinkPlugin_logic_down_d_ready = (LsuL1Plugin_logic_bus_toTilelink_nonCoherent_onD_sel ? LsuL1Plugin_logic_bus_read_rsp_ready : 1'b1);
  always @(*) begin
    TrapPlugin_logic_harts_0_crsPorts_write_valid = 1'b0;
    case(TrapPlugin_logic_harts_0_trap_fsm_stateReg)
      TrapPlugin_logic_harts_0_trap_fsm_enumDef_RUNNING : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_enumDef_PROCESS_1 : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_enumDef_TRAP_EPC : begin
        TrapPlugin_logic_harts_0_crsPorts_write_valid = 1'b1;
      end
      TrapPlugin_logic_harts_0_trap_fsm_enumDef_TRAP_TVAL : begin
        TrapPlugin_logic_harts_0_crsPorts_write_valid = 1'b1;
      end
      TrapPlugin_logic_harts_0_trap_fsm_enumDef_TRAP_TVEC : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_enumDef_TRAP_APPLY : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_enumDef_XRET_EPC : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_enumDef_XRET_APPLY : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_enumDef_ATS_RSP : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_enumDef_JUMP : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_enumDef_LSU_FLUSH : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_enumDef_FETCH_FLUSH : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    TrapPlugin_logic_harts_0_crsPorts_write_address = 3'bxxx;
    case(TrapPlugin_logic_harts_0_trap_fsm_stateReg)
      TrapPlugin_logic_harts_0_trap_fsm_enumDef_RUNNING : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_enumDef_PROCESS_1 : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_enumDef_TRAP_EPC : begin
        TrapPlugin_logic_harts_0_crsPorts_write_address = _zz_TrapPlugin_logic_harts_0_crsPorts_write_address;
      end
      TrapPlugin_logic_harts_0_trap_fsm_enumDef_TRAP_TVAL : begin
        TrapPlugin_logic_harts_0_crsPorts_write_address = _zz_TrapPlugin_logic_harts_0_crsPorts_write_address_1;
      end
      TrapPlugin_logic_harts_0_trap_fsm_enumDef_TRAP_TVEC : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_enumDef_TRAP_APPLY : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_enumDef_XRET_EPC : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_enumDef_XRET_APPLY : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_enumDef_ATS_RSP : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_enumDef_JUMP : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_enumDef_LSU_FLUSH : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_enumDef_FETCH_FLUSH : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    TrapPlugin_logic_harts_0_crsPorts_write_data = 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
    case(TrapPlugin_logic_harts_0_trap_fsm_stateReg)
      TrapPlugin_logic_harts_0_trap_fsm_enumDef_RUNNING : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_enumDef_PROCESS_1 : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_enumDef_TRAP_EPC : begin
        TrapPlugin_logic_harts_0_crsPorts_write_data = TrapPlugin_logic_harts_0_trap_pending_pc;
      end
      TrapPlugin_logic_harts_0_trap_fsm_enumDef_TRAP_TVAL : begin
        TrapPlugin_logic_harts_0_crsPorts_write_data = TrapPlugin_logic_harts_0_trap_fsm_buffer_trap_tval;
        if(TrapPlugin_logic_harts_0_trap_fsm_triggerEbreakReg) begin
          TrapPlugin_logic_harts_0_crsPorts_write_data = TrapPlugin_logic_harts_0_trap_pending_pc;
        end
      end
      TrapPlugin_logic_harts_0_trap_fsm_enumDef_TRAP_TVEC : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_enumDef_TRAP_APPLY : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_enumDef_XRET_EPC : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_enumDef_XRET_APPLY : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_enumDef_ATS_RSP : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_enumDef_JUMP : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_enumDef_LSU_FLUSH : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_enumDef_FETCH_FLUSH : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    TrapPlugin_logic_harts_0_interrupt_valid = 1'b0;
    if(when_TrapPlugin_l189_1) begin
      if(when_TrapPlugin_l195) begin
        TrapPlugin_logic_harts_0_interrupt_valid = 1'b1;
      end
      if(when_TrapPlugin_l195_1) begin
        TrapPlugin_logic_harts_0_interrupt_valid = 1'b1;
      end
      if(when_TrapPlugin_l195_2) begin
        TrapPlugin_logic_harts_0_interrupt_valid = 1'b1;
      end
    end
    if(when_TrapPlugin_l189) begin
      if(when_TrapPlugin_l195_3) begin
        TrapPlugin_logic_harts_0_interrupt_valid = 1'b1;
      end
      if(when_TrapPlugin_l195_4) begin
        TrapPlugin_logic_harts_0_interrupt_valid = 1'b1;
      end
      if(when_TrapPlugin_l195_5) begin
        TrapPlugin_logic_harts_0_interrupt_valid = 1'b1;
      end
      if(when_TrapPlugin_l195_6) begin
        TrapPlugin_logic_harts_0_interrupt_valid = 1'b1;
      end
      if(when_TrapPlugin_l195_7) begin
        TrapPlugin_logic_harts_0_interrupt_valid = 1'b1;
      end
      if(when_TrapPlugin_l195_8) begin
        TrapPlugin_logic_harts_0_interrupt_valid = 1'b1;
      end
    end
  end

  always @(*) begin
    TrapPlugin_logic_harts_0_interrupt_code = 4'bxxxx;
    if(when_TrapPlugin_l189_1) begin
      if(when_TrapPlugin_l195) begin
        TrapPlugin_logic_harts_0_interrupt_code = 4'b0001;
      end
      if(when_TrapPlugin_l195_1) begin
        TrapPlugin_logic_harts_0_interrupt_code = 4'b0101;
      end
      if(when_TrapPlugin_l195_2) begin
        TrapPlugin_logic_harts_0_interrupt_code = 4'b1001;
      end
    end
    if(when_TrapPlugin_l189) begin
      if(when_TrapPlugin_l195_3) begin
        TrapPlugin_logic_harts_0_interrupt_code = 4'b0111;
      end
      if(when_TrapPlugin_l195_4) begin
        TrapPlugin_logic_harts_0_interrupt_code = 4'b0011;
      end
      if(when_TrapPlugin_l195_5) begin
        TrapPlugin_logic_harts_0_interrupt_code = 4'b1011;
      end
      if(when_TrapPlugin_l195_6) begin
        TrapPlugin_logic_harts_0_interrupt_code = 4'b0001;
      end
      if(when_TrapPlugin_l195_7) begin
        TrapPlugin_logic_harts_0_interrupt_code = 4'b0101;
      end
      if(when_TrapPlugin_l195_8) begin
        TrapPlugin_logic_harts_0_interrupt_code = 4'b1001;
      end
    end
  end

  always @(*) begin
    TrapPlugin_logic_harts_0_interrupt_targetPrivilege = 2'bxx;
    if(when_TrapPlugin_l189_1) begin
      if(when_TrapPlugin_l195) begin
        TrapPlugin_logic_harts_0_interrupt_targetPrivilege = 2'b01;
      end
      if(when_TrapPlugin_l195_1) begin
        TrapPlugin_logic_harts_0_interrupt_targetPrivilege = 2'b01;
      end
      if(when_TrapPlugin_l195_2) begin
        TrapPlugin_logic_harts_0_interrupt_targetPrivilege = 2'b01;
      end
    end
    if(when_TrapPlugin_l189) begin
      if(when_TrapPlugin_l195_3) begin
        TrapPlugin_logic_harts_0_interrupt_targetPrivilege = 2'b11;
      end
      if(when_TrapPlugin_l195_4) begin
        TrapPlugin_logic_harts_0_interrupt_targetPrivilege = 2'b11;
      end
      if(when_TrapPlugin_l195_5) begin
        TrapPlugin_logic_harts_0_interrupt_targetPrivilege = 2'b11;
      end
      if(when_TrapPlugin_l195_6) begin
        TrapPlugin_logic_harts_0_interrupt_targetPrivilege = 2'b11;
      end
      if(when_TrapPlugin_l195_7) begin
        TrapPlugin_logic_harts_0_interrupt_targetPrivilege = 2'b11;
      end
      if(when_TrapPlugin_l195_8) begin
        TrapPlugin_logic_harts_0_interrupt_targetPrivilege = 2'b11;
      end
    end
  end

  assign when_TrapPlugin_l189 = (PrivilegedPlugin_logic_harts_0_m_status_mie || (! PrivilegedPlugin_logic_harts_0_withMachinePrivilege));
  assign when_TrapPlugin_l189_1 = ((PrivilegedPlugin_logic_harts_0_s_status_sie && (! PrivilegedPlugin_logic_harts_0_withMachinePrivilege)) || (! PrivilegedPlugin_logic_harts_0_withSupervisorPrivilege));
  assign when_TrapPlugin_l195 = ((_zz_when_TrapPlugin_l195_3 && (1'b1 && PrivilegedPlugin_logic_harts_0_m_ideleg_ss)) && (! 1'b0));
  assign when_TrapPlugin_l195_1 = ((_zz_when_TrapPlugin_l195_4 && (1'b1 && PrivilegedPlugin_logic_harts_0_m_ideleg_st)) && (! 1'b0));
  assign when_TrapPlugin_l195_2 = ((_zz_when_TrapPlugin_l195_5 && (1'b1 && PrivilegedPlugin_logic_harts_0_m_ideleg_se)) && (! 1'b0));
  assign when_TrapPlugin_l195_3 = ((_zz_when_TrapPlugin_l195 && 1'b1) && (! 1'b0));
  assign when_TrapPlugin_l195_4 = ((_zz_when_TrapPlugin_l195_1 && 1'b1) && (! 1'b0));
  assign when_TrapPlugin_l195_5 = ((_zz_when_TrapPlugin_l195_2 && 1'b1) && (! 1'b0));
  assign when_TrapPlugin_l195_6 = ((_zz_when_TrapPlugin_l195_3 && 1'b1) && (! (|PrivilegedPlugin_logic_harts_0_m_ideleg_ss)));
  assign when_TrapPlugin_l195_7 = ((_zz_when_TrapPlugin_l195_4 && 1'b1) && (! (|PrivilegedPlugin_logic_harts_0_m_ideleg_st)));
  assign when_TrapPlugin_l195_8 = ((_zz_when_TrapPlugin_l195_5 && 1'b1) && (! (|PrivilegedPlugin_logic_harts_0_m_ideleg_se)));
  assign TrapPlugin_logic_harts_0_interrupt_pendingInterrupt = (TrapPlugin_logic_harts_0_interrupt_validBuffer && PrivilegedPlugin_api_harts_0_allowInterrupts);
  assign when_TrapPlugin_l214 = (|{_zz_when_TrapPlugin_l195_5,{_zz_when_TrapPlugin_l195_4,{_zz_when_TrapPlugin_l195_3,{_zz_when_TrapPlugin_l195_2,{_zz_when_TrapPlugin_l195_1,_zz_when_TrapPlugin_l195}}}}});
  assign _zz_TrapPlugin_logic_harts_0_trap_pending_arbiter_ports_1_valid = (early0_EnvPlugin_logic_trapPort_valid && 1'b1);
  assign _zz_TrapPlugin_logic_harts_0_trap_pending_arbiter_ports_3_valid = (FetchL1Plugin_logic_trapPort_valid && 1'b1);
  assign _zz_TrapPlugin_logic_harts_0_trap_pending_arbiter_ports_0_valid = (LsuPlugin_logic_trapPort_valid && 1'b1);
  assign _zz_TrapPlugin_logic_harts_0_trap_pending_arbiter_ports_1_valid_1 = (CsrAccessPlugin_logic_trapPort_valid && 1'b1);
  assign _zz_TrapPlugin_logic_harts_0_trap_pending_arbiter_ports_2_valid = (DecoderPlugin_logic_laneLogic_0_trapPort_valid && 1'b1);
  assign _zz_TrapPlugin_logic_harts_0_trap_pending_arbiter_ports_2_valid_1 = (DecoderPlugin_logic_laneLogic_1_trapPort_valid && 1'b1);
  assign TrapPlugin_logic_harts_0_trap_pending_arbiter_ports_0_valid = (|_zz_TrapPlugin_logic_harts_0_trap_pending_arbiter_ports_0_valid);
  assign TrapPlugin_logic_harts_0_trap_pending_arbiter_ports_0_payload_exception = LsuPlugin_logic_trapPort_payload_exception;
  assign TrapPlugin_logic_harts_0_trap_pending_arbiter_ports_0_payload_tval = LsuPlugin_logic_trapPort_payload_tval;
  assign TrapPlugin_logic_harts_0_trap_pending_arbiter_ports_0_payload_code = LsuPlugin_logic_trapPort_payload_code;
  assign TrapPlugin_logic_harts_0_trap_pending_arbiter_ports_0_payload_arg = LsuPlugin_logic_trapPort_payload_arg;
  assign _zz_TrapPlugin_logic_harts_0_trap_pending_arbiter_ports_1_payload_exception = {(_zz_TrapPlugin_logic_harts_0_trap_pending_arbiter_ports_1_valid_1 && (&(! (_zz_TrapPlugin_logic_harts_0_trap_pending_arbiter_ports_1_valid && (early0_EnvPlugin_logic_trapPort_payload_laneAge < CsrAccessPlugin_logic_trapPort_payload_laneAge))))),(_zz_TrapPlugin_logic_harts_0_trap_pending_arbiter_ports_1_valid && (&(! (_zz_TrapPlugin_logic_harts_0_trap_pending_arbiter_ports_1_valid_1 && (CsrAccessPlugin_logic_trapPort_payload_laneAge < early0_EnvPlugin_logic_trapPort_payload_laneAge)))))};
  assign TrapPlugin_logic_harts_0_trap_pending_arbiter_ports_1_valid = (|{_zz_TrapPlugin_logic_harts_0_trap_pending_arbiter_ports_1_valid_1,_zz_TrapPlugin_logic_harts_0_trap_pending_arbiter_ports_1_valid});
  assign _zz_TrapPlugin_logic_harts_0_trap_pending_arbiter_ports_1_payload_exception_1 = ((_zz_TrapPlugin_logic_harts_0_trap_pending_arbiter_ports_1_payload_exception[0] ? {early0_EnvPlugin_logic_trapPort_payload_arg,{early0_EnvPlugin_logic_trapPort_payload_code,{early0_EnvPlugin_logic_trapPort_payload_tval,early0_EnvPlugin_logic_trapPort_payload_exception}}} : 40'h0) | (_zz_TrapPlugin_logic_harts_0_trap_pending_arbiter_ports_1_payload_exception[1] ? {CsrAccessPlugin_logic_trapPort_payload_arg,{CsrAccessPlugin_logic_trapPort_payload_code,{CsrAccessPlugin_logic_trapPort_payload_tval,CsrAccessPlugin_logic_trapPort_payload_exception}}} : 40'h0));
  assign TrapPlugin_logic_harts_0_trap_pending_arbiter_ports_1_payload_exception = _zz_TrapPlugin_logic_harts_0_trap_pending_arbiter_ports_1_payload_exception_1[0];
  assign TrapPlugin_logic_harts_0_trap_pending_arbiter_ports_1_payload_tval = _zz_TrapPlugin_logic_harts_0_trap_pending_arbiter_ports_1_payload_exception_1[32 : 1];
  assign TrapPlugin_logic_harts_0_trap_pending_arbiter_ports_1_payload_code = _zz_TrapPlugin_logic_harts_0_trap_pending_arbiter_ports_1_payload_exception_1[36 : 33];
  assign TrapPlugin_logic_harts_0_trap_pending_arbiter_ports_1_payload_arg = _zz_TrapPlugin_logic_harts_0_trap_pending_arbiter_ports_1_payload_exception_1[39 : 37];
  assign _zz_TrapPlugin_logic_harts_0_trap_pending_arbiter_ports_2_payload_exception = {(_zz_TrapPlugin_logic_harts_0_trap_pending_arbiter_ports_2_valid_1 && (&(! (_zz_TrapPlugin_logic_harts_0_trap_pending_arbiter_ports_2_valid && (DecoderPlugin_logic_laneLogic_0_trapPort_payload_laneAge < DecoderPlugin_logic_laneLogic_1_trapPort_payload_laneAge))))),(_zz_TrapPlugin_logic_harts_0_trap_pending_arbiter_ports_2_valid && (&(! (_zz_TrapPlugin_logic_harts_0_trap_pending_arbiter_ports_2_valid_1 && (DecoderPlugin_logic_laneLogic_1_trapPort_payload_laneAge < DecoderPlugin_logic_laneLogic_0_trapPort_payload_laneAge)))))};
  assign TrapPlugin_logic_harts_0_trap_pending_arbiter_ports_2_valid = (|{_zz_TrapPlugin_logic_harts_0_trap_pending_arbiter_ports_2_valid_1,_zz_TrapPlugin_logic_harts_0_trap_pending_arbiter_ports_2_valid});
  assign _zz_TrapPlugin_logic_harts_0_trap_pending_arbiter_ports_2_payload_exception_1 = ((_zz_TrapPlugin_logic_harts_0_trap_pending_arbiter_ports_2_payload_exception[0] ? {DecoderPlugin_logic_laneLogic_0_trapPort_payload_arg,{DecoderPlugin_logic_laneLogic_0_trapPort_payload_code,{DecoderPlugin_logic_laneLogic_0_trapPort_payload_tval,DecoderPlugin_logic_laneLogic_0_trapPort_payload_exception}}} : 40'h0) | (_zz_TrapPlugin_logic_harts_0_trap_pending_arbiter_ports_2_payload_exception[1] ? {DecoderPlugin_logic_laneLogic_1_trapPort_payload_arg,{DecoderPlugin_logic_laneLogic_1_trapPort_payload_code,{DecoderPlugin_logic_laneLogic_1_trapPort_payload_tval,DecoderPlugin_logic_laneLogic_1_trapPort_payload_exception}}} : 40'h0));
  assign TrapPlugin_logic_harts_0_trap_pending_arbiter_ports_2_payload_exception = _zz_TrapPlugin_logic_harts_0_trap_pending_arbiter_ports_2_payload_exception_1[0];
  assign TrapPlugin_logic_harts_0_trap_pending_arbiter_ports_2_payload_tval = _zz_TrapPlugin_logic_harts_0_trap_pending_arbiter_ports_2_payload_exception_1[32 : 1];
  assign TrapPlugin_logic_harts_0_trap_pending_arbiter_ports_2_payload_code = _zz_TrapPlugin_logic_harts_0_trap_pending_arbiter_ports_2_payload_exception_1[36 : 33];
  assign TrapPlugin_logic_harts_0_trap_pending_arbiter_ports_2_payload_arg = _zz_TrapPlugin_logic_harts_0_trap_pending_arbiter_ports_2_payload_exception_1[39 : 37];
  assign TrapPlugin_logic_harts_0_trap_pending_arbiter_ports_3_valid = (|_zz_TrapPlugin_logic_harts_0_trap_pending_arbiter_ports_3_valid);
  assign TrapPlugin_logic_harts_0_trap_pending_arbiter_ports_3_payload_exception = FetchL1Plugin_logic_trapPort_payload_exception;
  assign TrapPlugin_logic_harts_0_trap_pending_arbiter_ports_3_payload_tval = FetchL1Plugin_logic_trapPort_payload_tval;
  assign TrapPlugin_logic_harts_0_trap_pending_arbiter_ports_3_payload_code = FetchL1Plugin_logic_trapPort_payload_code;
  assign TrapPlugin_logic_harts_0_trap_pending_arbiter_ports_3_payload_arg = FetchL1Plugin_logic_trapPort_payload_arg;
  assign _zz_TrapPlugin_logic_harts_0_trap_pending_arbiter_oh = {TrapPlugin_logic_harts_0_trap_pending_arbiter_ports_3_valid,{TrapPlugin_logic_harts_0_trap_pending_arbiter_ports_2_valid,{TrapPlugin_logic_harts_0_trap_pending_arbiter_ports_1_valid,TrapPlugin_logic_harts_0_trap_pending_arbiter_ports_0_valid}}};
  assign _zz_TrapPlugin_logic_harts_0_trap_pending_arbiter_oh_1 = _zz_TrapPlugin_logic_harts_0_trap_pending_arbiter_oh[0];
  assign _zz_TrapPlugin_logic_harts_0_trap_pending_arbiter_oh_2 = _zz_TrapPlugin_logic_harts_0_trap_pending_arbiter_oh[1];
  assign _zz_TrapPlugin_logic_harts_0_trap_pending_arbiter_oh_3 = _zz_TrapPlugin_logic_harts_0_trap_pending_arbiter_oh[2];
  always @(*) begin
    _zz_TrapPlugin_logic_harts_0_trap_pending_arbiter_oh_4[0] = (_zz_TrapPlugin_logic_harts_0_trap_pending_arbiter_oh_1 && (! 1'b0));
    _zz_TrapPlugin_logic_harts_0_trap_pending_arbiter_oh_4[1] = (_zz_TrapPlugin_logic_harts_0_trap_pending_arbiter_oh_2 && (! _zz_TrapPlugin_logic_harts_0_trap_pending_arbiter_oh_1));
    _zz_TrapPlugin_logic_harts_0_trap_pending_arbiter_oh_4[2] = (_zz_TrapPlugin_logic_harts_0_trap_pending_arbiter_oh_3 && (! (|{_zz_TrapPlugin_logic_harts_0_trap_pending_arbiter_oh_2,_zz_TrapPlugin_logic_harts_0_trap_pending_arbiter_oh_1})));
    _zz_TrapPlugin_logic_harts_0_trap_pending_arbiter_oh_4[3] = (_zz_TrapPlugin_logic_harts_0_trap_pending_arbiter_oh[3] && (! (|{_zz_TrapPlugin_logic_harts_0_trap_pending_arbiter_oh_3,{_zz_TrapPlugin_logic_harts_0_trap_pending_arbiter_oh_2,_zz_TrapPlugin_logic_harts_0_trap_pending_arbiter_oh_1}})));
  end

  assign TrapPlugin_logic_harts_0_trap_pending_arbiter_oh = _zz_TrapPlugin_logic_harts_0_trap_pending_arbiter_oh_4;
  assign TrapPlugin_logic_harts_0_trap_pending_arbiter_down_valid = (|{_zz_TrapPlugin_logic_harts_0_trap_pending_arbiter_ports_2_valid_1,{_zz_TrapPlugin_logic_harts_0_trap_pending_arbiter_ports_2_valid,{_zz_TrapPlugin_logic_harts_0_trap_pending_arbiter_ports_1_valid_1,{_zz_TrapPlugin_logic_harts_0_trap_pending_arbiter_ports_0_valid,{_zz_TrapPlugin_logic_harts_0_trap_pending_arbiter_ports_3_valid,_zz_TrapPlugin_logic_harts_0_trap_pending_arbiter_ports_1_valid}}}}});
  assign _zz_TrapPlugin_logic_harts_0_trap_pending_arbiter_down_payload_exception = (((TrapPlugin_logic_harts_0_trap_pending_arbiter_oh[0] ? {TrapPlugin_logic_harts_0_trap_pending_arbiter_ports_0_payload_arg,{TrapPlugin_logic_harts_0_trap_pending_arbiter_ports_0_payload_code,_zz__zz_TrapPlugin_logic_harts_0_trap_pending_arbiter_down_payload_exception}} : 40'h0) | (TrapPlugin_logic_harts_0_trap_pending_arbiter_oh[1] ? {TrapPlugin_logic_harts_0_trap_pending_arbiter_ports_1_payload_arg,{TrapPlugin_logic_harts_0_trap_pending_arbiter_ports_1_payload_code,_zz__zz_TrapPlugin_logic_harts_0_trap_pending_arbiter_down_payload_exception_1}} : 40'h0)) | ((TrapPlugin_logic_harts_0_trap_pending_arbiter_oh[2] ? {TrapPlugin_logic_harts_0_trap_pending_arbiter_ports_2_payload_arg,{TrapPlugin_logic_harts_0_trap_pending_arbiter_ports_2_payload_code,_zz__zz_TrapPlugin_logic_harts_0_trap_pending_arbiter_down_payload_exception_2}} : 40'h0) | (TrapPlugin_logic_harts_0_trap_pending_arbiter_oh[3] ? {TrapPlugin_logic_harts_0_trap_pending_arbiter_ports_3_payload_arg,{TrapPlugin_logic_harts_0_trap_pending_arbiter_ports_3_payload_code,_zz__zz_TrapPlugin_logic_harts_0_trap_pending_arbiter_down_payload_exception_3}} : 40'h0)));
  assign TrapPlugin_logic_harts_0_trap_pending_arbiter_down_payload_exception = _zz_TrapPlugin_logic_harts_0_trap_pending_arbiter_down_payload_exception[0];
  assign TrapPlugin_logic_harts_0_trap_pending_arbiter_down_payload_tval = _zz_TrapPlugin_logic_harts_0_trap_pending_arbiter_down_payload_exception[32 : 1];
  assign TrapPlugin_logic_harts_0_trap_pending_arbiter_down_payload_code = _zz_TrapPlugin_logic_harts_0_trap_pending_arbiter_down_payload_exception[36 : 33];
  assign TrapPlugin_logic_harts_0_trap_pending_arbiter_down_payload_arg = _zz_TrapPlugin_logic_harts_0_trap_pending_arbiter_down_payload_exception[39 : 37];
  assign TrapPlugin_logic_harts_0_trap_pending_xret_sourcePrivilege = TrapPlugin_logic_harts_0_trap_pending_state_arg[1 : 0];
  always @(*) begin
    TrapPlugin_logic_harts_0_trap_pending_xret_targetPrivilege = PrivilegedPlugin_logic_harts_0_m_status_mpp;
    case(TrapPlugin_logic_harts_0_trap_pending_xret_sourcePrivilege)
      2'b01 : begin
        TrapPlugin_logic_harts_0_trap_pending_xret_targetPrivilege = {1'b0,PrivilegedPlugin_logic_harts_0_s_status_spp};
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    TrapPlugin_logic_harts_0_trap_exception_exceptionTargetPrivilegeUncapped = 2'b11;
    case(TrapPlugin_logic_harts_0_trap_exception_code)
      4'b0000 : begin
        if(when_TrapPlugin_l251) begin
          TrapPlugin_logic_harts_0_trap_exception_exceptionTargetPrivilegeUncapped = 2'b01;
        end
      end
      4'b0011 : begin
        if(when_TrapPlugin_l251_1) begin
          TrapPlugin_logic_harts_0_trap_exception_exceptionTargetPrivilegeUncapped = 2'b01;
        end
      end
      4'b1000 : begin
        if(when_TrapPlugin_l251_2) begin
          TrapPlugin_logic_harts_0_trap_exception_exceptionTargetPrivilegeUncapped = 2'b01;
        end
      end
      4'b1001 : begin
        if(when_TrapPlugin_l251_3) begin
          TrapPlugin_logic_harts_0_trap_exception_exceptionTargetPrivilegeUncapped = 2'b01;
        end
      end
      4'b1100 : begin
        if(when_TrapPlugin_l251_4) begin
          TrapPlugin_logic_harts_0_trap_exception_exceptionTargetPrivilegeUncapped = 2'b01;
        end
      end
      4'b1101 : begin
        if(when_TrapPlugin_l251_5) begin
          TrapPlugin_logic_harts_0_trap_exception_exceptionTargetPrivilegeUncapped = 2'b01;
        end
      end
      4'b1111 : begin
        if(when_TrapPlugin_l251_6) begin
          TrapPlugin_logic_harts_0_trap_exception_exceptionTargetPrivilegeUncapped = 2'b01;
        end
      end
      default : begin
      end
    endcase
  end

  assign TrapPlugin_logic_harts_0_trap_exception_code = TrapPlugin_logic_harts_0_trap_pending_state_code;
  assign when_TrapPlugin_l251 = ((1'b1 && PrivilegedPlugin_logic_harts_0_m_edeleg_iam) && (! 1'b0));
  assign when_TrapPlugin_l251_1 = ((1'b1 && PrivilegedPlugin_logic_harts_0_m_edeleg_bp) && (! 1'b0));
  assign when_TrapPlugin_l251_2 = ((1'b1 && PrivilegedPlugin_logic_harts_0_m_edeleg_eu) && (! 1'b0));
  assign when_TrapPlugin_l251_3 = ((1'b1 && PrivilegedPlugin_logic_harts_0_m_edeleg_es) && (! 1'b0));
  assign when_TrapPlugin_l251_4 = ((1'b1 && PrivilegedPlugin_logic_harts_0_m_edeleg_ipf) && (! 1'b0));
  assign when_TrapPlugin_l251_5 = ((1'b1 && PrivilegedPlugin_logic_harts_0_m_edeleg_lpf) && (! 1'b0));
  assign when_TrapPlugin_l251_6 = ((1'b1 && PrivilegedPlugin_logic_harts_0_m_edeleg_spf) && (! 1'b0));
  assign TrapPlugin_logic_harts_0_trap_exception_targetPrivilege = ((PrivilegedPlugin_logic_harts_0_privilege < TrapPlugin_logic_harts_0_trap_exception_exceptionTargetPrivilegeUncapped) ? TrapPlugin_logic_harts_0_trap_exception_exceptionTargetPrivilegeUncapped : PrivilegedPlugin_logic_harts_0_privilege);
  assign PrivilegedPlugin_logic_harts_0_commitMask = {(((toplevel_execute_ctrl5_down_LANE_SEL_lane1 && toplevel_execute_ctrl5_down_isReady) && (! toplevel_execute_lane1_ctrls_5_downIsCancel)) && toplevel_execute_ctrl5_down_COMMIT_lane1),(((toplevel_execute_ctrl5_down_LANE_SEL_lane0 && toplevel_execute_ctrl5_down_isReady) && (! toplevel_execute_lane0_ctrls_5_downIsCancel)) && toplevel_execute_ctrl5_down_COMMIT_lane0)};
  assign TrapPlugin_logic_harts_0_trap_trigger_oh = {(((toplevel_execute_ctrl4_down_LANE_SEL_lane1 && toplevel_execute_ctrl4_down_isReady) && (! toplevel_execute_lane1_ctrls_4_downIsCancel)) && toplevel_execute_ctrl4_down_TRAP_lane1),(((toplevel_execute_ctrl4_down_LANE_SEL_lane0 && toplevel_execute_ctrl4_down_isReady) && (! toplevel_execute_lane0_ctrls_4_downIsCancel)) && toplevel_execute_ctrl4_down_TRAP_lane0)};
  assign TrapPlugin_logic_harts_0_trap_trigger_valid = (|TrapPlugin_logic_harts_0_trap_trigger_oh);
  assign _zz_TrapPlugin_logic_harts_0_trap_pending_pc = TrapPlugin_logic_harts_0_trap_trigger_oh[0];
  assign _zz_TrapPlugin_logic_harts_0_trap_pending_pc_1 = TrapPlugin_logic_harts_0_trap_trigger_oh[1];
  always @(*) begin
    TrapPlugin_logic_harts_0_trap_whitebox_trap = 1'b0;
    case(TrapPlugin_logic_harts_0_trap_fsm_stateReg)
      TrapPlugin_logic_harts_0_trap_fsm_enumDef_RUNNING : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_enumDef_PROCESS_1 : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_enumDef_TRAP_EPC : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_enumDef_TRAP_TVAL : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_enumDef_TRAP_TVEC : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_enumDef_TRAP_APPLY : begin
        TrapPlugin_logic_harts_0_trap_whitebox_trap = 1'b1;
      end
      TrapPlugin_logic_harts_0_trap_fsm_enumDef_XRET_EPC : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_enumDef_XRET_APPLY : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_enumDef_ATS_RSP : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_enumDef_JUMP : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_enumDef_LSU_FLUSH : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_enumDef_FETCH_FLUSH : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    TrapPlugin_logic_harts_0_trap_whitebox_interrupt = 1'bx;
    case(TrapPlugin_logic_harts_0_trap_fsm_stateReg)
      TrapPlugin_logic_harts_0_trap_fsm_enumDef_RUNNING : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_enumDef_PROCESS_1 : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_enumDef_TRAP_EPC : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_enumDef_TRAP_TVAL : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_enumDef_TRAP_TVEC : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_enumDef_TRAP_APPLY : begin
        TrapPlugin_logic_harts_0_trap_whitebox_interrupt = TrapPlugin_logic_harts_0_trap_fsm_buffer_trap_interrupt;
      end
      TrapPlugin_logic_harts_0_trap_fsm_enumDef_XRET_EPC : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_enumDef_XRET_APPLY : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_enumDef_ATS_RSP : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_enumDef_JUMP : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_enumDef_LSU_FLUSH : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_enumDef_FETCH_FLUSH : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    TrapPlugin_logic_harts_0_trap_whitebox_code = 4'bxxxx;
    case(TrapPlugin_logic_harts_0_trap_fsm_stateReg)
      TrapPlugin_logic_harts_0_trap_fsm_enumDef_RUNNING : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_enumDef_PROCESS_1 : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_enumDef_TRAP_EPC : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_enumDef_TRAP_TVAL : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_enumDef_TRAP_TVEC : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_enumDef_TRAP_APPLY : begin
        TrapPlugin_logic_harts_0_trap_whitebox_code = TrapPlugin_logic_harts_0_trap_fsm_buffer_trap_code;
      end
      TrapPlugin_logic_harts_0_trap_fsm_enumDef_XRET_EPC : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_enumDef_XRET_APPLY : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_enumDef_ATS_RSP : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_enumDef_JUMP : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_enumDef_LSU_FLUSH : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_enumDef_FETCH_FLUSH : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    TrapPlugin_logic_harts_0_trap_historyPort_valid = 1'b0;
    case(TrapPlugin_logic_harts_0_trap_fsm_stateReg)
      TrapPlugin_logic_harts_0_trap_fsm_enumDef_RUNNING : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_enumDef_PROCESS_1 : begin
        TrapPlugin_logic_harts_0_trap_historyPort_valid = 1'b1;
      end
      TrapPlugin_logic_harts_0_trap_fsm_enumDef_TRAP_EPC : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_enumDef_TRAP_TVAL : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_enumDef_TRAP_TVEC : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_enumDef_TRAP_APPLY : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_enumDef_XRET_EPC : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_enumDef_XRET_APPLY : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_enumDef_ATS_RSP : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_enumDef_JUMP : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_enumDef_LSU_FLUSH : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_enumDef_FETCH_FLUSH : begin
      end
      default : begin
      end
    endcase
  end

  assign TrapPlugin_logic_harts_0_trap_historyPort_payload_history = TrapPlugin_logic_harts_0_trap_pending_history;
  always @(*) begin
    TrapPlugin_logic_harts_0_trap_pcPort_valid = 1'b0;
    case(TrapPlugin_logic_harts_0_trap_fsm_stateReg)
      TrapPlugin_logic_harts_0_trap_fsm_enumDef_RUNNING : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_enumDef_PROCESS_1 : begin
        if(!when_TrapPlugin_l393) begin
          case(TrapPlugin_logic_harts_0_trap_pending_state_code)
            4'b0000 : begin
              TrapPlugin_logic_harts_0_trap_pcPort_valid = 1'b1;
            end
            4'b0001 : begin
            end
            4'b0010 : begin
            end
            4'b0100 : begin
            end
            4'b0101 : begin
            end
            4'b1000 : begin
            end
            4'b0110 : begin
            end
            4'b0111 : begin
            end
            default : begin
            end
          endcase
        end
      end
      TrapPlugin_logic_harts_0_trap_fsm_enumDef_TRAP_EPC : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_enumDef_TRAP_TVAL : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_enumDef_TRAP_TVEC : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_enumDef_TRAP_APPLY : begin
        TrapPlugin_logic_harts_0_trap_pcPort_valid = 1'b1;
      end
      TrapPlugin_logic_harts_0_trap_fsm_enumDef_XRET_EPC : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_enumDef_XRET_APPLY : begin
        TrapPlugin_logic_harts_0_trap_pcPort_valid = 1'b1;
      end
      TrapPlugin_logic_harts_0_trap_fsm_enumDef_ATS_RSP : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_enumDef_JUMP : begin
        TrapPlugin_logic_harts_0_trap_pcPort_valid = 1'b1;
      end
      TrapPlugin_logic_harts_0_trap_fsm_enumDef_LSU_FLUSH : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_enumDef_FETCH_FLUSH : begin
      end
      default : begin
      end
    endcase
  end

  assign TrapPlugin_logic_harts_0_trap_pcPort_payload_fault = 1'b0;
  always @(*) begin
    TrapPlugin_logic_harts_0_trap_pcPort_payload_pc = 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
    case(TrapPlugin_logic_harts_0_trap_fsm_stateReg)
      TrapPlugin_logic_harts_0_trap_fsm_enumDef_RUNNING : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_enumDef_PROCESS_1 : begin
        if(!when_TrapPlugin_l393) begin
          case(TrapPlugin_logic_harts_0_trap_pending_state_code)
            4'b0000 : begin
              TrapPlugin_logic_harts_0_trap_pcPort_payload_pc = TrapPlugin_logic_harts_0_trap_pending_pc;
            end
            4'b0001 : begin
            end
            4'b0010 : begin
            end
            4'b0100 : begin
            end
            4'b0101 : begin
            end
            4'b1000 : begin
            end
            4'b0110 : begin
            end
            4'b0111 : begin
            end
            default : begin
            end
          endcase
        end
      end
      TrapPlugin_logic_harts_0_trap_fsm_enumDef_TRAP_EPC : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_enumDef_TRAP_TVAL : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_enumDef_TRAP_TVEC : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_enumDef_TRAP_APPLY : begin
        TrapPlugin_logic_harts_0_trap_pcPort_payload_pc = TrapPlugin_logic_harts_0_trap_fsm_readed;
      end
      TrapPlugin_logic_harts_0_trap_fsm_enumDef_XRET_EPC : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_enumDef_XRET_APPLY : begin
        TrapPlugin_logic_harts_0_trap_pcPort_payload_pc = TrapPlugin_logic_harts_0_trap_fsm_readed;
      end
      TrapPlugin_logic_harts_0_trap_fsm_enumDef_ATS_RSP : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_enumDef_JUMP : begin
        TrapPlugin_logic_harts_0_trap_pcPort_payload_pc = TrapPlugin_logic_harts_0_trap_fsm_jumpTarget;
      end
      TrapPlugin_logic_harts_0_trap_fsm_enumDef_LSU_FLUSH : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_enumDef_FETCH_FLUSH : begin
      end
      default : begin
      end
    endcase
  end

  assign TrapPlugin_logic_harts_0_trap_fsm_wantExit = 1'b0;
  always @(*) begin
    TrapPlugin_logic_harts_0_trap_fsm_wantStart = 1'b0;
    case(TrapPlugin_logic_harts_0_trap_fsm_stateReg)
      TrapPlugin_logic_harts_0_trap_fsm_enumDef_RUNNING : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_enumDef_PROCESS_1 : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_enumDef_TRAP_EPC : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_enumDef_TRAP_TVAL : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_enumDef_TRAP_TVEC : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_enumDef_TRAP_APPLY : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_enumDef_XRET_EPC : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_enumDef_XRET_APPLY : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_enumDef_ATS_RSP : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_enumDef_JUMP : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_enumDef_LSU_FLUSH : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_enumDef_FETCH_FLUSH : begin
      end
      default : begin
        TrapPlugin_logic_harts_0_trap_fsm_wantStart = 1'b1;
      end
    endcase
  end

  assign TrapPlugin_logic_harts_0_trap_fsm_wantKill = 1'b0;
  assign TrapPlugin_logic_harts_0_trap_fsm_inflightTrap = (|{execute_lane1_logic_trapPending[0],{execute_lane0_logic_trapPending[0],{DispatchPlugin_logic_trapPendings[0],decode_logic_trapPending[0]}}});
  assign TrapPlugin_logic_harts_0_trap_fsm_holdPort = (TrapPlugin_logic_harts_0_trap_fsm_inflightTrap || (! (TrapPlugin_logic_harts_0_trap_fsm_stateReg == TrapPlugin_logic_harts_0_trap_fsm_enumDef_RUNNING)));
  assign TrapPlugin_api_harts_0_fsmBusy = (! (TrapPlugin_logic_harts_0_trap_fsm_stateReg == TrapPlugin_logic_harts_0_trap_fsm_enumDef_RUNNING));
  always @(*) begin
    TrapPlugin_logic_harts_0_trap_fsm_wfi = 1'b0;
    case(TrapPlugin_logic_harts_0_trap_fsm_stateReg)
      TrapPlugin_logic_harts_0_trap_fsm_enumDef_RUNNING : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_enumDef_PROCESS_1 : begin
        if(!when_TrapPlugin_l393) begin
          case(TrapPlugin_logic_harts_0_trap_pending_state_code)
            4'b0000 : begin
            end
            4'b0001 : begin
            end
            4'b0010 : begin
            end
            4'b0100 : begin
            end
            4'b0101 : begin
            end
            4'b1000 : begin
              TrapPlugin_logic_harts_0_trap_fsm_wfi = 1'b1;
            end
            4'b0110 : begin
            end
            4'b0111 : begin
            end
            default : begin
            end
          endcase
        end
      end
      TrapPlugin_logic_harts_0_trap_fsm_enumDef_TRAP_EPC : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_enumDef_TRAP_TVAL : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_enumDef_TRAP_TVEC : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_enumDef_TRAP_APPLY : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_enumDef_XRET_EPC : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_enumDef_XRET_APPLY : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_enumDef_ATS_RSP : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_enumDef_JUMP : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_enumDef_LSU_FLUSH : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_enumDef_FETCH_FLUSH : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    TrapPlugin_logic_harts_0_trap_fsm_buffer_sampleIt = 1'b0;
    case(TrapPlugin_logic_harts_0_trap_fsm_stateReg)
      TrapPlugin_logic_harts_0_trap_fsm_enumDef_RUNNING : begin
        if(TrapPlugin_logic_harts_0_trap_trigger_valid) begin
          TrapPlugin_logic_harts_0_trap_fsm_buffer_sampleIt = 1'b1;
        end
      end
      TrapPlugin_logic_harts_0_trap_fsm_enumDef_PROCESS_1 : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_enumDef_TRAP_EPC : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_enumDef_TRAP_TVAL : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_enumDef_TRAP_TVEC : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_enumDef_TRAP_APPLY : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_enumDef_XRET_EPC : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_enumDef_XRET_APPLY : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_enumDef_ATS_RSP : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_enumDef_JUMP : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_enumDef_LSU_FLUSH : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_enumDef_FETCH_FLUSH : begin
      end
      default : begin
      end
    endcase
  end

  assign TrapPlugin_logic_harts_0_trap_fsm_buffer_trap_interrupt = ((TrapPlugin_logic_harts_0_trap_pending_state_code == 4'b0000) && TrapPlugin_logic_harts_0_trap_fsm_buffer_i_valid);
  assign TrapPlugin_logic_harts_0_trap_fsm_buffer_trap_targetPrivilege = (TrapPlugin_logic_harts_0_trap_fsm_buffer_trap_interrupt ? TrapPlugin_logic_harts_0_trap_fsm_buffer_i_targetPrivilege : TrapPlugin_logic_harts_0_trap_exception_targetPrivilege);
  assign TrapPlugin_logic_harts_0_trap_fsm_buffer_trap_tval = ((! TrapPlugin_logic_harts_0_trap_fsm_buffer_trap_interrupt) ? TrapPlugin_logic_harts_0_trap_pending_state_tval : 32'h0);
  assign TrapPlugin_logic_harts_0_trap_fsm_buffer_trap_code = (TrapPlugin_logic_harts_0_trap_fsm_buffer_trap_interrupt ? TrapPlugin_logic_harts_0_trap_fsm_buffer_i_code : TrapPlugin_logic_harts_0_trap_pending_state_code);
  assign TrapPlugin_logic_harts_0_trap_fsm_resetToRunConditions_0 = (! TrapPlugin_logic_initHold);
  always @(*) begin
    TrapPlugin_logic_harts_0_trap_fsm_atsPorts_refill_cmd_valid = 1'b0;
    case(TrapPlugin_logic_harts_0_trap_fsm_stateReg)
      TrapPlugin_logic_harts_0_trap_fsm_enumDef_RUNNING : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_enumDef_PROCESS_1 : begin
        if(!when_TrapPlugin_l393) begin
          case(TrapPlugin_logic_harts_0_trap_pending_state_code)
            4'b0000 : begin
            end
            4'b0001 : begin
            end
            4'b0010 : begin
            end
            4'b0100 : begin
            end
            4'b0101 : begin
            end
            4'b1000 : begin
            end
            4'b0110 : begin
            end
            4'b0111 : begin
              TrapPlugin_logic_harts_0_trap_fsm_atsPorts_refill_cmd_valid = 1'b1;
            end
            default : begin
            end
          endcase
        end
      end
      TrapPlugin_logic_harts_0_trap_fsm_enumDef_TRAP_EPC : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_enumDef_TRAP_TVAL : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_enumDef_TRAP_TVEC : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_enumDef_TRAP_APPLY : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_enumDef_XRET_EPC : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_enumDef_XRET_APPLY : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_enumDef_ATS_RSP : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_enumDef_JUMP : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_enumDef_LSU_FLUSH : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_enumDef_FETCH_FLUSH : begin
      end
      default : begin
      end
    endcase
  end

  assign TrapPlugin_logic_harts_0_trap_fsm_atsPorts_refill_cmd_payload_address = TrapPlugin_logic_harts_0_trap_pending_state_tval;
  assign TrapPlugin_logic_harts_0_trap_fsm_atsPorts_refill_cmd_payload_storageId = TrapPlugin_logic_harts_0_trap_pending_state_arg[2 : 2];
  always @(*) begin
    TrapPlugin_logic_harts_0_trap_fsm_atsPorts_invalidate_cmd_valid = 1'b0;
    if(when_TrapPlugin_l340) begin
      TrapPlugin_logic_harts_0_trap_fsm_atsPorts_invalidate_cmd_valid = 1'b1;
    end
    case(TrapPlugin_logic_harts_0_trap_fsm_stateReg)
      TrapPlugin_logic_harts_0_trap_fsm_enumDef_RUNNING : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_enumDef_PROCESS_1 : begin
        if(!when_TrapPlugin_l393) begin
          case(TrapPlugin_logic_harts_0_trap_pending_state_code)
            4'b0000 : begin
            end
            4'b0001 : begin
            end
            4'b0010 : begin
            end
            4'b0100 : begin
            end
            4'b0101 : begin
            end
            4'b1000 : begin
            end
            4'b0110 : begin
              TrapPlugin_logic_harts_0_trap_fsm_atsPorts_invalidate_cmd_valid = 1'b1;
            end
            4'b0111 : begin
            end
            default : begin
            end
          endcase
        end
      end
      TrapPlugin_logic_harts_0_trap_fsm_enumDef_TRAP_EPC : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_enumDef_TRAP_TVAL : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_enumDef_TRAP_TVEC : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_enumDef_TRAP_APPLY : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_enumDef_XRET_EPC : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_enumDef_XRET_APPLY : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_enumDef_ATS_RSP : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_enumDef_JUMP : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_enumDef_LSU_FLUSH : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_enumDef_FETCH_FLUSH : begin
      end
      default : begin
      end
    endcase
  end

  assign TrapPlugin_logic_harts_0_trap_fsm_atsPorts_invalidate_cmd_fire = (TrapPlugin_logic_harts_0_trap_fsm_atsPorts_invalidate_cmd_valid && TrapPlugin_logic_harts_0_trap_fsm_atsPorts_invalidate_cmd_ready);
  assign when_TrapPlugin_l340 = (! TrapPlugin_logic_harts_0_trap_fsm_atsPorts_invalidated);
  assign TrapPlugin_logic_harts_0_trap_fsm_jumpOffset = ((|{(TrapPlugin_logic_harts_0_trap_pending_state_code == 4'b1000),{(TrapPlugin_logic_harts_0_trap_pending_state_code == 4'b0110),{(TrapPlugin_logic_harts_0_trap_pending_state_code == 4'b0010),(TrapPlugin_logic_harts_0_trap_pending_state_code == 4'b0101)}}}) ? TrapPlugin_logic_harts_0_trap_pending_slices : 2'b00);
  always @(*) begin
    TrapPlugin_logic_fetchL1Invalidate_0_cmd_valid = 1'b0;
    case(TrapPlugin_logic_harts_0_trap_fsm_stateReg)
      TrapPlugin_logic_harts_0_trap_fsm_enumDef_RUNNING : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_enumDef_PROCESS_1 : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_enumDef_TRAP_EPC : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_enumDef_TRAP_TVAL : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_enumDef_TRAP_TVEC : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_enumDef_TRAP_APPLY : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_enumDef_XRET_EPC : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_enumDef_XRET_APPLY : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_enumDef_ATS_RSP : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_enumDef_JUMP : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_enumDef_LSU_FLUSH : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_enumDef_FETCH_FLUSH : begin
        TrapPlugin_logic_fetchL1Invalidate_0_cmd_valid = 1'b1;
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    TrapPlugin_logic_lsuL1Invalidate_0_cmd_valid = 1'b0;
    case(TrapPlugin_logic_harts_0_trap_fsm_stateReg)
      TrapPlugin_logic_harts_0_trap_fsm_enumDef_RUNNING : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_enumDef_PROCESS_1 : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_enumDef_TRAP_EPC : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_enumDef_TRAP_TVAL : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_enumDef_TRAP_TVEC : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_enumDef_TRAP_APPLY : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_enumDef_XRET_EPC : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_enumDef_XRET_APPLY : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_enumDef_ATS_RSP : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_enumDef_JUMP : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_enumDef_LSU_FLUSH : begin
        TrapPlugin_logic_lsuL1Invalidate_0_cmd_valid = 1'b1;
      end
      TrapPlugin_logic_harts_0_trap_fsm_enumDef_FETCH_FLUSH : begin
      end
      default : begin
      end
    endcase
  end

  assign TrapPlugin_logic_harts_0_trap_fsm_triggerEbreak = 1'b0;
  assign when_TrapPlugin_l539 = (TrapPlugin_logic_harts_0_crsPorts_read_valid && TrapPlugin_logic_harts_0_crsPorts_read_ready);
  assign TrapPlugin_logic_harts_0_trap_fsm_xretPrivilege = TrapPlugin_logic_harts_0_trap_pending_state_arg[1 : 0];
  always @(*) begin
    FetchL1Plugin_logic_translationStorage_logic_sl_0_write_mask = 2'b00;
    if(!when_MmuPlugin_l496) begin
      FetchL1Plugin_logic_translationStorage_logic_sl_0_write_mask = 2'b11;
    end
    case(MmuPlugin_logic_refill_stateReg)
      MmuPlugin_logic_refill_enumDef_IDLE : begin
      end
      MmuPlugin_logic_refill_enumDef_CMD_0 : begin
      end
      MmuPlugin_logic_refill_enumDef_CMD_1 : begin
      end
      MmuPlugin_logic_refill_enumDef_RSP_0 : begin
        if(MmuPlugin_logic_refill_load_rsp_valid) begin
          if(!MmuPlugin_logic_refill_load_rsp_payload_redo) begin
            FetchL1Plugin_logic_translationStorage_logic_sl_0_write_mask = (MmuPlugin_logic_refill_storageOhReg[0] ? _zz_FetchL1Plugin_logic_translationStorage_logic_sl_0_write_mask : 2'b00);
            if(when_MmuPlugin_l439) begin
              FetchL1Plugin_logic_translationStorage_logic_sl_0_write_mask = 2'b00;
            end
          end
        end
      end
      MmuPlugin_logic_refill_enumDef_RSP_1 : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    FetchL1Plugin_logic_translationStorage_logic_sl_0_write_address = 6'bxxxxxx;
    if(!when_MmuPlugin_l496) begin
      FetchL1Plugin_logic_translationStorage_logic_sl_0_write_address = MmuPlugin_logic_invalidate_counter;
    end
    case(MmuPlugin_logic_refill_stateReg)
      MmuPlugin_logic_refill_enumDef_IDLE : begin
      end
      MmuPlugin_logic_refill_enumDef_CMD_0 : begin
      end
      MmuPlugin_logic_refill_enumDef_CMD_1 : begin
      end
      MmuPlugin_logic_refill_enumDef_RSP_0 : begin
        if(MmuPlugin_logic_refill_load_rsp_valid) begin
          if(!MmuPlugin_logic_refill_load_rsp_payload_redo) begin
            FetchL1Plugin_logic_translationStorage_logic_sl_0_write_address = MmuPlugin_logic_refill_virtual[17 : 12];
          end
        end
      end
      MmuPlugin_logic_refill_enumDef_RSP_1 : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    FetchL1Plugin_logic_translationStorage_logic_sl_0_write_data_valid = 1'bx;
    if(!when_MmuPlugin_l496) begin
      FetchL1Plugin_logic_translationStorage_logic_sl_0_write_data_valid = 1'b0;
    end
    case(MmuPlugin_logic_refill_stateReg)
      MmuPlugin_logic_refill_enumDef_IDLE : begin
      end
      MmuPlugin_logic_refill_enumDef_CMD_0 : begin
      end
      MmuPlugin_logic_refill_enumDef_CMD_1 : begin
      end
      MmuPlugin_logic_refill_enumDef_RSP_0 : begin
        if(MmuPlugin_logic_refill_load_rsp_valid) begin
          if(!MmuPlugin_logic_refill_load_rsp_payload_redo) begin
            FetchL1Plugin_logic_translationStorage_logic_sl_0_write_data_valid = 1'b1;
          end
        end
      end
      MmuPlugin_logic_refill_enumDef_RSP_1 : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    FetchL1Plugin_logic_translationStorage_logic_sl_0_write_data_virtualAddress = 14'bxxxxxxxxxxxxxx;
    case(MmuPlugin_logic_refill_stateReg)
      MmuPlugin_logic_refill_enumDef_IDLE : begin
      end
      MmuPlugin_logic_refill_enumDef_CMD_0 : begin
      end
      MmuPlugin_logic_refill_enumDef_CMD_1 : begin
      end
      MmuPlugin_logic_refill_enumDef_RSP_0 : begin
        if(MmuPlugin_logic_refill_load_rsp_valid) begin
          if(!MmuPlugin_logic_refill_load_rsp_payload_redo) begin
            FetchL1Plugin_logic_translationStorage_logic_sl_0_write_data_virtualAddress = MmuPlugin_logic_refill_virtual[31 : 18];
          end
        end
      end
      MmuPlugin_logic_refill_enumDef_RSP_1 : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    FetchL1Plugin_logic_translationStorage_logic_sl_0_write_data_physicalAddress = 20'bxxxxxxxxxxxxxxxxxxxx;
    case(MmuPlugin_logic_refill_stateReg)
      MmuPlugin_logic_refill_enumDef_IDLE : begin
      end
      MmuPlugin_logic_refill_enumDef_CMD_0 : begin
      end
      MmuPlugin_logic_refill_enumDef_CMD_1 : begin
      end
      MmuPlugin_logic_refill_enumDef_RSP_0 : begin
        if(MmuPlugin_logic_refill_load_rsp_valid) begin
          if(!MmuPlugin_logic_refill_load_rsp_payload_redo) begin
            FetchL1Plugin_logic_translationStorage_logic_sl_0_write_data_physicalAddress = (MmuPlugin_logic_refill_load_levelToPhysicalAddress_0 >>> 4'd12);
          end
        end
      end
      MmuPlugin_logic_refill_enumDef_RSP_1 : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    FetchL1Plugin_logic_translationStorage_logic_sl_0_write_data_allowRead = 1'bx;
    case(MmuPlugin_logic_refill_stateReg)
      MmuPlugin_logic_refill_enumDef_IDLE : begin
      end
      MmuPlugin_logic_refill_enumDef_CMD_0 : begin
      end
      MmuPlugin_logic_refill_enumDef_CMD_1 : begin
      end
      MmuPlugin_logic_refill_enumDef_RSP_0 : begin
        if(MmuPlugin_logic_refill_load_rsp_valid) begin
          if(!MmuPlugin_logic_refill_load_rsp_payload_redo) begin
            FetchL1Plugin_logic_translationStorage_logic_sl_0_write_data_allowRead = MmuPlugin_logic_refill_load_flags_R;
          end
        end
      end
      MmuPlugin_logic_refill_enumDef_RSP_1 : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    FetchL1Plugin_logic_translationStorage_logic_sl_0_write_data_allowWrite = 1'bx;
    case(MmuPlugin_logic_refill_stateReg)
      MmuPlugin_logic_refill_enumDef_IDLE : begin
      end
      MmuPlugin_logic_refill_enumDef_CMD_0 : begin
      end
      MmuPlugin_logic_refill_enumDef_CMD_1 : begin
      end
      MmuPlugin_logic_refill_enumDef_RSP_0 : begin
        if(MmuPlugin_logic_refill_load_rsp_valid) begin
          if(!MmuPlugin_logic_refill_load_rsp_payload_redo) begin
            FetchL1Plugin_logic_translationStorage_logic_sl_0_write_data_allowWrite = (MmuPlugin_logic_refill_load_flags_W && MmuPlugin_logic_refill_load_flags_D);
          end
        end
      end
      MmuPlugin_logic_refill_enumDef_RSP_1 : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    FetchL1Plugin_logic_translationStorage_logic_sl_0_write_data_allowExecute = 1'bx;
    case(MmuPlugin_logic_refill_stateReg)
      MmuPlugin_logic_refill_enumDef_IDLE : begin
      end
      MmuPlugin_logic_refill_enumDef_CMD_0 : begin
      end
      MmuPlugin_logic_refill_enumDef_CMD_1 : begin
      end
      MmuPlugin_logic_refill_enumDef_RSP_0 : begin
        if(MmuPlugin_logic_refill_load_rsp_valid) begin
          if(!MmuPlugin_logic_refill_load_rsp_payload_redo) begin
            FetchL1Plugin_logic_translationStorage_logic_sl_0_write_data_allowExecute = MmuPlugin_logic_refill_load_flags_X;
          end
        end
      end
      MmuPlugin_logic_refill_enumDef_RSP_1 : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    FetchL1Plugin_logic_translationStorage_logic_sl_0_write_data_allowUser = 1'bx;
    case(MmuPlugin_logic_refill_stateReg)
      MmuPlugin_logic_refill_enumDef_IDLE : begin
      end
      MmuPlugin_logic_refill_enumDef_CMD_0 : begin
      end
      MmuPlugin_logic_refill_enumDef_CMD_1 : begin
      end
      MmuPlugin_logic_refill_enumDef_RSP_0 : begin
        if(MmuPlugin_logic_refill_load_rsp_valid) begin
          if(!MmuPlugin_logic_refill_load_rsp_payload_redo) begin
            FetchL1Plugin_logic_translationStorage_logic_sl_0_write_data_allowUser = MmuPlugin_logic_refill_load_flags_U;
          end
        end
      end
      MmuPlugin_logic_refill_enumDef_RSP_1 : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    FetchL1Plugin_logic_translationStorage_logic_sl_0_allocId_willIncrement = 1'b0;
    case(MmuPlugin_logic_refill_stateReg)
      MmuPlugin_logic_refill_enumDef_IDLE : begin
      end
      MmuPlugin_logic_refill_enumDef_CMD_0 : begin
      end
      MmuPlugin_logic_refill_enumDef_CMD_1 : begin
      end
      MmuPlugin_logic_refill_enumDef_RSP_0 : begin
        if(MmuPlugin_logic_refill_load_rsp_valid) begin
          if(!MmuPlugin_logic_refill_load_rsp_payload_redo) begin
            FetchL1Plugin_logic_translationStorage_logic_sl_0_allocId_willIncrement = 1'b1;
          end
        end
      end
      MmuPlugin_logic_refill_enumDef_RSP_1 : begin
      end
      default : begin
      end
    endcase
  end

  assign FetchL1Plugin_logic_translationStorage_logic_sl_0_allocId_willClear = 1'b0;
  assign FetchL1Plugin_logic_translationStorage_logic_sl_0_allocId_willOverflowIfInc = (FetchL1Plugin_logic_translationStorage_logic_sl_0_allocId_value == 1'b1);
  assign FetchL1Plugin_logic_translationStorage_logic_sl_0_allocId_willOverflow = (FetchL1Plugin_logic_translationStorage_logic_sl_0_allocId_willOverflowIfInc && FetchL1Plugin_logic_translationStorage_logic_sl_0_allocId_willIncrement);
  always @(*) begin
    FetchL1Plugin_logic_translationStorage_logic_sl_0_allocId_valueNext = (FetchL1Plugin_logic_translationStorage_logic_sl_0_allocId_value + FetchL1Plugin_logic_translationStorage_logic_sl_0_allocId_willIncrement);
    if(FetchL1Plugin_logic_translationStorage_logic_sl_0_allocId_willClear) begin
      FetchL1Plugin_logic_translationStorage_logic_sl_0_allocId_valueNext = 1'b0;
    end
  end

  always @(*) begin
    FetchL1Plugin_logic_translationStorage_logic_sl_1_write_mask = 1'b0;
    if(!when_MmuPlugin_l496) begin
      FetchL1Plugin_logic_translationStorage_logic_sl_1_write_mask = 1'b1;
    end
    case(MmuPlugin_logic_refill_stateReg)
      MmuPlugin_logic_refill_enumDef_IDLE : begin
      end
      MmuPlugin_logic_refill_enumDef_CMD_0 : begin
      end
      MmuPlugin_logic_refill_enumDef_CMD_1 : begin
      end
      MmuPlugin_logic_refill_enumDef_RSP_0 : begin
      end
      MmuPlugin_logic_refill_enumDef_RSP_1 : begin
        if(MmuPlugin_logic_refill_load_rsp_valid) begin
          if(!MmuPlugin_logic_refill_load_rsp_payload_redo) begin
            if(when_MmuPlugin_l471) begin
              FetchL1Plugin_logic_translationStorage_logic_sl_1_write_mask = (MmuPlugin_logic_refill_storageOhReg[0] ? 1'b1 : 1'b0);
              if(when_MmuPlugin_l439_2) begin
                FetchL1Plugin_logic_translationStorage_logic_sl_1_write_mask = 1'b0;
              end
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    FetchL1Plugin_logic_translationStorage_logic_sl_1_write_address = 6'bxxxxxx;
    if(!when_MmuPlugin_l496) begin
      FetchL1Plugin_logic_translationStorage_logic_sl_1_write_address = MmuPlugin_logic_invalidate_counter;
    end
    case(MmuPlugin_logic_refill_stateReg)
      MmuPlugin_logic_refill_enumDef_IDLE : begin
      end
      MmuPlugin_logic_refill_enumDef_CMD_0 : begin
      end
      MmuPlugin_logic_refill_enumDef_CMD_1 : begin
      end
      MmuPlugin_logic_refill_enumDef_RSP_0 : begin
      end
      MmuPlugin_logic_refill_enumDef_RSP_1 : begin
        if(MmuPlugin_logic_refill_load_rsp_valid) begin
          if(!MmuPlugin_logic_refill_load_rsp_payload_redo) begin
            if(when_MmuPlugin_l471) begin
              FetchL1Plugin_logic_translationStorage_logic_sl_1_write_address = MmuPlugin_logic_refill_virtual[27 : 22];
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    FetchL1Plugin_logic_translationStorage_logic_sl_1_write_data_valid = 1'bx;
    if(!when_MmuPlugin_l496) begin
      FetchL1Plugin_logic_translationStorage_logic_sl_1_write_data_valid = 1'b0;
    end
    case(MmuPlugin_logic_refill_stateReg)
      MmuPlugin_logic_refill_enumDef_IDLE : begin
      end
      MmuPlugin_logic_refill_enumDef_CMD_0 : begin
      end
      MmuPlugin_logic_refill_enumDef_CMD_1 : begin
      end
      MmuPlugin_logic_refill_enumDef_RSP_0 : begin
      end
      MmuPlugin_logic_refill_enumDef_RSP_1 : begin
        if(MmuPlugin_logic_refill_load_rsp_valid) begin
          if(!MmuPlugin_logic_refill_load_rsp_payload_redo) begin
            if(when_MmuPlugin_l471) begin
              FetchL1Plugin_logic_translationStorage_logic_sl_1_write_data_valid = 1'b1;
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    FetchL1Plugin_logic_translationStorage_logic_sl_1_write_data_virtualAddress = 4'bxxxx;
    case(MmuPlugin_logic_refill_stateReg)
      MmuPlugin_logic_refill_enumDef_IDLE : begin
      end
      MmuPlugin_logic_refill_enumDef_CMD_0 : begin
      end
      MmuPlugin_logic_refill_enumDef_CMD_1 : begin
      end
      MmuPlugin_logic_refill_enumDef_RSP_0 : begin
      end
      MmuPlugin_logic_refill_enumDef_RSP_1 : begin
        if(MmuPlugin_logic_refill_load_rsp_valid) begin
          if(!MmuPlugin_logic_refill_load_rsp_payload_redo) begin
            if(when_MmuPlugin_l471) begin
              FetchL1Plugin_logic_translationStorage_logic_sl_1_write_data_virtualAddress = MmuPlugin_logic_refill_virtual[31 : 28];
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    FetchL1Plugin_logic_translationStorage_logic_sl_1_write_data_physicalAddress = 10'bxxxxxxxxxx;
    case(MmuPlugin_logic_refill_stateReg)
      MmuPlugin_logic_refill_enumDef_IDLE : begin
      end
      MmuPlugin_logic_refill_enumDef_CMD_0 : begin
      end
      MmuPlugin_logic_refill_enumDef_CMD_1 : begin
      end
      MmuPlugin_logic_refill_enumDef_RSP_0 : begin
      end
      MmuPlugin_logic_refill_enumDef_RSP_1 : begin
        if(MmuPlugin_logic_refill_load_rsp_valid) begin
          if(!MmuPlugin_logic_refill_load_rsp_payload_redo) begin
            if(when_MmuPlugin_l471) begin
              FetchL1Plugin_logic_translationStorage_logic_sl_1_write_data_physicalAddress = (MmuPlugin_logic_refill_load_levelToPhysicalAddress_1 >>> 5'd22);
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    FetchL1Plugin_logic_translationStorage_logic_sl_1_write_data_allowRead = 1'bx;
    case(MmuPlugin_logic_refill_stateReg)
      MmuPlugin_logic_refill_enumDef_IDLE : begin
      end
      MmuPlugin_logic_refill_enumDef_CMD_0 : begin
      end
      MmuPlugin_logic_refill_enumDef_CMD_1 : begin
      end
      MmuPlugin_logic_refill_enumDef_RSP_0 : begin
      end
      MmuPlugin_logic_refill_enumDef_RSP_1 : begin
        if(MmuPlugin_logic_refill_load_rsp_valid) begin
          if(!MmuPlugin_logic_refill_load_rsp_payload_redo) begin
            if(when_MmuPlugin_l471) begin
              FetchL1Plugin_logic_translationStorage_logic_sl_1_write_data_allowRead = MmuPlugin_logic_refill_load_flags_R;
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    FetchL1Plugin_logic_translationStorage_logic_sl_1_write_data_allowWrite = 1'bx;
    case(MmuPlugin_logic_refill_stateReg)
      MmuPlugin_logic_refill_enumDef_IDLE : begin
      end
      MmuPlugin_logic_refill_enumDef_CMD_0 : begin
      end
      MmuPlugin_logic_refill_enumDef_CMD_1 : begin
      end
      MmuPlugin_logic_refill_enumDef_RSP_0 : begin
      end
      MmuPlugin_logic_refill_enumDef_RSP_1 : begin
        if(MmuPlugin_logic_refill_load_rsp_valid) begin
          if(!MmuPlugin_logic_refill_load_rsp_payload_redo) begin
            if(when_MmuPlugin_l471) begin
              FetchL1Plugin_logic_translationStorage_logic_sl_1_write_data_allowWrite = (MmuPlugin_logic_refill_load_flags_W && MmuPlugin_logic_refill_load_flags_D);
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    FetchL1Plugin_logic_translationStorage_logic_sl_1_write_data_allowExecute = 1'bx;
    case(MmuPlugin_logic_refill_stateReg)
      MmuPlugin_logic_refill_enumDef_IDLE : begin
      end
      MmuPlugin_logic_refill_enumDef_CMD_0 : begin
      end
      MmuPlugin_logic_refill_enumDef_CMD_1 : begin
      end
      MmuPlugin_logic_refill_enumDef_RSP_0 : begin
      end
      MmuPlugin_logic_refill_enumDef_RSP_1 : begin
        if(MmuPlugin_logic_refill_load_rsp_valid) begin
          if(!MmuPlugin_logic_refill_load_rsp_payload_redo) begin
            if(when_MmuPlugin_l471) begin
              FetchL1Plugin_logic_translationStorage_logic_sl_1_write_data_allowExecute = MmuPlugin_logic_refill_load_flags_X;
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    FetchL1Plugin_logic_translationStorage_logic_sl_1_write_data_allowUser = 1'bx;
    case(MmuPlugin_logic_refill_stateReg)
      MmuPlugin_logic_refill_enumDef_IDLE : begin
      end
      MmuPlugin_logic_refill_enumDef_CMD_0 : begin
      end
      MmuPlugin_logic_refill_enumDef_CMD_1 : begin
      end
      MmuPlugin_logic_refill_enumDef_RSP_0 : begin
      end
      MmuPlugin_logic_refill_enumDef_RSP_1 : begin
        if(MmuPlugin_logic_refill_load_rsp_valid) begin
          if(!MmuPlugin_logic_refill_load_rsp_payload_redo) begin
            if(when_MmuPlugin_l471) begin
              FetchL1Plugin_logic_translationStorage_logic_sl_1_write_data_allowUser = MmuPlugin_logic_refill_load_flags_U;
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    FetchL1Plugin_logic_translationStorage_logic_sl_1_allocId_willIncrement = 1'b0;
    case(MmuPlugin_logic_refill_stateReg)
      MmuPlugin_logic_refill_enumDef_IDLE : begin
      end
      MmuPlugin_logic_refill_enumDef_CMD_0 : begin
      end
      MmuPlugin_logic_refill_enumDef_CMD_1 : begin
      end
      MmuPlugin_logic_refill_enumDef_RSP_0 : begin
      end
      MmuPlugin_logic_refill_enumDef_RSP_1 : begin
        if(MmuPlugin_logic_refill_load_rsp_valid) begin
          if(!MmuPlugin_logic_refill_load_rsp_payload_redo) begin
            if(when_MmuPlugin_l471) begin
              FetchL1Plugin_logic_translationStorage_logic_sl_1_allocId_willIncrement = 1'b1;
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  assign FetchL1Plugin_logic_translationStorage_logic_sl_1_allocId_willClear = 1'b0;
  assign FetchL1Plugin_logic_translationStorage_logic_sl_1_allocId_willOverflowIfInc = 1'b1;
  assign FetchL1Plugin_logic_translationStorage_logic_sl_1_allocId_willOverflow = (FetchL1Plugin_logic_translationStorage_logic_sl_1_allocId_willOverflowIfInc && FetchL1Plugin_logic_translationStorage_logic_sl_1_allocId_willIncrement);
  always @(*) begin
    LsuPlugin_logic_translationStorage_logic_sl_0_write_mask = 2'b00;
    if(!when_MmuPlugin_l496) begin
      LsuPlugin_logic_translationStorage_logic_sl_0_write_mask = 2'b11;
    end
    case(MmuPlugin_logic_refill_stateReg)
      MmuPlugin_logic_refill_enumDef_IDLE : begin
      end
      MmuPlugin_logic_refill_enumDef_CMD_0 : begin
      end
      MmuPlugin_logic_refill_enumDef_CMD_1 : begin
      end
      MmuPlugin_logic_refill_enumDef_RSP_0 : begin
        if(MmuPlugin_logic_refill_load_rsp_valid) begin
          if(!MmuPlugin_logic_refill_load_rsp_payload_redo) begin
            LsuPlugin_logic_translationStorage_logic_sl_0_write_mask = (MmuPlugin_logic_refill_storageOhReg[1] ? _zz_LsuPlugin_logic_translationStorage_logic_sl_0_write_mask : 2'b00);
            if(when_MmuPlugin_l439_1) begin
              LsuPlugin_logic_translationStorage_logic_sl_0_write_mask = 2'b00;
            end
          end
        end
      end
      MmuPlugin_logic_refill_enumDef_RSP_1 : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    LsuPlugin_logic_translationStorage_logic_sl_0_write_address = 6'bxxxxxx;
    if(!when_MmuPlugin_l496) begin
      LsuPlugin_logic_translationStorage_logic_sl_0_write_address = MmuPlugin_logic_invalidate_counter;
    end
    case(MmuPlugin_logic_refill_stateReg)
      MmuPlugin_logic_refill_enumDef_IDLE : begin
      end
      MmuPlugin_logic_refill_enumDef_CMD_0 : begin
      end
      MmuPlugin_logic_refill_enumDef_CMD_1 : begin
      end
      MmuPlugin_logic_refill_enumDef_RSP_0 : begin
        if(MmuPlugin_logic_refill_load_rsp_valid) begin
          if(!MmuPlugin_logic_refill_load_rsp_payload_redo) begin
            LsuPlugin_logic_translationStorage_logic_sl_0_write_address = MmuPlugin_logic_refill_virtual[17 : 12];
          end
        end
      end
      MmuPlugin_logic_refill_enumDef_RSP_1 : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    LsuPlugin_logic_translationStorage_logic_sl_0_write_data_valid = 1'bx;
    if(!when_MmuPlugin_l496) begin
      LsuPlugin_logic_translationStorage_logic_sl_0_write_data_valid = 1'b0;
    end
    case(MmuPlugin_logic_refill_stateReg)
      MmuPlugin_logic_refill_enumDef_IDLE : begin
      end
      MmuPlugin_logic_refill_enumDef_CMD_0 : begin
      end
      MmuPlugin_logic_refill_enumDef_CMD_1 : begin
      end
      MmuPlugin_logic_refill_enumDef_RSP_0 : begin
        if(MmuPlugin_logic_refill_load_rsp_valid) begin
          if(!MmuPlugin_logic_refill_load_rsp_payload_redo) begin
            LsuPlugin_logic_translationStorage_logic_sl_0_write_data_valid = 1'b1;
          end
        end
      end
      MmuPlugin_logic_refill_enumDef_RSP_1 : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    LsuPlugin_logic_translationStorage_logic_sl_0_write_data_virtualAddress = 14'bxxxxxxxxxxxxxx;
    case(MmuPlugin_logic_refill_stateReg)
      MmuPlugin_logic_refill_enumDef_IDLE : begin
      end
      MmuPlugin_logic_refill_enumDef_CMD_0 : begin
      end
      MmuPlugin_logic_refill_enumDef_CMD_1 : begin
      end
      MmuPlugin_logic_refill_enumDef_RSP_0 : begin
        if(MmuPlugin_logic_refill_load_rsp_valid) begin
          if(!MmuPlugin_logic_refill_load_rsp_payload_redo) begin
            LsuPlugin_logic_translationStorage_logic_sl_0_write_data_virtualAddress = MmuPlugin_logic_refill_virtual[31 : 18];
          end
        end
      end
      MmuPlugin_logic_refill_enumDef_RSP_1 : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    LsuPlugin_logic_translationStorage_logic_sl_0_write_data_physicalAddress = 20'bxxxxxxxxxxxxxxxxxxxx;
    case(MmuPlugin_logic_refill_stateReg)
      MmuPlugin_logic_refill_enumDef_IDLE : begin
      end
      MmuPlugin_logic_refill_enumDef_CMD_0 : begin
      end
      MmuPlugin_logic_refill_enumDef_CMD_1 : begin
      end
      MmuPlugin_logic_refill_enumDef_RSP_0 : begin
        if(MmuPlugin_logic_refill_load_rsp_valid) begin
          if(!MmuPlugin_logic_refill_load_rsp_payload_redo) begin
            LsuPlugin_logic_translationStorage_logic_sl_0_write_data_physicalAddress = (MmuPlugin_logic_refill_load_levelToPhysicalAddress_0 >>> 4'd12);
          end
        end
      end
      MmuPlugin_logic_refill_enumDef_RSP_1 : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    LsuPlugin_logic_translationStorage_logic_sl_0_write_data_allowRead = 1'bx;
    case(MmuPlugin_logic_refill_stateReg)
      MmuPlugin_logic_refill_enumDef_IDLE : begin
      end
      MmuPlugin_logic_refill_enumDef_CMD_0 : begin
      end
      MmuPlugin_logic_refill_enumDef_CMD_1 : begin
      end
      MmuPlugin_logic_refill_enumDef_RSP_0 : begin
        if(MmuPlugin_logic_refill_load_rsp_valid) begin
          if(!MmuPlugin_logic_refill_load_rsp_payload_redo) begin
            LsuPlugin_logic_translationStorage_logic_sl_0_write_data_allowRead = MmuPlugin_logic_refill_load_flags_R;
          end
        end
      end
      MmuPlugin_logic_refill_enumDef_RSP_1 : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    LsuPlugin_logic_translationStorage_logic_sl_0_write_data_allowWrite = 1'bx;
    case(MmuPlugin_logic_refill_stateReg)
      MmuPlugin_logic_refill_enumDef_IDLE : begin
      end
      MmuPlugin_logic_refill_enumDef_CMD_0 : begin
      end
      MmuPlugin_logic_refill_enumDef_CMD_1 : begin
      end
      MmuPlugin_logic_refill_enumDef_RSP_0 : begin
        if(MmuPlugin_logic_refill_load_rsp_valid) begin
          if(!MmuPlugin_logic_refill_load_rsp_payload_redo) begin
            LsuPlugin_logic_translationStorage_logic_sl_0_write_data_allowWrite = (MmuPlugin_logic_refill_load_flags_W && MmuPlugin_logic_refill_load_flags_D);
          end
        end
      end
      MmuPlugin_logic_refill_enumDef_RSP_1 : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    LsuPlugin_logic_translationStorage_logic_sl_0_write_data_allowExecute = 1'bx;
    case(MmuPlugin_logic_refill_stateReg)
      MmuPlugin_logic_refill_enumDef_IDLE : begin
      end
      MmuPlugin_logic_refill_enumDef_CMD_0 : begin
      end
      MmuPlugin_logic_refill_enumDef_CMD_1 : begin
      end
      MmuPlugin_logic_refill_enumDef_RSP_0 : begin
        if(MmuPlugin_logic_refill_load_rsp_valid) begin
          if(!MmuPlugin_logic_refill_load_rsp_payload_redo) begin
            LsuPlugin_logic_translationStorage_logic_sl_0_write_data_allowExecute = MmuPlugin_logic_refill_load_flags_X;
          end
        end
      end
      MmuPlugin_logic_refill_enumDef_RSP_1 : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    LsuPlugin_logic_translationStorage_logic_sl_0_write_data_allowUser = 1'bx;
    case(MmuPlugin_logic_refill_stateReg)
      MmuPlugin_logic_refill_enumDef_IDLE : begin
      end
      MmuPlugin_logic_refill_enumDef_CMD_0 : begin
      end
      MmuPlugin_logic_refill_enumDef_CMD_1 : begin
      end
      MmuPlugin_logic_refill_enumDef_RSP_0 : begin
        if(MmuPlugin_logic_refill_load_rsp_valid) begin
          if(!MmuPlugin_logic_refill_load_rsp_payload_redo) begin
            LsuPlugin_logic_translationStorage_logic_sl_0_write_data_allowUser = MmuPlugin_logic_refill_load_flags_U;
          end
        end
      end
      MmuPlugin_logic_refill_enumDef_RSP_1 : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    LsuPlugin_logic_translationStorage_logic_sl_0_allocId_willIncrement = 1'b0;
    case(MmuPlugin_logic_refill_stateReg)
      MmuPlugin_logic_refill_enumDef_IDLE : begin
      end
      MmuPlugin_logic_refill_enumDef_CMD_0 : begin
      end
      MmuPlugin_logic_refill_enumDef_CMD_1 : begin
      end
      MmuPlugin_logic_refill_enumDef_RSP_0 : begin
        if(MmuPlugin_logic_refill_load_rsp_valid) begin
          if(!MmuPlugin_logic_refill_load_rsp_payload_redo) begin
            LsuPlugin_logic_translationStorage_logic_sl_0_allocId_willIncrement = 1'b1;
          end
        end
      end
      MmuPlugin_logic_refill_enumDef_RSP_1 : begin
      end
      default : begin
      end
    endcase
  end

  assign LsuPlugin_logic_translationStorage_logic_sl_0_allocId_willClear = 1'b0;
  assign LsuPlugin_logic_translationStorage_logic_sl_0_allocId_willOverflowIfInc = (LsuPlugin_logic_translationStorage_logic_sl_0_allocId_value == 1'b1);
  assign LsuPlugin_logic_translationStorage_logic_sl_0_allocId_willOverflow = (LsuPlugin_logic_translationStorage_logic_sl_0_allocId_willOverflowIfInc && LsuPlugin_logic_translationStorage_logic_sl_0_allocId_willIncrement);
  always @(*) begin
    LsuPlugin_logic_translationStorage_logic_sl_0_allocId_valueNext = (LsuPlugin_logic_translationStorage_logic_sl_0_allocId_value + LsuPlugin_logic_translationStorage_logic_sl_0_allocId_willIncrement);
    if(LsuPlugin_logic_translationStorage_logic_sl_0_allocId_willClear) begin
      LsuPlugin_logic_translationStorage_logic_sl_0_allocId_valueNext = 1'b0;
    end
  end

  always @(*) begin
    LsuPlugin_logic_translationStorage_logic_sl_1_write_mask = 1'b0;
    if(!when_MmuPlugin_l496) begin
      LsuPlugin_logic_translationStorage_logic_sl_1_write_mask = 1'b1;
    end
    case(MmuPlugin_logic_refill_stateReg)
      MmuPlugin_logic_refill_enumDef_IDLE : begin
      end
      MmuPlugin_logic_refill_enumDef_CMD_0 : begin
      end
      MmuPlugin_logic_refill_enumDef_CMD_1 : begin
      end
      MmuPlugin_logic_refill_enumDef_RSP_0 : begin
      end
      MmuPlugin_logic_refill_enumDef_RSP_1 : begin
        if(MmuPlugin_logic_refill_load_rsp_valid) begin
          if(!MmuPlugin_logic_refill_load_rsp_payload_redo) begin
            if(when_MmuPlugin_l471) begin
              LsuPlugin_logic_translationStorage_logic_sl_1_write_mask = (MmuPlugin_logic_refill_storageOhReg[1] ? 1'b1 : 1'b0);
              if(when_MmuPlugin_l439_3) begin
                LsuPlugin_logic_translationStorage_logic_sl_1_write_mask = 1'b0;
              end
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    LsuPlugin_logic_translationStorage_logic_sl_1_write_address = 6'bxxxxxx;
    if(!when_MmuPlugin_l496) begin
      LsuPlugin_logic_translationStorage_logic_sl_1_write_address = MmuPlugin_logic_invalidate_counter;
    end
    case(MmuPlugin_logic_refill_stateReg)
      MmuPlugin_logic_refill_enumDef_IDLE : begin
      end
      MmuPlugin_logic_refill_enumDef_CMD_0 : begin
      end
      MmuPlugin_logic_refill_enumDef_CMD_1 : begin
      end
      MmuPlugin_logic_refill_enumDef_RSP_0 : begin
      end
      MmuPlugin_logic_refill_enumDef_RSP_1 : begin
        if(MmuPlugin_logic_refill_load_rsp_valid) begin
          if(!MmuPlugin_logic_refill_load_rsp_payload_redo) begin
            if(when_MmuPlugin_l471) begin
              LsuPlugin_logic_translationStorage_logic_sl_1_write_address = MmuPlugin_logic_refill_virtual[27 : 22];
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    LsuPlugin_logic_translationStorage_logic_sl_1_write_data_valid = 1'bx;
    if(!when_MmuPlugin_l496) begin
      LsuPlugin_logic_translationStorage_logic_sl_1_write_data_valid = 1'b0;
    end
    case(MmuPlugin_logic_refill_stateReg)
      MmuPlugin_logic_refill_enumDef_IDLE : begin
      end
      MmuPlugin_logic_refill_enumDef_CMD_0 : begin
      end
      MmuPlugin_logic_refill_enumDef_CMD_1 : begin
      end
      MmuPlugin_logic_refill_enumDef_RSP_0 : begin
      end
      MmuPlugin_logic_refill_enumDef_RSP_1 : begin
        if(MmuPlugin_logic_refill_load_rsp_valid) begin
          if(!MmuPlugin_logic_refill_load_rsp_payload_redo) begin
            if(when_MmuPlugin_l471) begin
              LsuPlugin_logic_translationStorage_logic_sl_1_write_data_valid = 1'b1;
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    LsuPlugin_logic_translationStorage_logic_sl_1_write_data_virtualAddress = 4'bxxxx;
    case(MmuPlugin_logic_refill_stateReg)
      MmuPlugin_logic_refill_enumDef_IDLE : begin
      end
      MmuPlugin_logic_refill_enumDef_CMD_0 : begin
      end
      MmuPlugin_logic_refill_enumDef_CMD_1 : begin
      end
      MmuPlugin_logic_refill_enumDef_RSP_0 : begin
      end
      MmuPlugin_logic_refill_enumDef_RSP_1 : begin
        if(MmuPlugin_logic_refill_load_rsp_valid) begin
          if(!MmuPlugin_logic_refill_load_rsp_payload_redo) begin
            if(when_MmuPlugin_l471) begin
              LsuPlugin_logic_translationStorage_logic_sl_1_write_data_virtualAddress = MmuPlugin_logic_refill_virtual[31 : 28];
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    LsuPlugin_logic_translationStorage_logic_sl_1_write_data_physicalAddress = 10'bxxxxxxxxxx;
    case(MmuPlugin_logic_refill_stateReg)
      MmuPlugin_logic_refill_enumDef_IDLE : begin
      end
      MmuPlugin_logic_refill_enumDef_CMD_0 : begin
      end
      MmuPlugin_logic_refill_enumDef_CMD_1 : begin
      end
      MmuPlugin_logic_refill_enumDef_RSP_0 : begin
      end
      MmuPlugin_logic_refill_enumDef_RSP_1 : begin
        if(MmuPlugin_logic_refill_load_rsp_valid) begin
          if(!MmuPlugin_logic_refill_load_rsp_payload_redo) begin
            if(when_MmuPlugin_l471) begin
              LsuPlugin_logic_translationStorage_logic_sl_1_write_data_physicalAddress = (MmuPlugin_logic_refill_load_levelToPhysicalAddress_1 >>> 5'd22);
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    LsuPlugin_logic_translationStorage_logic_sl_1_write_data_allowRead = 1'bx;
    case(MmuPlugin_logic_refill_stateReg)
      MmuPlugin_logic_refill_enumDef_IDLE : begin
      end
      MmuPlugin_logic_refill_enumDef_CMD_0 : begin
      end
      MmuPlugin_logic_refill_enumDef_CMD_1 : begin
      end
      MmuPlugin_logic_refill_enumDef_RSP_0 : begin
      end
      MmuPlugin_logic_refill_enumDef_RSP_1 : begin
        if(MmuPlugin_logic_refill_load_rsp_valid) begin
          if(!MmuPlugin_logic_refill_load_rsp_payload_redo) begin
            if(when_MmuPlugin_l471) begin
              LsuPlugin_logic_translationStorage_logic_sl_1_write_data_allowRead = MmuPlugin_logic_refill_load_flags_R;
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    LsuPlugin_logic_translationStorage_logic_sl_1_write_data_allowWrite = 1'bx;
    case(MmuPlugin_logic_refill_stateReg)
      MmuPlugin_logic_refill_enumDef_IDLE : begin
      end
      MmuPlugin_logic_refill_enumDef_CMD_0 : begin
      end
      MmuPlugin_logic_refill_enumDef_CMD_1 : begin
      end
      MmuPlugin_logic_refill_enumDef_RSP_0 : begin
      end
      MmuPlugin_logic_refill_enumDef_RSP_1 : begin
        if(MmuPlugin_logic_refill_load_rsp_valid) begin
          if(!MmuPlugin_logic_refill_load_rsp_payload_redo) begin
            if(when_MmuPlugin_l471) begin
              LsuPlugin_logic_translationStorage_logic_sl_1_write_data_allowWrite = (MmuPlugin_logic_refill_load_flags_W && MmuPlugin_logic_refill_load_flags_D);
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    LsuPlugin_logic_translationStorage_logic_sl_1_write_data_allowExecute = 1'bx;
    case(MmuPlugin_logic_refill_stateReg)
      MmuPlugin_logic_refill_enumDef_IDLE : begin
      end
      MmuPlugin_logic_refill_enumDef_CMD_0 : begin
      end
      MmuPlugin_logic_refill_enumDef_CMD_1 : begin
      end
      MmuPlugin_logic_refill_enumDef_RSP_0 : begin
      end
      MmuPlugin_logic_refill_enumDef_RSP_1 : begin
        if(MmuPlugin_logic_refill_load_rsp_valid) begin
          if(!MmuPlugin_logic_refill_load_rsp_payload_redo) begin
            if(when_MmuPlugin_l471) begin
              LsuPlugin_logic_translationStorage_logic_sl_1_write_data_allowExecute = MmuPlugin_logic_refill_load_flags_X;
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    LsuPlugin_logic_translationStorage_logic_sl_1_write_data_allowUser = 1'bx;
    case(MmuPlugin_logic_refill_stateReg)
      MmuPlugin_logic_refill_enumDef_IDLE : begin
      end
      MmuPlugin_logic_refill_enumDef_CMD_0 : begin
      end
      MmuPlugin_logic_refill_enumDef_CMD_1 : begin
      end
      MmuPlugin_logic_refill_enumDef_RSP_0 : begin
      end
      MmuPlugin_logic_refill_enumDef_RSP_1 : begin
        if(MmuPlugin_logic_refill_load_rsp_valid) begin
          if(!MmuPlugin_logic_refill_load_rsp_payload_redo) begin
            if(when_MmuPlugin_l471) begin
              LsuPlugin_logic_translationStorage_logic_sl_1_write_data_allowUser = MmuPlugin_logic_refill_load_flags_U;
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    LsuPlugin_logic_translationStorage_logic_sl_1_allocId_willIncrement = 1'b0;
    case(MmuPlugin_logic_refill_stateReg)
      MmuPlugin_logic_refill_enumDef_IDLE : begin
      end
      MmuPlugin_logic_refill_enumDef_CMD_0 : begin
      end
      MmuPlugin_logic_refill_enumDef_CMD_1 : begin
      end
      MmuPlugin_logic_refill_enumDef_RSP_0 : begin
      end
      MmuPlugin_logic_refill_enumDef_RSP_1 : begin
        if(MmuPlugin_logic_refill_load_rsp_valid) begin
          if(!MmuPlugin_logic_refill_load_rsp_payload_redo) begin
            if(when_MmuPlugin_l471) begin
              LsuPlugin_logic_translationStorage_logic_sl_1_allocId_willIncrement = 1'b1;
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  assign LsuPlugin_logic_translationStorage_logic_sl_1_allocId_willClear = 1'b0;
  assign LsuPlugin_logic_translationStorage_logic_sl_1_allocId_willOverflowIfInc = 1'b1;
  assign LsuPlugin_logic_translationStorage_logic_sl_1_allocId_willOverflow = (LsuPlugin_logic_translationStorage_logic_sl_1_allocId_willOverflowIfInc && LsuPlugin_logic_translationStorage_logic_sl_1_allocId_willIncrement);
  assign MmuPlugin_logic_isMachine = (PrivilegedPlugin_logic_harts_0_privilege == 2'b11);
  assign MmuPlugin_logic_isSupervisor = (PrivilegedPlugin_logic_harts_0_privilege == 2'b01);
  assign MmuPlugin_logic_isUser = (PrivilegedPlugin_logic_harts_0_privilege == 2'b00);
  always @(*) begin
    MmuPlugin_api_fetchTranslationEnable = (MmuPlugin_logic_satp_mode == 1'b1);
    if(MmuPlugin_logic_isMachine) begin
      MmuPlugin_api_fetchTranslationEnable = 1'b0;
    end
  end

  always @(*) begin
    MmuPlugin_api_lsuTranslationEnable = (MmuPlugin_logic_satp_mode == 1'b1);
    if(when_MmuPlugin_l264) begin
      MmuPlugin_api_lsuTranslationEnable = 1'b0;
    end
    if(MmuPlugin_logic_isMachine) begin
      if(when_MmuPlugin_l266) begin
        MmuPlugin_api_lsuTranslationEnable = 1'b0;
      end
    end
  end

  assign when_MmuPlugin_l264 = ((! MmuPlugin_logic_status_mprv) && MmuPlugin_logic_isMachine);
  assign when_MmuPlugin_l266 = ((! MmuPlugin_logic_status_mprv) || (PrivilegedPlugin_logic_harts_0_m_status_mpp == 2'b11));
  assign LsuPlugin_logic_onAddress0_translationPort_logic_read_0_readAddress = toplevel_execute_ctrl3_down_LsuL1_MIXED_ADDRESS_lane0[17 : 12];
  assign _zz_toplevel_execute_ctrl3_down_MMU_L0_ENTRIES_lane0_0_valid = LsuPlugin_logic_translationStorage_logic_sl_0_ways_0_spinal_port1;
  assign toplevel_execute_ctrl3_down_MMU_L0_ENTRIES_lane0_0_valid = _zz_toplevel_execute_ctrl3_down_MMU_L0_ENTRIES_lane0_0_valid[0];
  assign toplevel_execute_ctrl3_down_MMU_L0_ENTRIES_lane0_0_virtualAddress = _zz_toplevel_execute_ctrl3_down_MMU_L0_ENTRIES_lane0_0_valid[14 : 1];
  assign toplevel_execute_ctrl3_down_MMU_L0_ENTRIES_lane0_0_physicalAddress = _zz_toplevel_execute_ctrl3_down_MMU_L0_ENTRIES_lane0_0_valid[34 : 15];
  assign toplevel_execute_ctrl3_down_MMU_L0_ENTRIES_lane0_0_allowRead = _zz_toplevel_execute_ctrl3_down_MMU_L0_ENTRIES_lane0_0_valid[35];
  assign toplevel_execute_ctrl3_down_MMU_L0_ENTRIES_lane0_0_allowWrite = _zz_toplevel_execute_ctrl3_down_MMU_L0_ENTRIES_lane0_0_valid[36];
  assign toplevel_execute_ctrl3_down_MMU_L0_ENTRIES_lane0_0_allowExecute = _zz_toplevel_execute_ctrl3_down_MMU_L0_ENTRIES_lane0_0_valid[37];
  assign toplevel_execute_ctrl3_down_MMU_L0_ENTRIES_lane0_0_allowUser = _zz_toplevel_execute_ctrl3_down_MMU_L0_ENTRIES_lane0_0_valid[38];
  always @(*) begin
    toplevel_execute_ctrl3_down_MMU_L0_HITS_PRE_VALID_lane0[0] = (toplevel_execute_ctrl3_down_MMU_L0_ENTRIES_lane0_0_virtualAddress == toplevel_execute_ctrl3_down_LsuL1_MIXED_ADDRESS_lane0[31 : 18]);
    toplevel_execute_ctrl3_down_MMU_L0_HITS_PRE_VALID_lane0[1] = (toplevel_execute_ctrl3_down_MMU_L0_ENTRIES_lane0_1_virtualAddress == toplevel_execute_ctrl3_down_LsuL1_MIXED_ADDRESS_lane0[31 : 18]);
  end

  always @(*) begin
    toplevel_execute_ctrl3_down_MMU_L0_HITS_lane0[0] = (toplevel_execute_ctrl3_down_MMU_L0_HITS_PRE_VALID_lane0[0] && toplevel_execute_ctrl3_down_MMU_L0_ENTRIES_lane0_0_valid);
    toplevel_execute_ctrl3_down_MMU_L0_HITS_lane0[1] = (toplevel_execute_ctrl3_down_MMU_L0_HITS_PRE_VALID_lane0[1] && toplevel_execute_ctrl3_down_MMU_L0_ENTRIES_lane0_1_valid);
  end

  assign _zz_toplevel_execute_ctrl3_down_MMU_L0_ENTRIES_lane0_1_valid = LsuPlugin_logic_translationStorage_logic_sl_0_ways_1_spinal_port1;
  assign toplevel_execute_ctrl3_down_MMU_L0_ENTRIES_lane0_1_valid = _zz_toplevel_execute_ctrl3_down_MMU_L0_ENTRIES_lane0_1_valid[0];
  assign toplevel_execute_ctrl3_down_MMU_L0_ENTRIES_lane0_1_virtualAddress = _zz_toplevel_execute_ctrl3_down_MMU_L0_ENTRIES_lane0_1_valid[14 : 1];
  assign toplevel_execute_ctrl3_down_MMU_L0_ENTRIES_lane0_1_physicalAddress = _zz_toplevel_execute_ctrl3_down_MMU_L0_ENTRIES_lane0_1_valid[34 : 15];
  assign toplevel_execute_ctrl3_down_MMU_L0_ENTRIES_lane0_1_allowRead = _zz_toplevel_execute_ctrl3_down_MMU_L0_ENTRIES_lane0_1_valid[35];
  assign toplevel_execute_ctrl3_down_MMU_L0_ENTRIES_lane0_1_allowWrite = _zz_toplevel_execute_ctrl3_down_MMU_L0_ENTRIES_lane0_1_valid[36];
  assign toplevel_execute_ctrl3_down_MMU_L0_ENTRIES_lane0_1_allowExecute = _zz_toplevel_execute_ctrl3_down_MMU_L0_ENTRIES_lane0_1_valid[37];
  assign toplevel_execute_ctrl3_down_MMU_L0_ENTRIES_lane0_1_allowUser = _zz_toplevel_execute_ctrl3_down_MMU_L0_ENTRIES_lane0_1_valid[38];
  assign LsuPlugin_logic_onAddress0_translationPort_logic_read_1_readAddress = toplevel_execute_ctrl3_down_LsuL1_MIXED_ADDRESS_lane0[27 : 22];
  assign _zz_toplevel_execute_ctrl3_down_MMU_L1_ENTRIES_lane0_0_valid = LsuPlugin_logic_translationStorage_logic_sl_1_ways_0_spinal_port1;
  assign toplevel_execute_ctrl3_down_MMU_L1_ENTRIES_lane0_0_valid = _zz_toplevel_execute_ctrl3_down_MMU_L1_ENTRIES_lane0_0_valid[0];
  assign toplevel_execute_ctrl3_down_MMU_L1_ENTRIES_lane0_0_virtualAddress = _zz_toplevel_execute_ctrl3_down_MMU_L1_ENTRIES_lane0_0_valid[4 : 1];
  assign toplevel_execute_ctrl3_down_MMU_L1_ENTRIES_lane0_0_physicalAddress = _zz_toplevel_execute_ctrl3_down_MMU_L1_ENTRIES_lane0_0_valid[14 : 5];
  assign toplevel_execute_ctrl3_down_MMU_L1_ENTRIES_lane0_0_allowRead = _zz_toplevel_execute_ctrl3_down_MMU_L1_ENTRIES_lane0_0_valid[15];
  assign toplevel_execute_ctrl3_down_MMU_L1_ENTRIES_lane0_0_allowWrite = _zz_toplevel_execute_ctrl3_down_MMU_L1_ENTRIES_lane0_0_valid[16];
  assign toplevel_execute_ctrl3_down_MMU_L1_ENTRIES_lane0_0_allowExecute = _zz_toplevel_execute_ctrl3_down_MMU_L1_ENTRIES_lane0_0_valid[17];
  assign toplevel_execute_ctrl3_down_MMU_L1_ENTRIES_lane0_0_allowUser = _zz_toplevel_execute_ctrl3_down_MMU_L1_ENTRIES_lane0_0_valid[18];
  assign toplevel_execute_ctrl3_down_MMU_L1_HITS_PRE_VALID_lane0[0] = (toplevel_execute_ctrl3_down_MMU_L1_ENTRIES_lane0_0_virtualAddress == toplevel_execute_ctrl3_down_LsuL1_MIXED_ADDRESS_lane0[31 : 28]);
  assign toplevel_execute_ctrl3_down_MMU_L1_HITS_lane0[0] = (toplevel_execute_ctrl3_down_MMU_L1_HITS_PRE_VALID_lane0[0] && toplevel_execute_ctrl3_down_MMU_L1_ENTRIES_lane0_0_valid);
  assign LsuPlugin_logic_onAddress0_translationPort_logic_ctrl_hits = {toplevel_execute_ctrl3_down_MMU_L1_HITS_lane0,toplevel_execute_ctrl3_down_MMU_L0_HITS_lane0};
  assign LsuPlugin_logic_onAddress0_translationPort_logic_ctrl_hit = (|LsuPlugin_logic_onAddress0_translationPort_logic_ctrl_hits);
  assign _zz_LsuPlugin_logic_onAddress0_translationPort_logic_ctrl_hits_bools_0 = LsuPlugin_logic_onAddress0_translationPort_logic_ctrl_hits;
  assign LsuPlugin_logic_onAddress0_translationPort_logic_ctrl_hits_bools_0 = _zz_LsuPlugin_logic_onAddress0_translationPort_logic_ctrl_hits_bools_0[0];
  assign LsuPlugin_logic_onAddress0_translationPort_logic_ctrl_hits_bools_1 = _zz_LsuPlugin_logic_onAddress0_translationPort_logic_ctrl_hits_bools_0[1];
  assign LsuPlugin_logic_onAddress0_translationPort_logic_ctrl_hits_bools_2 = _zz_LsuPlugin_logic_onAddress0_translationPort_logic_ctrl_hits_bools_0[2];
  always @(*) begin
    _zz_LsuPlugin_logic_onAddress0_translationPort_logic_ctrl_oh[0] = (LsuPlugin_logic_onAddress0_translationPort_logic_ctrl_hits_bools_0 && (! 1'b0));
    _zz_LsuPlugin_logic_onAddress0_translationPort_logic_ctrl_oh[1] = (LsuPlugin_logic_onAddress0_translationPort_logic_ctrl_hits_bools_1 && (! LsuPlugin_logic_onAddress0_translationPort_logic_ctrl_hits_bools_0));
    _zz_LsuPlugin_logic_onAddress0_translationPort_logic_ctrl_oh[2] = (LsuPlugin_logic_onAddress0_translationPort_logic_ctrl_hits_bools_2 && (! LsuPlugin_logic_onAddress0_translationPort_logic_ctrl_hits_range_0_to_1));
  end

  assign LsuPlugin_logic_onAddress0_translationPort_logic_ctrl_hits_range_0_to_1 = (|{LsuPlugin_logic_onAddress0_translationPort_logic_ctrl_hits_bools_1,LsuPlugin_logic_onAddress0_translationPort_logic_ctrl_hits_bools_0});
  assign LsuPlugin_logic_onAddress0_translationPort_logic_ctrl_oh = _zz_LsuPlugin_logic_onAddress0_translationPort_logic_ctrl_oh;
  assign _zz_LsuPlugin_logic_onAddress0_translationPort_logic_ctrl_lineAllowExecute = LsuPlugin_logic_onAddress0_translationPort_logic_ctrl_oh[0];
  assign _zz_LsuPlugin_logic_onAddress0_translationPort_logic_ctrl_lineAllowExecute_1 = LsuPlugin_logic_onAddress0_translationPort_logic_ctrl_oh[1];
  assign _zz_LsuPlugin_logic_onAddress0_translationPort_logic_ctrl_lineAllowExecute_2 = LsuPlugin_logic_onAddress0_translationPort_logic_ctrl_oh[2];
  assign LsuPlugin_logic_onAddress0_translationPort_logic_ctrl_lineAllowExecute = _zz_LsuPlugin_logic_onAddress0_translationPort_logic_ctrl_lineAllowExecute_3[0];
  assign LsuPlugin_logic_onAddress0_translationPort_logic_ctrl_lineAllowRead = _zz_LsuPlugin_logic_onAddress0_translationPort_logic_ctrl_lineAllowRead[0];
  assign LsuPlugin_logic_onAddress0_translationPort_logic_ctrl_lineAllowWrite = _zz_LsuPlugin_logic_onAddress0_translationPort_logic_ctrl_lineAllowWrite[0];
  assign LsuPlugin_logic_onAddress0_translationPort_logic_ctrl_lineAllowUser = _zz_LsuPlugin_logic_onAddress0_translationPort_logic_ctrl_lineAllowUser[0];
  assign LsuPlugin_logic_onAddress0_translationPort_logic_ctrl_lineTranslated = (((_zz_LsuPlugin_logic_onAddress0_translationPort_logic_ctrl_lineAllowExecute ? {toplevel_execute_ctrl3_down_MMU_L0_ENTRIES_lane0_0_physicalAddress,_zz_LsuPlugin_logic_onAddress0_translationPort_logic_ctrl_lineTranslated} : 32'h0) | (_zz_LsuPlugin_logic_onAddress0_translationPort_logic_ctrl_lineAllowExecute_1 ? {toplevel_execute_ctrl3_down_MMU_L0_ENTRIES_lane0_1_physicalAddress,_zz_LsuPlugin_logic_onAddress0_translationPort_logic_ctrl_lineTranslated_1} : 32'h0)) | (_zz_LsuPlugin_logic_onAddress0_translationPort_logic_ctrl_lineAllowExecute_2 ? {toplevel_execute_ctrl3_down_MMU_L1_ENTRIES_lane0_0_physicalAddress,toplevel_execute_ctrl3_down_LsuL1_MIXED_ADDRESS_lane0[21 : 0]} : 32'h0));
  always @(*) begin
    LsuPlugin_logic_onAddress0_translationPort_logic_ctrl_requireMmuLockup = MmuPlugin_api_lsuTranslationEnable;
    if(toplevel_execute_ctrl3_down_LsuPlugin_logic_FORCE_PHYSICAL_lane0) begin
      LsuPlugin_logic_onAddress0_translationPort_logic_ctrl_requireMmuLockup = 1'b0;
    end
  end

  always @(*) begin
    if(LsuPlugin_logic_onAddress0_translationPort_logic_ctrl_requireMmuLockup) begin
      toplevel_execute_ctrl3_down_MMU_HAZARD_lane0 = 1'b0;
    end else begin
      toplevel_execute_ctrl3_down_MMU_HAZARD_lane0 = 1'b0;
    end
  end

  always @(*) begin
    if(LsuPlugin_logic_onAddress0_translationPort_logic_ctrl_requireMmuLockup) begin
      toplevel_execute_ctrl3_down_MMU_REFILL_lane0 = (! LsuPlugin_logic_onAddress0_translationPort_logic_ctrl_hit);
    end else begin
      toplevel_execute_ctrl3_down_MMU_REFILL_lane0 = 1'b0;
    end
  end

  always @(*) begin
    if(LsuPlugin_logic_onAddress0_translationPort_logic_ctrl_requireMmuLockup) begin
      toplevel_execute_ctrl3_down_MMU_TRANSLATED_lane0 = LsuPlugin_logic_onAddress0_translationPort_logic_ctrl_lineTranslated;
    end else begin
      toplevel_execute_ctrl3_down_MMU_TRANSLATED_lane0 = toplevel_execute_ctrl3_down_LsuL1_MIXED_ADDRESS_lane0;
    end
  end

  always @(*) begin
    if(LsuPlugin_logic_onAddress0_translationPort_logic_ctrl_requireMmuLockup) begin
      toplevel_execute_ctrl3_down_MMU_ALLOW_EXECUTE_lane0 = (LsuPlugin_logic_onAddress0_translationPort_logic_ctrl_lineAllowExecute && (! (LsuPlugin_logic_onAddress0_translationPort_logic_ctrl_lineAllowUser && MmuPlugin_logic_isSupervisor)));
    end else begin
      toplevel_execute_ctrl3_down_MMU_ALLOW_EXECUTE_lane0 = 1'b1;
    end
  end

  always @(*) begin
    if(LsuPlugin_logic_onAddress0_translationPort_logic_ctrl_requireMmuLockup) begin
      toplevel_execute_ctrl3_down_MMU_ALLOW_READ_lane0 = (LsuPlugin_logic_onAddress0_translationPort_logic_ctrl_lineAllowRead || (MmuPlugin_logic_status_mxr && LsuPlugin_logic_onAddress0_translationPort_logic_ctrl_lineAllowExecute));
    end else begin
      toplevel_execute_ctrl3_down_MMU_ALLOW_READ_lane0 = 1'b1;
    end
  end

  always @(*) begin
    if(LsuPlugin_logic_onAddress0_translationPort_logic_ctrl_requireMmuLockup) begin
      toplevel_execute_ctrl3_down_MMU_ALLOW_WRITE_lane0 = LsuPlugin_logic_onAddress0_translationPort_logic_ctrl_lineAllowWrite;
    end else begin
      toplevel_execute_ctrl3_down_MMU_ALLOW_WRITE_lane0 = 1'b1;
    end
  end

  always @(*) begin
    if(LsuPlugin_logic_onAddress0_translationPort_logic_ctrl_requireMmuLockup) begin
      toplevel_execute_ctrl3_down_MMU_PAGE_FAULT_lane0 = (((LsuPlugin_logic_onAddress0_translationPort_logic_ctrl_lineAllowUser && MmuPlugin_logic_isSupervisor) && (! MmuPlugin_logic_status_sum)) || ((! LsuPlugin_logic_onAddress0_translationPort_logic_ctrl_lineAllowUser) && MmuPlugin_logic_isUser));
    end else begin
      toplevel_execute_ctrl3_down_MMU_PAGE_FAULT_lane0 = 1'b0;
    end
  end

  always @(*) begin
    if(LsuPlugin_logic_onAddress0_translationPort_logic_ctrl_requireMmuLockup) begin
      toplevel_execute_ctrl3_down_MMU_ACCESS_FAULT_lane0 = 1'b0;
    end else begin
      toplevel_execute_ctrl3_down_MMU_ACCESS_FAULT_lane0 = 1'b0;
    end
  end

  assign toplevel_execute_ctrl3_down_MMU_BYPASS_TRANSLATION_lane0 = (! LsuPlugin_logic_onAddress0_translationPort_logic_ctrl_requireMmuLockup);
  assign toplevel_execute_ctrl3_down_MMU_WAYS_OH_lane0 = LsuPlugin_logic_onAddress0_translationPort_logic_ctrl_oh;
  assign toplevel_execute_ctrl3_down_MMU_WAYS_PHYSICAL_lane0_0 = {toplevel_execute_ctrl3_down_MMU_L0_ENTRIES_lane0_0_physicalAddress,toplevel_execute_ctrl3_down_LsuL1_MIXED_ADDRESS_lane0[11 : 0]};
  assign toplevel_execute_ctrl3_down_MMU_WAYS_PHYSICAL_lane0_1 = {toplevel_execute_ctrl3_down_MMU_L0_ENTRIES_lane0_1_physicalAddress,toplevel_execute_ctrl3_down_LsuL1_MIXED_ADDRESS_lane0[11 : 0]};
  assign toplevel_execute_ctrl3_down_MMU_WAYS_PHYSICAL_lane0_2 = {toplevel_execute_ctrl3_down_MMU_L1_ENTRIES_lane0_0_physicalAddress,toplevel_execute_ctrl3_down_LsuL1_MIXED_ADDRESS_lane0[21 : 0]};
  assign FetchL1Plugin_logic_translationPort_logic_read_0_readAddress = fetch_logic_ctrls_1_down_Fetch_WORD_PC[17 : 12];
  assign _zz_fetch_logic_ctrls_1_down_MMU_L0_ENTRIES_0_valid = FetchL1Plugin_logic_translationStorage_logic_sl_0_ways_0_spinal_port1;
  assign fetch_logic_ctrls_1_down_MMU_L0_ENTRIES_0_valid = _zz_fetch_logic_ctrls_1_down_MMU_L0_ENTRIES_0_valid[0];
  assign fetch_logic_ctrls_1_down_MMU_L0_ENTRIES_0_virtualAddress = _zz_fetch_logic_ctrls_1_down_MMU_L0_ENTRIES_0_valid[14 : 1];
  assign fetch_logic_ctrls_1_down_MMU_L0_ENTRIES_0_physicalAddress = _zz_fetch_logic_ctrls_1_down_MMU_L0_ENTRIES_0_valid[34 : 15];
  assign fetch_logic_ctrls_1_down_MMU_L0_ENTRIES_0_allowRead = _zz_fetch_logic_ctrls_1_down_MMU_L0_ENTRIES_0_valid[35];
  assign fetch_logic_ctrls_1_down_MMU_L0_ENTRIES_0_allowWrite = _zz_fetch_logic_ctrls_1_down_MMU_L0_ENTRIES_0_valid[36];
  assign fetch_logic_ctrls_1_down_MMU_L0_ENTRIES_0_allowExecute = _zz_fetch_logic_ctrls_1_down_MMU_L0_ENTRIES_0_valid[37];
  assign fetch_logic_ctrls_1_down_MMU_L0_ENTRIES_0_allowUser = _zz_fetch_logic_ctrls_1_down_MMU_L0_ENTRIES_0_valid[38];
  always @(*) begin
    fetch_logic_ctrls_1_down_MMU_L0_HITS_PRE_VALID[0] = (fetch_logic_ctrls_1_down_MMU_L0_ENTRIES_0_virtualAddress == fetch_logic_ctrls_1_down_Fetch_WORD_PC[31 : 18]);
    fetch_logic_ctrls_1_down_MMU_L0_HITS_PRE_VALID[1] = (fetch_logic_ctrls_1_down_MMU_L0_ENTRIES_1_virtualAddress == fetch_logic_ctrls_1_down_Fetch_WORD_PC[31 : 18]);
  end

  always @(*) begin
    fetch_logic_ctrls_1_down_MMU_L0_HITS[0] = (fetch_logic_ctrls_1_down_MMU_L0_HITS_PRE_VALID[0] && fetch_logic_ctrls_1_down_MMU_L0_ENTRIES_0_valid);
    fetch_logic_ctrls_1_down_MMU_L0_HITS[1] = (fetch_logic_ctrls_1_down_MMU_L0_HITS_PRE_VALID[1] && fetch_logic_ctrls_1_down_MMU_L0_ENTRIES_1_valid);
  end

  assign _zz_fetch_logic_ctrls_1_down_MMU_L0_ENTRIES_1_valid = FetchL1Plugin_logic_translationStorage_logic_sl_0_ways_1_spinal_port1;
  assign fetch_logic_ctrls_1_down_MMU_L0_ENTRIES_1_valid = _zz_fetch_logic_ctrls_1_down_MMU_L0_ENTRIES_1_valid[0];
  assign fetch_logic_ctrls_1_down_MMU_L0_ENTRIES_1_virtualAddress = _zz_fetch_logic_ctrls_1_down_MMU_L0_ENTRIES_1_valid[14 : 1];
  assign fetch_logic_ctrls_1_down_MMU_L0_ENTRIES_1_physicalAddress = _zz_fetch_logic_ctrls_1_down_MMU_L0_ENTRIES_1_valid[34 : 15];
  assign fetch_logic_ctrls_1_down_MMU_L0_ENTRIES_1_allowRead = _zz_fetch_logic_ctrls_1_down_MMU_L0_ENTRIES_1_valid[35];
  assign fetch_logic_ctrls_1_down_MMU_L0_ENTRIES_1_allowWrite = _zz_fetch_logic_ctrls_1_down_MMU_L0_ENTRIES_1_valid[36];
  assign fetch_logic_ctrls_1_down_MMU_L0_ENTRIES_1_allowExecute = _zz_fetch_logic_ctrls_1_down_MMU_L0_ENTRIES_1_valid[37];
  assign fetch_logic_ctrls_1_down_MMU_L0_ENTRIES_1_allowUser = _zz_fetch_logic_ctrls_1_down_MMU_L0_ENTRIES_1_valid[38];
  assign FetchL1Plugin_logic_translationPort_logic_read_1_readAddress = fetch_logic_ctrls_1_down_Fetch_WORD_PC[27 : 22];
  assign _zz_fetch_logic_ctrls_1_down_MMU_L1_ENTRIES_0_valid = FetchL1Plugin_logic_translationStorage_logic_sl_1_ways_0_spinal_port1;
  assign fetch_logic_ctrls_1_down_MMU_L1_ENTRIES_0_valid = _zz_fetch_logic_ctrls_1_down_MMU_L1_ENTRIES_0_valid[0];
  assign fetch_logic_ctrls_1_down_MMU_L1_ENTRIES_0_virtualAddress = _zz_fetch_logic_ctrls_1_down_MMU_L1_ENTRIES_0_valid[4 : 1];
  assign fetch_logic_ctrls_1_down_MMU_L1_ENTRIES_0_physicalAddress = _zz_fetch_logic_ctrls_1_down_MMU_L1_ENTRIES_0_valid[14 : 5];
  assign fetch_logic_ctrls_1_down_MMU_L1_ENTRIES_0_allowRead = _zz_fetch_logic_ctrls_1_down_MMU_L1_ENTRIES_0_valid[15];
  assign fetch_logic_ctrls_1_down_MMU_L1_ENTRIES_0_allowWrite = _zz_fetch_logic_ctrls_1_down_MMU_L1_ENTRIES_0_valid[16];
  assign fetch_logic_ctrls_1_down_MMU_L1_ENTRIES_0_allowExecute = _zz_fetch_logic_ctrls_1_down_MMU_L1_ENTRIES_0_valid[17];
  assign fetch_logic_ctrls_1_down_MMU_L1_ENTRIES_0_allowUser = _zz_fetch_logic_ctrls_1_down_MMU_L1_ENTRIES_0_valid[18];
  assign fetch_logic_ctrls_1_down_MMU_L1_HITS_PRE_VALID[0] = (fetch_logic_ctrls_1_down_MMU_L1_ENTRIES_0_virtualAddress == fetch_logic_ctrls_1_down_Fetch_WORD_PC[31 : 28]);
  assign fetch_logic_ctrls_1_down_MMU_L1_HITS[0] = (fetch_logic_ctrls_1_down_MMU_L1_HITS_PRE_VALID[0] && fetch_logic_ctrls_1_down_MMU_L1_ENTRIES_0_valid);
  assign FetchL1Plugin_logic_translationPort_logic_ctrl_hits = {fetch_logic_ctrls_1_down_MMU_L1_HITS,fetch_logic_ctrls_1_down_MMU_L0_HITS};
  assign FetchL1Plugin_logic_translationPort_logic_ctrl_hit = (|FetchL1Plugin_logic_translationPort_logic_ctrl_hits);
  assign _zz_FetchL1Plugin_logic_translationPort_logic_ctrl_hits_bools_0 = FetchL1Plugin_logic_translationPort_logic_ctrl_hits;
  assign FetchL1Plugin_logic_translationPort_logic_ctrl_hits_bools_0 = _zz_FetchL1Plugin_logic_translationPort_logic_ctrl_hits_bools_0[0];
  assign FetchL1Plugin_logic_translationPort_logic_ctrl_hits_bools_1 = _zz_FetchL1Plugin_logic_translationPort_logic_ctrl_hits_bools_0[1];
  assign FetchL1Plugin_logic_translationPort_logic_ctrl_hits_bools_2 = _zz_FetchL1Plugin_logic_translationPort_logic_ctrl_hits_bools_0[2];
  always @(*) begin
    _zz_FetchL1Plugin_logic_translationPort_logic_ctrl_oh[0] = (FetchL1Plugin_logic_translationPort_logic_ctrl_hits_bools_0 && (! 1'b0));
    _zz_FetchL1Plugin_logic_translationPort_logic_ctrl_oh[1] = (FetchL1Plugin_logic_translationPort_logic_ctrl_hits_bools_1 && (! FetchL1Plugin_logic_translationPort_logic_ctrl_hits_bools_0));
    _zz_FetchL1Plugin_logic_translationPort_logic_ctrl_oh[2] = (FetchL1Plugin_logic_translationPort_logic_ctrl_hits_bools_2 && (! FetchL1Plugin_logic_translationPort_logic_ctrl_hits_range_0_to_1));
  end

  assign FetchL1Plugin_logic_translationPort_logic_ctrl_hits_range_0_to_1 = (|{FetchL1Plugin_logic_translationPort_logic_ctrl_hits_bools_1,FetchL1Plugin_logic_translationPort_logic_ctrl_hits_bools_0});
  assign FetchL1Plugin_logic_translationPort_logic_ctrl_oh = _zz_FetchL1Plugin_logic_translationPort_logic_ctrl_oh;
  assign _zz_FetchL1Plugin_logic_translationPort_logic_ctrl_lineAllowExecute = FetchL1Plugin_logic_translationPort_logic_ctrl_oh[0];
  assign _zz_FetchL1Plugin_logic_translationPort_logic_ctrl_lineAllowExecute_1 = FetchL1Plugin_logic_translationPort_logic_ctrl_oh[1];
  assign _zz_FetchL1Plugin_logic_translationPort_logic_ctrl_lineAllowExecute_2 = FetchL1Plugin_logic_translationPort_logic_ctrl_oh[2];
  assign FetchL1Plugin_logic_translationPort_logic_ctrl_lineAllowExecute = _zz_FetchL1Plugin_logic_translationPort_logic_ctrl_lineAllowExecute_3[0];
  assign FetchL1Plugin_logic_translationPort_logic_ctrl_lineAllowRead = _zz_FetchL1Plugin_logic_translationPort_logic_ctrl_lineAllowRead[0];
  assign FetchL1Plugin_logic_translationPort_logic_ctrl_lineAllowWrite = _zz_FetchL1Plugin_logic_translationPort_logic_ctrl_lineAllowWrite[0];
  assign FetchL1Plugin_logic_translationPort_logic_ctrl_lineAllowUser = _zz_FetchL1Plugin_logic_translationPort_logic_ctrl_lineAllowUser[0];
  assign FetchL1Plugin_logic_translationPort_logic_ctrl_lineTranslated = (((_zz_FetchL1Plugin_logic_translationPort_logic_ctrl_lineAllowExecute ? {fetch_logic_ctrls_1_down_MMU_L0_ENTRIES_0_physicalAddress,_zz_FetchL1Plugin_logic_translationPort_logic_ctrl_lineTranslated} : 32'h0) | (_zz_FetchL1Plugin_logic_translationPort_logic_ctrl_lineAllowExecute_1 ? {fetch_logic_ctrls_1_down_MMU_L0_ENTRIES_1_physicalAddress,_zz_FetchL1Plugin_logic_translationPort_logic_ctrl_lineTranslated_1} : 32'h0)) | (_zz_FetchL1Plugin_logic_translationPort_logic_ctrl_lineAllowExecute_2 ? {fetch_logic_ctrls_1_down_MMU_L1_ENTRIES_0_physicalAddress,fetch_logic_ctrls_1_down_Fetch_WORD_PC[21 : 0]} : 32'h0));
  always @(*) begin
    FetchL1Plugin_logic_translationPort_logic_ctrl_requireMmuLockup = MmuPlugin_api_fetchTranslationEnable;
    if(_zz_1) begin
      FetchL1Plugin_logic_translationPort_logic_ctrl_requireMmuLockup = 1'b0;
    end
  end

  always @(*) begin
    if(FetchL1Plugin_logic_translationPort_logic_ctrl_requireMmuLockup) begin
      fetch_logic_ctrls_1_down_MMU_HAZARD = 1'b0;
    end else begin
      fetch_logic_ctrls_1_down_MMU_HAZARD = 1'b0;
    end
  end

  always @(*) begin
    if(FetchL1Plugin_logic_translationPort_logic_ctrl_requireMmuLockup) begin
      fetch_logic_ctrls_1_down_MMU_REFILL = (! FetchL1Plugin_logic_translationPort_logic_ctrl_hit);
    end else begin
      fetch_logic_ctrls_1_down_MMU_REFILL = 1'b0;
    end
  end

  always @(*) begin
    if(FetchL1Plugin_logic_translationPort_logic_ctrl_requireMmuLockup) begin
      fetch_logic_ctrls_1_down_MMU_TRANSLATED = FetchL1Plugin_logic_translationPort_logic_ctrl_lineTranslated;
    end else begin
      fetch_logic_ctrls_1_down_MMU_TRANSLATED = fetch_logic_ctrls_1_down_Fetch_WORD_PC;
    end
  end

  always @(*) begin
    if(FetchL1Plugin_logic_translationPort_logic_ctrl_requireMmuLockup) begin
      fetch_logic_ctrls_1_down_MMU_ALLOW_EXECUTE = (FetchL1Plugin_logic_translationPort_logic_ctrl_lineAllowExecute && (! (FetchL1Plugin_logic_translationPort_logic_ctrl_lineAllowUser && MmuPlugin_logic_isSupervisor)));
    end else begin
      fetch_logic_ctrls_1_down_MMU_ALLOW_EXECUTE = 1'b1;
    end
  end

  always @(*) begin
    if(FetchL1Plugin_logic_translationPort_logic_ctrl_requireMmuLockup) begin
      fetch_logic_ctrls_1_down_MMU_ALLOW_READ = (FetchL1Plugin_logic_translationPort_logic_ctrl_lineAllowRead || (MmuPlugin_logic_status_mxr && FetchL1Plugin_logic_translationPort_logic_ctrl_lineAllowExecute));
    end else begin
      fetch_logic_ctrls_1_down_MMU_ALLOW_READ = 1'b1;
    end
  end

  always @(*) begin
    if(FetchL1Plugin_logic_translationPort_logic_ctrl_requireMmuLockup) begin
      fetch_logic_ctrls_1_down_MMU_ALLOW_WRITE = FetchL1Plugin_logic_translationPort_logic_ctrl_lineAllowWrite;
    end else begin
      fetch_logic_ctrls_1_down_MMU_ALLOW_WRITE = 1'b1;
    end
  end

  always @(*) begin
    if(FetchL1Plugin_logic_translationPort_logic_ctrl_requireMmuLockup) begin
      fetch_logic_ctrls_1_down_MMU_PAGE_FAULT = (((FetchL1Plugin_logic_translationPort_logic_ctrl_lineAllowUser && MmuPlugin_logic_isSupervisor) && (! MmuPlugin_logic_status_sum)) || ((! FetchL1Plugin_logic_translationPort_logic_ctrl_lineAllowUser) && MmuPlugin_logic_isUser));
    end else begin
      fetch_logic_ctrls_1_down_MMU_PAGE_FAULT = 1'b0;
    end
  end

  always @(*) begin
    if(FetchL1Plugin_logic_translationPort_logic_ctrl_requireMmuLockup) begin
      fetch_logic_ctrls_1_down_MMU_ACCESS_FAULT = 1'b0;
    end else begin
      fetch_logic_ctrls_1_down_MMU_ACCESS_FAULT = 1'b0;
    end
  end

  assign fetch_logic_ctrls_1_down_MMU_BYPASS_TRANSLATION = (! FetchL1Plugin_logic_translationPort_logic_ctrl_requireMmuLockup);
  assign fetch_logic_ctrls_1_down_MMU_WAYS_OH = FetchL1Plugin_logic_translationPort_logic_ctrl_oh;
  assign fetch_logic_ctrls_1_down_MMU_WAYS_PHYSICAL_0 = {fetch_logic_ctrls_1_down_MMU_L0_ENTRIES_0_physicalAddress,fetch_logic_ctrls_1_down_Fetch_WORD_PC[11 : 0]};
  assign fetch_logic_ctrls_1_down_MMU_WAYS_PHYSICAL_1 = {fetch_logic_ctrls_1_down_MMU_L0_ENTRIES_1_physicalAddress,fetch_logic_ctrls_1_down_Fetch_WORD_PC[11 : 0]};
  assign fetch_logic_ctrls_1_down_MMU_WAYS_PHYSICAL_2 = {fetch_logic_ctrls_1_down_MMU_L1_ENTRIES_0_physicalAddress,fetch_logic_ctrls_1_down_Fetch_WORD_PC[21 : 0]};
  assign MmuPlugin_logic_refill_wantExit = 1'b0;
  always @(*) begin
    MmuPlugin_logic_refill_wantStart = 1'b0;
    case(MmuPlugin_logic_refill_stateReg)
      MmuPlugin_logic_refill_enumDef_IDLE : begin
      end
      MmuPlugin_logic_refill_enumDef_CMD_0 : begin
      end
      MmuPlugin_logic_refill_enumDef_CMD_1 : begin
      end
      MmuPlugin_logic_refill_enumDef_RSP_0 : begin
      end
      MmuPlugin_logic_refill_enumDef_RSP_1 : begin
      end
      default : begin
        MmuPlugin_logic_refill_wantStart = 1'b1;
      end
    endcase
  end

  assign MmuPlugin_logic_refill_wantKill = 1'b0;
  assign MmuPlugin_logic_refill_busy = (! (MmuPlugin_logic_refill_stateReg == MmuPlugin_logic_refill_enumDef_IDLE));
  always @(*) begin
    MmuPlugin_logic_refill_cacheRefillAnySet = 1'b0;
    if(when_MmuPlugin_l383) begin
      MmuPlugin_logic_refill_cacheRefillAnySet = MmuPlugin_logic_accessBus_rsp_payload_waitAny;
    end
  end

  assign TrapPlugin_logic_harts_0_trap_fsm_atsPorts_refill_cmd_ready = MmuPlugin_logic_refill_arbiter_io_inputs_0_ready;
  always @(*) begin
    MmuPlugin_logic_refill_arbiter_io_output_ready = 1'b0;
    case(MmuPlugin_logic_refill_stateReg)
      MmuPlugin_logic_refill_enumDef_IDLE : begin
        if(MmuPlugin_logic_refill_arbiter_io_output_valid) begin
          MmuPlugin_logic_refill_arbiter_io_output_ready = 1'b1;
        end
      end
      MmuPlugin_logic_refill_enumDef_CMD_0 : begin
      end
      MmuPlugin_logic_refill_enumDef_CMD_1 : begin
      end
      MmuPlugin_logic_refill_enumDef_RSP_0 : begin
      end
      MmuPlugin_logic_refill_enumDef_RSP_1 : begin
      end
      default : begin
      end
    endcase
  end

  assign MmuPlugin_logic_refill_load_readed = MmuPlugin_logic_refill_load_rsp_payload_data[31 : 0];
  assign when_MmuPlugin_l383 = (MmuPlugin_logic_accessBus_rsp_valid && MmuPlugin_logic_accessBus_rsp_payload_redo);
  always @(*) begin
    MmuPlugin_logic_accessBus_cmd_valid = 1'b0;
    case(MmuPlugin_logic_refill_stateReg)
      MmuPlugin_logic_refill_enumDef_IDLE : begin
      end
      MmuPlugin_logic_refill_enumDef_CMD_0 : begin
        if(when_MmuPlugin_l454) begin
          MmuPlugin_logic_accessBus_cmd_valid = 1'b1;
        end
      end
      MmuPlugin_logic_refill_enumDef_CMD_1 : begin
        if(when_MmuPlugin_l454_1) begin
          MmuPlugin_logic_accessBus_cmd_valid = 1'b1;
        end
      end
      MmuPlugin_logic_refill_enumDef_RSP_0 : begin
      end
      MmuPlugin_logic_refill_enumDef_RSP_1 : begin
      end
      default : begin
      end
    endcase
  end

  assign MmuPlugin_logic_accessBus_cmd_payload_address = MmuPlugin_logic_refill_load_address;
  assign MmuPlugin_logic_accessBus_cmd_payload_size = 2'b10;
  assign _zz_MmuPlugin_logic_refill_load_flags_V = MmuPlugin_logic_refill_load_readed;
  assign MmuPlugin_logic_refill_load_flags_V = _zz_MmuPlugin_logic_refill_load_flags_V[0];
  assign MmuPlugin_logic_refill_load_flags_R = _zz_MmuPlugin_logic_refill_load_flags_V[1];
  assign MmuPlugin_logic_refill_load_flags_W = _zz_MmuPlugin_logic_refill_load_flags_V[2];
  assign MmuPlugin_logic_refill_load_flags_X = _zz_MmuPlugin_logic_refill_load_flags_V[3];
  assign MmuPlugin_logic_refill_load_flags_U = _zz_MmuPlugin_logic_refill_load_flags_V[4];
  assign MmuPlugin_logic_refill_load_flags_G = _zz_MmuPlugin_logic_refill_load_flags_V[5];
  assign MmuPlugin_logic_refill_load_flags_A = _zz_MmuPlugin_logic_refill_load_flags_V[6];
  assign MmuPlugin_logic_refill_load_flags_D = _zz_MmuPlugin_logic_refill_load_flags_V[7];
  assign MmuPlugin_logic_refill_load_leaf = (MmuPlugin_logic_refill_load_flags_R || MmuPlugin_logic_refill_load_flags_X);
  always @(*) begin
    MmuPlugin_logic_refill_load_exception = ((((! MmuPlugin_logic_refill_load_flags_V) || ((! MmuPlugin_logic_refill_load_flags_R) && MmuPlugin_logic_refill_load_flags_W)) || MmuPlugin_logic_refill_load_rsp_payload_error) || ((! MmuPlugin_logic_refill_load_leaf) && ((MmuPlugin_logic_refill_load_flags_D || MmuPlugin_logic_refill_load_flags_A) || MmuPlugin_logic_refill_load_flags_U)));
    case(MmuPlugin_logic_refill_stateReg)
      MmuPlugin_logic_refill_enumDef_IDLE : begin
      end
      MmuPlugin_logic_refill_enumDef_CMD_0 : begin
      end
      MmuPlugin_logic_refill_enumDef_CMD_1 : begin
      end
      MmuPlugin_logic_refill_enumDef_RSP_0 : begin
        if(when_MmuPlugin_l463) begin
          MmuPlugin_logic_refill_load_exception = 1'b1;
        end
      end
      MmuPlugin_logic_refill_enumDef_RSP_1 : begin
      end
      default : begin
      end
    endcase
  end

  assign MmuPlugin_logic_refill_load_levelException_0 = 1'b0;
  always @(*) begin
    MmuPlugin_logic_refill_load_levelException_1 = 1'b0;
    if(when_MmuPlugin_l403) begin
      MmuPlugin_logic_refill_load_levelException_1 = 1'b1;
    end
  end

  always @(*) begin
    MmuPlugin_logic_refill_load_nextLevelBase = 32'h0;
    MmuPlugin_logic_refill_load_nextLevelBase[21 : 12] = MmuPlugin_logic_refill_load_readed[19 : 10];
    MmuPlugin_logic_refill_load_nextLevelBase[31 : 22] = MmuPlugin_logic_refill_load_readed[29 : 20];
  end

  always @(*) begin
    MmuPlugin_logic_refill_load_levelToPhysicalAddress_0 = 32'h0;
    MmuPlugin_logic_refill_load_levelToPhysicalAddress_0[21 : 12] = MmuPlugin_logic_refill_load_readed[19 : 10];
    MmuPlugin_logic_refill_load_levelToPhysicalAddress_0[31 : 22] = MmuPlugin_logic_refill_load_readed[29 : 20];
  end

  always @(*) begin
    MmuPlugin_logic_refill_load_levelToPhysicalAddress_1 = 32'h0;
    MmuPlugin_logic_refill_load_levelToPhysicalAddress_1[21 : 12] = MmuPlugin_logic_refill_virtual[21 : 12];
    MmuPlugin_logic_refill_load_levelToPhysicalAddress_1[31 : 22] = MmuPlugin_logic_refill_load_readed[29 : 20];
  end

  assign when_MmuPlugin_l403 = (MmuPlugin_logic_refill_load_readed[19 : 10] != 10'h0);
  always @(*) begin
    TrapPlugin_logic_harts_0_trap_fsm_atsPorts_refill_rsp_valid = 1'b0;
    case(MmuPlugin_logic_refill_stateReg)
      MmuPlugin_logic_refill_enumDef_IDLE : begin
      end
      MmuPlugin_logic_refill_enumDef_CMD_0 : begin
      end
      MmuPlugin_logic_refill_enumDef_CMD_1 : begin
      end
      MmuPlugin_logic_refill_enumDef_RSP_0 : begin
        if(MmuPlugin_logic_refill_load_rsp_valid) begin
          if(!MmuPlugin_logic_refill_load_rsp_payload_redo) begin
            if(_zz_54) begin
              TrapPlugin_logic_harts_0_trap_fsm_atsPorts_refill_rsp_valid = 1'b1;
            end
            if(_zz_54) begin
              TrapPlugin_logic_harts_0_trap_fsm_atsPorts_refill_rsp_valid = 1'b1;
            end
          end
        end
      end
      MmuPlugin_logic_refill_enumDef_RSP_1 : begin
        if(MmuPlugin_logic_refill_load_rsp_valid) begin
          if(!MmuPlugin_logic_refill_load_rsp_payload_redo) begin
            if(when_MmuPlugin_l471) begin
              if(_zz_54) begin
                TrapPlugin_logic_harts_0_trap_fsm_atsPorts_refill_rsp_valid = 1'b1;
              end
              if(_zz_54) begin
                TrapPlugin_logic_harts_0_trap_fsm_atsPorts_refill_rsp_valid = 1'b1;
              end
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    TrapPlugin_logic_harts_0_trap_fsm_atsPorts_refill_rsp_payload_pageFault = 1'bx;
    case(MmuPlugin_logic_refill_stateReg)
      MmuPlugin_logic_refill_enumDef_IDLE : begin
      end
      MmuPlugin_logic_refill_enumDef_CMD_0 : begin
      end
      MmuPlugin_logic_refill_enumDef_CMD_1 : begin
      end
      MmuPlugin_logic_refill_enumDef_RSP_0 : begin
        if(MmuPlugin_logic_refill_load_rsp_valid) begin
          if(!MmuPlugin_logic_refill_load_rsp_payload_redo) begin
            if(_zz_54) begin
              TrapPlugin_logic_harts_0_trap_fsm_atsPorts_refill_rsp_payload_pageFault = MmuPlugin_logic_refill_fetch_0_pageFault;
            end
            if(_zz_54) begin
              TrapPlugin_logic_harts_0_trap_fsm_atsPorts_refill_rsp_payload_pageFault = MmuPlugin_logic_refill_fetch_0_pageFault;
            end
          end
        end
      end
      MmuPlugin_logic_refill_enumDef_RSP_1 : begin
        if(MmuPlugin_logic_refill_load_rsp_valid) begin
          if(!MmuPlugin_logic_refill_load_rsp_payload_redo) begin
            if(when_MmuPlugin_l471) begin
              if(_zz_54) begin
                TrapPlugin_logic_harts_0_trap_fsm_atsPorts_refill_rsp_payload_pageFault = MmuPlugin_logic_refill_fetch_1_pageFault;
              end
              if(_zz_54) begin
                TrapPlugin_logic_harts_0_trap_fsm_atsPorts_refill_rsp_payload_pageFault = MmuPlugin_logic_refill_fetch_1_pageFault;
              end
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    TrapPlugin_logic_harts_0_trap_fsm_atsPorts_refill_rsp_payload_accessFault = 1'bx;
    case(MmuPlugin_logic_refill_stateReg)
      MmuPlugin_logic_refill_enumDef_IDLE : begin
      end
      MmuPlugin_logic_refill_enumDef_CMD_0 : begin
      end
      MmuPlugin_logic_refill_enumDef_CMD_1 : begin
      end
      MmuPlugin_logic_refill_enumDef_RSP_0 : begin
        if(MmuPlugin_logic_refill_load_rsp_valid) begin
          if(!MmuPlugin_logic_refill_load_rsp_payload_redo) begin
            if(_zz_54) begin
              TrapPlugin_logic_harts_0_trap_fsm_atsPorts_refill_rsp_payload_accessFault = MmuPlugin_logic_refill_fetch_0_accessFault;
            end
            if(_zz_54) begin
              TrapPlugin_logic_harts_0_trap_fsm_atsPorts_refill_rsp_payload_accessFault = MmuPlugin_logic_refill_fetch_0_accessFault;
            end
          end
        end
      end
      MmuPlugin_logic_refill_enumDef_RSP_1 : begin
        if(MmuPlugin_logic_refill_load_rsp_valid) begin
          if(!MmuPlugin_logic_refill_load_rsp_payload_redo) begin
            if(when_MmuPlugin_l471) begin
              if(_zz_54) begin
                TrapPlugin_logic_harts_0_trap_fsm_atsPorts_refill_rsp_payload_accessFault = MmuPlugin_logic_refill_fetch_1_accessFault;
              end
              if(_zz_54) begin
                TrapPlugin_logic_harts_0_trap_fsm_atsPorts_refill_rsp_payload_accessFault = MmuPlugin_logic_refill_fetch_1_accessFault;
              end
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  assign MmuPlugin_logic_refill_fetch_0_pageFault = ((MmuPlugin_logic_refill_load_exception || MmuPlugin_logic_refill_load_levelException_0) || (! MmuPlugin_logic_refill_load_flags_A));
  assign MmuPlugin_logic_refill_fetch_0_accessFault = ((! MmuPlugin_logic_refill_fetch_0_pageFault) && 1'b0);
  assign MmuPlugin_logic_refill_fetch_1_pageFault = ((MmuPlugin_logic_refill_load_exception || MmuPlugin_logic_refill_load_levelException_1) || (! MmuPlugin_logic_refill_load_flags_A));
  assign MmuPlugin_logic_refill_fetch_1_accessFault = ((! MmuPlugin_logic_refill_fetch_1_pageFault) && 1'b0);
  assign TrapPlugin_logic_harts_0_trap_fsm_atsPorts_invalidate_cmd_ready = MmuPlugin_logic_invalidate_arbiter_io_inputs_0_ready;
  always @(*) begin
    MmuPlugin_logic_invalidate_arbiter_io_output_ready = 1'b0;
    if(!when_MmuPlugin_l496) begin
      if(when_MmuPlugin_l510) begin
        MmuPlugin_logic_invalidate_arbiter_io_output_ready = 1'b1;
      end
    end
  end

  assign when_MmuPlugin_l496 = (! MmuPlugin_logic_invalidate_busy);
  assign when_MmuPlugin_l510 = (&MmuPlugin_logic_invalidate_counter);
  assign LsuTileLinkPlugin_logic_bridge_cmdHash = LsuPlugin_logic_bus_cmd_payload_address[9 : 2];
  assign LsuTileLinkPlugin_logic_bridge_pendings_0_hazard = (LsuTileLinkPlugin_logic_bridge_pendings_0_valid && (((LsuTileLinkPlugin_logic_bridge_pendings_0_hash == LsuTileLinkPlugin_logic_bridge_cmdHash) && (|(LsuTileLinkPlugin_logic_bridge_pendings_0_mask & LsuPlugin_logic_bus_cmd_payload_mask))) || (LsuTileLinkPlugin_logic_bridge_pendings_0_io && LsuPlugin_logic_bus_cmd_payload_io)));
  assign LsuTileLinkPlugin_logic_bridge_hazard = (|LsuTileLinkPlugin_logic_bridge_pendings_0_hazard);
  assign LsuTileLinkPlugin_logic_bridge_down_d_fire = (LsuTileLinkPlugin_logic_bridge_down_d_valid && LsuTileLinkPlugin_logic_bridge_down_d_ready);
  assign LsuTileLinkPlugin_logic_bridge_down_a_fire = (LsuTileLinkPlugin_logic_bridge_down_a_valid && LsuTileLinkPlugin_logic_bridge_down_a_ready);
  assign _zz_LsuPlugin_logic_bus_cmd_ready = (! LsuTileLinkPlugin_logic_bridge_hazard);
  assign LsuPlugin_logic_bus_cmd_ready = (LsuTileLinkPlugin_logic_bridge_down_a_ready && _zz_LsuPlugin_logic_bus_cmd_ready);
  assign LsuTileLinkPlugin_logic_bridge_down_a_valid = (LsuPlugin_logic_bus_cmd_valid && _zz_LsuPlugin_logic_bus_cmd_ready);
  assign _zz_LsuTileLinkPlugin_logic_bridge_down_a_payload_opcode = (LsuPlugin_logic_bus_cmd_payload_write ? A_PUT_FULL_DATA : A_GET);
  assign LsuTileLinkPlugin_logic_bridge_down_a_payload_opcode = _zz_LsuTileLinkPlugin_logic_bridge_down_a_payload_opcode;
  assign LsuTileLinkPlugin_logic_bridge_down_a_payload_param = 3'b000;
  assign LsuTileLinkPlugin_logic_bridge_down_a_payload_address = LsuPlugin_logic_bus_cmd_payload_address;
  assign LsuTileLinkPlugin_logic_bridge_down_a_payload_size = LsuPlugin_logic_bus_cmd_payload_size;
  assign LsuTileLinkPlugin_logic_bridge_down_a_payload_mask = LsuPlugin_logic_bus_cmd_payload_mask;
  assign LsuTileLinkPlugin_logic_bridge_down_a_payload_data = LsuPlugin_logic_bus_cmd_payload_data;
  assign LsuTileLinkPlugin_logic_bridge_down_a_payload_corrupt = 1'b0;
  assign LsuTileLinkPlugin_logic_bridge_down_d_ready = 1'b1;
  assign LsuPlugin_logic_bus_rsp_valid = LsuTileLinkPlugin_logic_bridge_down_d_valid;
  assign LsuPlugin_logic_bus_rsp_payload_error = LsuTileLinkPlugin_logic_bridge_down_d_payload_denied;
  assign LsuPlugin_logic_bus_rsp_payload_data = LsuTileLinkPlugin_logic_bridge_down_d_payload_data;
  assign PcPlugin_logic_forcedSpawn = (|{TrapPlugin_logic_harts_0_trap_pcPort_valid,{late1_BranchPlugin_logic_pcPort_valid,{early1_BranchPlugin_logic_pcPort_valid,{late0_BranchPlugin_logic_pcPort_valid,{early0_BranchPlugin_logic_pcPort_valid,BtbPlugin_logic_pcPort_valid}}}}});
  assign PcPlugin_logic_harts_0_self_pc = (PcPlugin_logic_harts_0_self_state + _zz_PcPlugin_logic_harts_0_self_pc);
  assign PcPlugin_logic_harts_0_self_flow_valid = 1'b1;
  assign PcPlugin_logic_harts_0_self_flow_payload_fault = PcPlugin_logic_harts_0_self_fault;
  assign PcPlugin_logic_harts_0_self_flow_payload_pc = PcPlugin_logic_harts_0_self_pc;
  assign PcPlugin_logic_harts_0_aggregator_sortedByPriority_5_laneValid = 1'b1;
  assign PcPlugin_logic_harts_0_aggregator_sortedByPriority_3_laneValid = (&((! early1_BranchPlugin_logic_pcPort_valid) || (early0_BranchPlugin_logic_pcPort_payload_laneAge < early1_BranchPlugin_logic_pcPort_payload_laneAge)));
  assign PcPlugin_logic_harts_0_aggregator_sortedByPriority_1_laneValid = (&((! late1_BranchPlugin_logic_pcPort_valid) || (late0_BranchPlugin_logic_pcPort_payload_laneAge < late1_BranchPlugin_logic_pcPort_payload_laneAge)));
  assign PcPlugin_logic_harts_0_aggregator_sortedByPriority_4_laneValid = (&((! early0_BranchPlugin_logic_pcPort_valid) || (early1_BranchPlugin_logic_pcPort_payload_laneAge < early0_BranchPlugin_logic_pcPort_payload_laneAge)));
  assign PcPlugin_logic_harts_0_aggregator_sortedByPriority_2_laneValid = (&((! late0_BranchPlugin_logic_pcPort_valid) || (late1_BranchPlugin_logic_pcPort_payload_laneAge < late0_BranchPlugin_logic_pcPort_payload_laneAge)));
  assign PcPlugin_logic_harts_0_aggregator_sortedByPriority_0_laneValid = 1'b1;
  assign PcPlugin_logic_harts_0_aggregator_sortedByPriority_6_laneValid = 1'b1;
  assign PcPlugin_logic_harts_0_aggregator_valids_0 = ((TrapPlugin_logic_harts_0_trap_pcPort_valid && 1'b1) && PcPlugin_logic_harts_0_aggregator_sortedByPriority_0_laneValid);
  assign PcPlugin_logic_harts_0_aggregator_valids_1 = ((late0_BranchPlugin_logic_pcPort_valid && 1'b1) && PcPlugin_logic_harts_0_aggregator_sortedByPriority_1_laneValid);
  assign PcPlugin_logic_harts_0_aggregator_valids_2 = ((late1_BranchPlugin_logic_pcPort_valid && 1'b1) && PcPlugin_logic_harts_0_aggregator_sortedByPriority_2_laneValid);
  assign PcPlugin_logic_harts_0_aggregator_valids_3 = ((early0_BranchPlugin_logic_pcPort_valid && 1'b1) && PcPlugin_logic_harts_0_aggregator_sortedByPriority_3_laneValid);
  assign PcPlugin_logic_harts_0_aggregator_valids_4 = ((early1_BranchPlugin_logic_pcPort_valid && 1'b1) && PcPlugin_logic_harts_0_aggregator_sortedByPriority_4_laneValid);
  assign PcPlugin_logic_harts_0_aggregator_valids_5 = ((BtbPlugin_logic_pcPort_valid && 1'b1) && PcPlugin_logic_harts_0_aggregator_sortedByPriority_5_laneValid);
  assign PcPlugin_logic_harts_0_aggregator_valids_6 = ((PcPlugin_logic_harts_0_self_flow_valid && 1'b1) && PcPlugin_logic_harts_0_aggregator_sortedByPriority_6_laneValid);
  assign _zz_PcPlugin_logic_harts_0_aggregator_oh = {PcPlugin_logic_harts_0_aggregator_valids_6,{PcPlugin_logic_harts_0_aggregator_valids_5,{PcPlugin_logic_harts_0_aggregator_valids_4,{PcPlugin_logic_harts_0_aggregator_valids_3,{PcPlugin_logic_harts_0_aggregator_valids_2,{PcPlugin_logic_harts_0_aggregator_valids_1,PcPlugin_logic_harts_0_aggregator_valids_0}}}}}};
  assign _zz_PcPlugin_logic_harts_0_aggregator_oh_1 = _zz_PcPlugin_logic_harts_0_aggregator_oh[0];
  assign _zz_PcPlugin_logic_harts_0_aggregator_oh_2 = _zz_PcPlugin_logic_harts_0_aggregator_oh[1];
  assign _zz_PcPlugin_logic_harts_0_aggregator_oh_3 = _zz_PcPlugin_logic_harts_0_aggregator_oh[2];
  assign _zz_PcPlugin_logic_harts_0_aggregator_oh_4 = _zz_PcPlugin_logic_harts_0_aggregator_oh[3];
  assign _zz_PcPlugin_logic_harts_0_aggregator_oh_5 = _zz_PcPlugin_logic_harts_0_aggregator_oh[4];
  assign _zz_PcPlugin_logic_harts_0_aggregator_oh_6 = _zz_PcPlugin_logic_harts_0_aggregator_oh[5];
  always @(*) begin
    _zz_PcPlugin_logic_harts_0_aggregator_oh_7[0] = (_zz_PcPlugin_logic_harts_0_aggregator_oh_1 && (! 1'b0));
    _zz_PcPlugin_logic_harts_0_aggregator_oh_7[1] = (_zz_PcPlugin_logic_harts_0_aggregator_oh_2 && (! _zz_PcPlugin_logic_harts_0_aggregator_oh_1));
    _zz_PcPlugin_logic_harts_0_aggregator_oh_7[2] = (_zz_PcPlugin_logic_harts_0_aggregator_oh_3 && (! (|{_zz_PcPlugin_logic_harts_0_aggregator_oh_2,_zz_PcPlugin_logic_harts_0_aggregator_oh_1})));
    _zz_PcPlugin_logic_harts_0_aggregator_oh_7[3] = (_zz_PcPlugin_logic_harts_0_aggregator_oh_4 && (! (|{_zz_PcPlugin_logic_harts_0_aggregator_oh_3,{_zz_PcPlugin_logic_harts_0_aggregator_oh_2,_zz_PcPlugin_logic_harts_0_aggregator_oh_1}})));
    _zz_PcPlugin_logic_harts_0_aggregator_oh_7[4] = (_zz_PcPlugin_logic_harts_0_aggregator_oh_5 && (! _zz_PcPlugin_logic_harts_0_aggregator_oh_8));
    _zz_PcPlugin_logic_harts_0_aggregator_oh_7[5] = (_zz_PcPlugin_logic_harts_0_aggregator_oh_6 && (! (_zz_PcPlugin_logic_harts_0_aggregator_oh_5 || _zz_PcPlugin_logic_harts_0_aggregator_oh_8)));
    _zz_PcPlugin_logic_harts_0_aggregator_oh_7[6] = (_zz_PcPlugin_logic_harts_0_aggregator_oh[6] && (! ((|{_zz_PcPlugin_logic_harts_0_aggregator_oh_6,_zz_PcPlugin_logic_harts_0_aggregator_oh_5}) || _zz_PcPlugin_logic_harts_0_aggregator_oh_8)));
  end

  assign _zz_PcPlugin_logic_harts_0_aggregator_oh_8 = (|{_zz_PcPlugin_logic_harts_0_aggregator_oh_4,{_zz_PcPlugin_logic_harts_0_aggregator_oh_3,{_zz_PcPlugin_logic_harts_0_aggregator_oh_2,_zz_PcPlugin_logic_harts_0_aggregator_oh_1}}});
  assign PcPlugin_logic_harts_0_aggregator_oh = _zz_PcPlugin_logic_harts_0_aggregator_oh_7;
  assign _zz_PcPlugin_logic_harts_0_aggregator_target = PcPlugin_logic_harts_0_aggregator_oh[0];
  assign _zz_PcPlugin_logic_harts_0_aggregator_target_1 = PcPlugin_logic_harts_0_aggregator_oh[1];
  assign _zz_PcPlugin_logic_harts_0_aggregator_target_2 = PcPlugin_logic_harts_0_aggregator_oh[2];
  assign _zz_PcPlugin_logic_harts_0_aggregator_target_3 = PcPlugin_logic_harts_0_aggregator_oh[3];
  assign _zz_PcPlugin_logic_harts_0_aggregator_target_4 = PcPlugin_logic_harts_0_aggregator_oh[4];
  assign _zz_PcPlugin_logic_harts_0_aggregator_target_5 = PcPlugin_logic_harts_0_aggregator_oh[5];
  assign _zz_PcPlugin_logic_harts_0_aggregator_target_6 = PcPlugin_logic_harts_0_aggregator_oh[6];
  assign PcPlugin_logic_harts_0_aggregator_target = ((((_zz_PcPlugin_logic_harts_0_aggregator_target ? _zz_PcPlugin_logic_harts_0_aggregator_target_7 : _zz_PcPlugin_logic_harts_0_aggregator_target_8) | (_zz_PcPlugin_logic_harts_0_aggregator_target_1 ? _zz_PcPlugin_logic_harts_0_aggregator_target_9 : _zz_PcPlugin_logic_harts_0_aggregator_target_10)) | ((_zz_PcPlugin_logic_harts_0_aggregator_target_2 ? _zz_PcPlugin_logic_harts_0_aggregator_target_11 : _zz_PcPlugin_logic_harts_0_aggregator_target_12) | (_zz_PcPlugin_logic_harts_0_aggregator_target_3 ? _zz_PcPlugin_logic_harts_0_aggregator_target_13 : _zz_PcPlugin_logic_harts_0_aggregator_target_14))) | (((_zz_PcPlugin_logic_harts_0_aggregator_target_4 ? _zz_PcPlugin_logic_harts_0_aggregator_target_15 : _zz_PcPlugin_logic_harts_0_aggregator_target_16) | (_zz_PcPlugin_logic_harts_0_aggregator_target_5 ? _zz_PcPlugin_logic_harts_0_aggregator_target_17 : _zz_PcPlugin_logic_harts_0_aggregator_target_18)) | (_zz_PcPlugin_logic_harts_0_aggregator_target_6 ? PcPlugin_logic_harts_0_self_flow_payload_pc : 32'h0)));
  assign PcPlugin_logic_harts_0_aggregator_fault = _zz_PcPlugin_logic_harts_0_aggregator_fault[0];
  assign PcPlugin_logic_harts_0_holdComb = (|TrapPlugin_logic_harts_0_trap_fsm_holdPort);
  assign PcPlugin_logic_harts_0_output_valid = (! PcPlugin_logic_harts_0_holdReg);
  assign PcPlugin_logic_harts_0_output_payload_fault = PcPlugin_logic_harts_0_aggregator_fault;
  always @(*) begin
    PcPlugin_logic_harts_0_output_payload_pc = PcPlugin_logic_harts_0_aggregator_target;
    PcPlugin_logic_harts_0_output_payload_pc[0 : 0] = 1'b0;
  end

  assign PcPlugin_logic_harts_0_output_fire = (PcPlugin_logic_harts_0_output_valid && PcPlugin_logic_harts_0_output_ready);
  assign fetch_logic_ctrls_0_up_valid = PcPlugin_logic_harts_0_output_valid;
  assign PcPlugin_logic_harts_0_output_ready = fetch_logic_ctrls_0_up_ready;
  assign fetch_logic_ctrls_0_up_Fetch_WORD_PC = PcPlugin_logic_harts_0_output_payload_pc;
  assign fetch_logic_ctrls_0_up_Fetch_PC_FAULT = PcPlugin_logic_harts_0_output_payload_fault;
  always @(*) begin
    fetch_logic_ctrls_0_up_Fetch_ID = 10'bxxxxxxxxxx;
    fetch_logic_ctrls_0_up_Fetch_ID = PcPlugin_logic_harts_0_self_id;
  end

  assign PcPlugin_logic_holdHalter_doIt = PcPlugin_logic_harts_0_holdComb;
  assign fetch_logic_ctrls_0_haltRequest_PcPlugin_l136 = PcPlugin_logic_holdHalter_doIt;
  assign CsrAccessPlugin_logic_fsm_wantExit = 1'b0;
  always @(*) begin
    CsrAccessPlugin_logic_fsm_wantStart = 1'b0;
    case(CsrAccessPlugin_logic_fsm_stateReg)
      CsrAccessPlugin_logic_fsm_enumDef_READ : begin
      end
      CsrAccessPlugin_logic_fsm_enumDef_WRITE : begin
      end
      CsrAccessPlugin_logic_fsm_enumDef_COMPLETION : begin
      end
      default : begin
        CsrAccessPlugin_logic_fsm_wantStart = 1'b1;
      end
    endcase
  end

  assign CsrAccessPlugin_logic_fsm_wantKill = 1'b0;
  always @(*) begin
    CsrAccessPlugin_logic_fsm_regs_fire = 1'b0;
    case(CsrAccessPlugin_logic_fsm_stateReg)
      CsrAccessPlugin_logic_fsm_enumDef_READ : begin
      end
      CsrAccessPlugin_logic_fsm_enumDef_WRITE : begin
      end
      CsrAccessPlugin_logic_fsm_enumDef_COMPLETION : begin
        if(toplevel_execute_ctrl2_down_isReady) begin
          CsrAccessPlugin_logic_fsm_regs_fire = 1'b1;
        end
      end
      default : begin
      end
    endcase
  end

  assign CsrAccessPlugin_logic_fsm_inject_csrAddress = toplevel_execute_ctrl2_down_Decode_UOP_lane0[31 : 20];
  assign CsrAccessPlugin_logic_fsm_inject_immZero = (toplevel_execute_ctrl2_down_Decode_UOP_lane0[19 : 15] == 5'h0);
  assign CsrAccessPlugin_logic_fsm_inject_srcZero = (toplevel_execute_ctrl2_down_CsrAccessPlugin_CSR_IMM_lane0 ? CsrAccessPlugin_logic_fsm_inject_immZero : (toplevel_execute_ctrl2_down_Decode_UOP_lane0[19 : 15] == 5'h0));
  assign CsrAccessPlugin_logic_fsm_inject_csrWrite = (! (toplevel_execute_ctrl2_down_CsrAccessPlugin_CSR_MASK_lane0 && CsrAccessPlugin_logic_fsm_inject_srcZero));
  assign CsrAccessPlugin_logic_fsm_inject_csrRead = (! ((! toplevel_execute_ctrl2_down_CsrAccessPlugin_CSR_MASK_lane0) && (! toplevel_execute_ctrl2_up_RD_ENABLE_lane0)));
  assign COMB_CSR_1952 = (CsrAccessPlugin_logic_fsm_inject_csrAddress == 12'h7a0);
  assign COMB_CSR_1953 = (CsrAccessPlugin_logic_fsm_inject_csrAddress == 12'h7a1);
  assign COMB_CSR_1954 = (CsrAccessPlugin_logic_fsm_inject_csrAddress == 12'h7a2);
  assign COMB_CSR_3857 = (CsrAccessPlugin_logic_fsm_inject_csrAddress == 12'hf11);
  assign COMB_CSR_3858 = (CsrAccessPlugin_logic_fsm_inject_csrAddress == 12'hf12);
  assign COMB_CSR_3859 = (CsrAccessPlugin_logic_fsm_inject_csrAddress == 12'hf13);
  assign COMB_CSR_3860 = (CsrAccessPlugin_logic_fsm_inject_csrAddress == 12'hf14);
  assign COMB_CSR_769 = (CsrAccessPlugin_logic_fsm_inject_csrAddress == 12'h301);
  assign COMB_CSR_768 = (CsrAccessPlugin_logic_fsm_inject_csrAddress == 12'h300);
  assign COMB_CSR_834 = (CsrAccessPlugin_logic_fsm_inject_csrAddress == 12'h342);
  assign COMB_CSR_836 = (CsrAccessPlugin_logic_fsm_inject_csrAddress == 12'h344);
  assign COMB_CSR_772 = (CsrAccessPlugin_logic_fsm_inject_csrAddress == 12'h304);
  assign COMB_CSR_770 = (CsrAccessPlugin_logic_fsm_inject_csrAddress == 12'h302);
  assign COMB_CSR_771 = (CsrAccessPlugin_logic_fsm_inject_csrAddress == 12'h303);
  assign COMB_CSR_322 = (CsrAccessPlugin_logic_fsm_inject_csrAddress == 12'h142);
  assign COMB_CSR_256 = (CsrAccessPlugin_logic_fsm_inject_csrAddress == 12'h100);
  assign COMB_CSR_260 = (CsrAccessPlugin_logic_fsm_inject_csrAddress == 12'h104);
  assign COMB_CSR_324 = (CsrAccessPlugin_logic_fsm_inject_csrAddress == 12'h144);
  assign COMB_CSR_3073 = (CsrAccessPlugin_logic_fsm_inject_csrAddress == 12'hc01);
  assign COMB_CSR_3201 = (CsrAccessPlugin_logic_fsm_inject_csrAddress == 12'hc81);
  assign COMB_CSR_PrivilegedPlugin_logic_readAnyWriteLegal_tvecFilter = (|{(CsrAccessPlugin_logic_fsm_inject_csrAddress == 12'h105),(CsrAccessPlugin_logic_fsm_inject_csrAddress == 12'h305)});
  assign COMB_CSR_PrivilegedPlugin_logic_readAnyWriteLegal_epcFilter = (|{(CsrAccessPlugin_logic_fsm_inject_csrAddress == 12'h141),(CsrAccessPlugin_logic_fsm_inject_csrAddress == 12'h341)});
  assign COMB_CSR_384 = (CsrAccessPlugin_logic_fsm_inject_csrAddress == 12'h180);
  assign COMB_CSR_CsrRamPlugin_csrMapper_selFilter = (|{(CsrAccessPlugin_logic_fsm_inject_csrAddress == 12'h140),{(CsrAccessPlugin_logic_fsm_inject_csrAddress == 12'h141),{(CsrAccessPlugin_logic_fsm_inject_csrAddress == 12'h143),{(CsrAccessPlugin_logic_fsm_inject_csrAddress == 12'h105),{(CsrAccessPlugin_logic_fsm_inject_csrAddress == _zz_COMB_CSR_CsrRamPlugin_csrMapper_selFilter),{_zz_COMB_CSR_CsrRamPlugin_csrMapper_selFilter_1,{_zz_COMB_CSR_CsrRamPlugin_csrMapper_selFilter_2,_zz_COMB_CSR_CsrRamPlugin_csrMapper_selFilter_3}}}}}}});
  assign COMB_CSR_CsrAccessPlugin_logic_trapNextOnWriteFilter = (|{(CsrAccessPlugin_logic_fsm_inject_csrAddress == 12'h100),(CsrAccessPlugin_logic_fsm_inject_csrAddress == 12'h300)});
  assign CsrAccessPlugin_logic_fsm_inject_implemented = (|{COMB_CSR_CsrAccessPlugin_logic_trapNextOnWriteFilter,{COMB_CSR_CsrRamPlugin_csrMapper_selFilter,{COMB_CSR_384,{COMB_CSR_PrivilegedPlugin_logic_readAnyWriteLegal_epcFilter,{COMB_CSR_PrivilegedPlugin_logic_readAnyWriteLegal_tvecFilter,{COMB_CSR_3201,{COMB_CSR_3073,{COMB_CSR_324,{COMB_CSR_260,{COMB_CSR_256,{_zz_CsrAccessPlugin_logic_fsm_inject_implemented,_zz_CsrAccessPlugin_logic_fsm_inject_implemented_1}}}}}}}}}}});
  assign CsrAccessPlugin_logic_fsm_inject_onDecodeDo = ((toplevel_execute_ctrl2_up_LANE_SEL_lane0 && toplevel_execute_ctrl2_down_CsrAccessPlugin_SEL_lane0) && (CsrAccessPlugin_logic_fsm_stateReg == CsrAccessPlugin_logic_fsm_enumDef_IDLE));
  assign when_CsrAccessPlugin_l155 = (CsrAccessPlugin_logic_fsm_inject_onDecodeDo && COMB_CSR_384);
  assign when_MmuPlugin_l212 = (PrivilegedPlugin_logic_harts_0_m_status_tvm && (PrivilegedPlugin_logic_harts_0_privilege == 2'b01));
  assign when_CsrAccessPlugin_l155_1 = (CsrAccessPlugin_logic_fsm_inject_onDecodeDo && COMB_CSR_CsrAccessPlugin_logic_trapNextOnWriteFilter);
  assign CsrAccessPlugin_logic_fsm_inject_trap = ((! CsrAccessPlugin_logic_fsm_inject_implemented) || CsrAccessPlugin_bus_decode_exception);
  assign CsrAccessPlugin_bus_decode_read = CsrAccessPlugin_logic_fsm_inject_csrRead;
  assign CsrAccessPlugin_bus_decode_write = CsrAccessPlugin_logic_fsm_inject_csrWrite;
  assign CsrAccessPlugin_bus_decode_address = CsrAccessPlugin_logic_fsm_inject_csrAddress;
  assign CsrAccessPlugin_logic_fsm_regs_uopId = toplevel_execute_ctrl2_down_Decode_UOP_ID_lane0;
  assign CsrAccessPlugin_logic_fsm_regs_rs1 = toplevel_execute_ctrl2_up_integer_RS1_lane0;
  assign CsrAccessPlugin_logic_fsm_regs_uop = toplevel_execute_ctrl2_down_Decode_UOP_lane0;
  assign CsrAccessPlugin_logic_fsm_regs_doImm = toplevel_execute_ctrl2_down_CsrAccessPlugin_CSR_IMM_lane0;
  assign CsrAccessPlugin_logic_fsm_regs_doMask = toplevel_execute_ctrl2_down_CsrAccessPlugin_CSR_MASK_lane0;
  assign CsrAccessPlugin_logic_fsm_regs_doClear = toplevel_execute_ctrl2_down_CsrAccessPlugin_CSR_CLEAR_lane0;
  assign CsrAccessPlugin_logic_fsm_regs_rdEnable = toplevel_execute_ctrl2_up_RD_ENABLE_lane0;
  assign CsrAccessPlugin_logic_fsm_regs_rdPhys = toplevel_execute_ctrl2_down_RD_PHYS_lane0;
  assign CsrAccessPlugin_logic_fsm_inject_iLogic_freeze = ((toplevel_execute_ctrl2_up_LANE_SEL_lane0 && toplevel_execute_ctrl2_down_CsrAccessPlugin_SEL_lane0) && (! CsrAccessPlugin_logic_fsm_inject_unfreeze));
  always @(*) begin
    CsrAccessPlugin_logic_flushPort_valid = 1'b0;
    if(CsrAccessPlugin_logic_fsm_inject_flushReg) begin
      CsrAccessPlugin_logic_flushPort_valid = 1'b1;
    end
    case(CsrAccessPlugin_logic_fsm_stateReg)
      CsrAccessPlugin_logic_fsm_enumDef_READ : begin
      end
      CsrAccessPlugin_logic_fsm_enumDef_WRITE : begin
      end
      CsrAccessPlugin_logic_fsm_enumDef_COMPLETION : begin
      end
      default : begin
        if(CsrAccessPlugin_logic_fsm_inject_onDecodeDo) begin
          if(CsrAccessPlugin_logic_fsm_inject_sampled) begin
            if(CsrAccessPlugin_logic_fsm_inject_trapReg) begin
              CsrAccessPlugin_logic_flushPort_valid = 1'b1;
            end else begin
              if(CsrAccessPlugin_logic_fsm_inject_busTrapReg) begin
                CsrAccessPlugin_logic_flushPort_valid = 1'b1;
              end
            end
          end
        end
      end
    endcase
  end

  assign CsrAccessPlugin_logic_flushPort_payload_uopId = toplevel_execute_ctrl2_down_Decode_UOP_ID_lane0;
  assign CsrAccessPlugin_logic_flushPort_payload_laneAge = toplevel_execute_ctrl2_down_LANE_AGE_lane0;
  assign CsrAccessPlugin_logic_flushPort_payload_self = 1'b0;
  always @(*) begin
    CsrAccessPlugin_logic_trapPort_valid = 1'b0;
    case(CsrAccessPlugin_logic_fsm_stateReg)
      CsrAccessPlugin_logic_fsm_enumDef_READ : begin
      end
      CsrAccessPlugin_logic_fsm_enumDef_WRITE : begin
      end
      CsrAccessPlugin_logic_fsm_enumDef_COMPLETION : begin
      end
      default : begin
        if(CsrAccessPlugin_logic_fsm_inject_onDecodeDo) begin
          if(CsrAccessPlugin_logic_fsm_inject_sampled) begin
            if(CsrAccessPlugin_logic_fsm_inject_trapReg) begin
              CsrAccessPlugin_logic_trapPort_valid = 1'b1;
            end else begin
              if(CsrAccessPlugin_logic_fsm_inject_busTrapReg) begin
                CsrAccessPlugin_logic_trapPort_valid = 1'b1;
              end
            end
          end
        end
      end
    endcase
  end

  always @(*) begin
    CsrAccessPlugin_logic_trapPort_payload_exception = 1'b1;
    case(CsrAccessPlugin_logic_fsm_stateReg)
      CsrAccessPlugin_logic_fsm_enumDef_READ : begin
      end
      CsrAccessPlugin_logic_fsm_enumDef_WRITE : begin
      end
      CsrAccessPlugin_logic_fsm_enumDef_COMPLETION : begin
      end
      default : begin
        if(CsrAccessPlugin_logic_fsm_inject_onDecodeDo) begin
          if(CsrAccessPlugin_logic_fsm_inject_sampled) begin
            if(!CsrAccessPlugin_logic_fsm_inject_trapReg) begin
              if(CsrAccessPlugin_logic_fsm_inject_busTrapReg) begin
                CsrAccessPlugin_logic_trapPort_payload_exception = 1'b0;
              end
            end
          end
        end
      end
    endcase
  end

  always @(*) begin
    CsrAccessPlugin_logic_trapPort_payload_code = 4'b0010;
    case(CsrAccessPlugin_logic_fsm_stateReg)
      CsrAccessPlugin_logic_fsm_enumDef_READ : begin
      end
      CsrAccessPlugin_logic_fsm_enumDef_WRITE : begin
      end
      CsrAccessPlugin_logic_fsm_enumDef_COMPLETION : begin
      end
      default : begin
        if(CsrAccessPlugin_logic_fsm_inject_onDecodeDo) begin
          if(CsrAccessPlugin_logic_fsm_inject_sampled) begin
            if(!CsrAccessPlugin_logic_fsm_inject_trapReg) begin
              if(CsrAccessPlugin_logic_fsm_inject_busTrapReg) begin
                CsrAccessPlugin_logic_trapPort_payload_code = CsrAccessPlugin_logic_fsm_inject_busTrapCodeReg;
              end
            end
          end
        end
      end
    endcase
  end

  assign CsrAccessPlugin_logic_trapPort_payload_tval = toplevel_execute_ctrl2_down_Decode_UOP_lane0;
  assign CsrAccessPlugin_logic_trapPort_payload_arg = 3'b000;
  assign CsrAccessPlugin_logic_trapPort_payload_laneAge = toplevel_execute_ctrl2_down_LANE_AGE_lane0;
  assign when_CsrAccessPlugin_l209 = (! execute_freeze_valid);
  always @(*) begin
    CsrAccessPlugin_logic_fsm_readLogic_onReadsDo = 1'b0;
    case(CsrAccessPlugin_logic_fsm_stateReg)
      CsrAccessPlugin_logic_fsm_enumDef_READ : begin
        CsrAccessPlugin_logic_fsm_readLogic_onReadsDo = CsrAccessPlugin_logic_fsm_regs_read;
      end
      CsrAccessPlugin_logic_fsm_enumDef_WRITE : begin
      end
      CsrAccessPlugin_logic_fsm_enumDef_COMPLETION : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    CsrAccessPlugin_logic_fsm_readLogic_onReadsFireDo = 1'b0;
    case(CsrAccessPlugin_logic_fsm_stateReg)
      CsrAccessPlugin_logic_fsm_enumDef_READ : begin
        if(when_CsrAccessPlugin_l308) begin
          CsrAccessPlugin_logic_fsm_readLogic_onReadsFireDo = CsrAccessPlugin_logic_fsm_regs_read;
        end
      end
      CsrAccessPlugin_logic_fsm_enumDef_WRITE : begin
      end
      CsrAccessPlugin_logic_fsm_enumDef_COMPLETION : begin
      end
      default : begin
      end
    endcase
  end

  assign CsrAccessPlugin_bus_read_valid = CsrAccessPlugin_logic_fsm_readLogic_onReadsDo;
  assign CsrAccessPlugin_bus_read_address = CsrAccessPlugin_logic_fsm_regs_uop[31 : 20];
  assign CsrAccessPlugin_bus_read_moving = (! CsrAccessPlugin_bus_read_halt);
  assign when_CsrAccessPlugin_l264 = (CsrAccessPlugin_logic_fsm_readLogic_onReadsDo && REG_CSR_CsrRamPlugin_csrMapper_selFilter);
  assign CsrAccessPlugin_logic_fsm_readLogic_csrValue = (((((_zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_13 | _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_16) | (_zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_17 | _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_20)) | ((_zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_25 | _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_29) | (_zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_34 | _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_38))) | (((_zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_43 | _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_48) | (_zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_53 | _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_58)) | ((_zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_63 | _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_68) | (_zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_73 | _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_78)))) | ((((_zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_82 | _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_86) | (_zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_91 | _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_96)) | ((_zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_101 | _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_106) | (_zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_111 | _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_116))) | (((_zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_121 | _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_126) | (_zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_131 | _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_134)) | ((_zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_137 | _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_142) | (_zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_147 | _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_151)))));
  assign CsrAccessPlugin_bus_read_data = CsrAccessPlugin_logic_fsm_readLogic_csrValue;
  always @(*) begin
    CsrAccessPlugin_bus_read_toWriteBits = CsrAccessPlugin_logic_fsm_readLogic_csrValue;
    if(when_CsrAccessPlugin_l291) begin
      if(when_CsrService_l188) begin
        CsrAccessPlugin_bus_read_toWriteBits[9 : 9] = PrivilegedPlugin_logic_harts_0_s_ip_seipSoft;
      end
    end
  end

  assign when_CsrAccessPlugin_l291 = (CsrAccessPlugin_logic_fsm_readLogic_onReadsDo && REG_CSR_836);
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue = REG_CSR_768;
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_8 = REG_CSR_256;
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_12 = REG_CSR_384;
  assign when_CsrService_l188 = 1'b1;
  assign CsrAccessPlugin_bus_write_moving = (! CsrAccessPlugin_bus_write_halt);
  assign CsrAccessPlugin_logic_fsm_writeLogic_alu_mask = (CsrAccessPlugin_logic_fsm_regs_doImm ? _zz_CsrAccessPlugin_logic_fsm_writeLogic_alu_mask : CsrAccessPlugin_logic_fsm_regs_rs1);
  assign CsrAccessPlugin_logic_fsm_writeLogic_alu_masked = (CsrAccessPlugin_logic_fsm_regs_doClear ? (CsrAccessPlugin_logic_fsm_regs_aluInput & (~ CsrAccessPlugin_logic_fsm_writeLogic_alu_mask)) : (CsrAccessPlugin_logic_fsm_regs_aluInput | CsrAccessPlugin_logic_fsm_writeLogic_alu_mask));
  assign CsrAccessPlugin_logic_fsm_writeLogic_alu_result = (CsrAccessPlugin_logic_fsm_regs_doMask ? CsrAccessPlugin_logic_fsm_writeLogic_alu_masked : CsrAccessPlugin_logic_fsm_writeLogic_alu_mask);
  always @(*) begin
    CsrAccessPlugin_bus_write_bits = CsrAccessPlugin_logic_fsm_writeLogic_alu_result;
    if(when_CsrAccessPlugin_l356) begin
      CsrAccessPlugin_bus_write_bits[1 : 0] = 2'b00;
    end
    if(when_CsrAccessPlugin_l356_1) begin
      CsrAccessPlugin_bus_write_bits[0 : 0] = 1'b0;
    end
  end

  assign CsrAccessPlugin_bus_write_address = CsrAccessPlugin_logic_fsm_regs_uop[31 : 20];
  always @(*) begin
    CsrAccessPlugin_logic_fsm_writeLogic_onWritesDo = 1'b0;
    case(CsrAccessPlugin_logic_fsm_stateReg)
      CsrAccessPlugin_logic_fsm_enumDef_READ : begin
      end
      CsrAccessPlugin_logic_fsm_enumDef_WRITE : begin
        CsrAccessPlugin_logic_fsm_writeLogic_onWritesDo = CsrAccessPlugin_logic_fsm_regs_write;
      end
      CsrAccessPlugin_logic_fsm_enumDef_COMPLETION : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    CsrAccessPlugin_logic_fsm_writeLogic_onWritesFireDo = 1'b0;
    case(CsrAccessPlugin_logic_fsm_stateReg)
      CsrAccessPlugin_logic_fsm_enumDef_READ : begin
      end
      CsrAccessPlugin_logic_fsm_enumDef_WRITE : begin
        if(when_CsrAccessPlugin_l338) begin
          CsrAccessPlugin_logic_fsm_writeLogic_onWritesFireDo = CsrAccessPlugin_logic_fsm_regs_write;
        end
      end
      CsrAccessPlugin_logic_fsm_enumDef_COMPLETION : begin
      end
      default : begin
      end
    endcase
  end

  assign CsrAccessPlugin_bus_write_valid = CsrAccessPlugin_logic_fsm_writeLogic_onWritesDo;
  assign when_CsrService_l166 = 1'b1;
  assign when_CsrAccessPlugin_l359 = (CsrAccessPlugin_logic_fsm_writeLogic_onWritesFireDo && REG_CSR_768);
  assign switch_PrivilegedPlugin_l540 = CsrAccessPlugin_bus_write_bits[12 : 11];
  assign when_CsrAccessPlugin_l359_1 = (CsrAccessPlugin_logic_fsm_writeLogic_onWritesFireDo && REG_CSR_834);
  assign when_CsrAccessPlugin_l359_2 = (CsrAccessPlugin_logic_fsm_writeLogic_onWritesFireDo && REG_CSR_836);
  assign when_CsrAccessPlugin_l359_3 = (CsrAccessPlugin_logic_fsm_writeLogic_onWritesFireDo && REG_CSR_772);
  assign when_CsrAccessPlugin_l359_4 = (CsrAccessPlugin_logic_fsm_writeLogic_onWritesFireDo && REG_CSR_770);
  assign when_CsrAccessPlugin_l359_5 = (CsrAccessPlugin_logic_fsm_writeLogic_onWritesFireDo && REG_CSR_771);
  assign when_CsrAccessPlugin_l359_6 = (CsrAccessPlugin_logic_fsm_writeLogic_onWritesFireDo && REG_CSR_322);
  assign when_CsrAccessPlugin_l359_7 = (CsrAccessPlugin_logic_fsm_writeLogic_onWritesFireDo && REG_CSR_256);
  assign when_CsrAccessPlugin_l359_8 = (CsrAccessPlugin_logic_fsm_writeLogic_onWritesFireDo && REG_CSR_260);
  assign when_CsrAccessPlugin_l359_9 = (CsrAccessPlugin_logic_fsm_writeLogic_onWritesFireDo && REG_CSR_324);
  assign when_CsrAccessPlugin_l356 = (CsrAccessPlugin_logic_fsm_writeLogic_onWritesDo && REG_CSR_PrivilegedPlugin_logic_readAnyWriteLegal_tvecFilter);
  assign when_CsrAccessPlugin_l356_1 = (CsrAccessPlugin_logic_fsm_writeLogic_onWritesDo && REG_CSR_PrivilegedPlugin_logic_readAnyWriteLegal_epcFilter);
  assign when_CsrAccessPlugin_l366 = ((|((MmuPlugin_logic_satpModeWrite != 1'b0) && (MmuPlugin_logic_satpModeWrite != 1'b1))) == 1'b0);
  assign when_CsrAccessPlugin_l359_10 = (CsrAccessPlugin_logic_fsm_writeLogic_onWritesFireDo && REG_CSR_384);
  assign when_CsrAccessPlugin_l356_2 = (CsrAccessPlugin_logic_fsm_writeLogic_onWritesDo && REG_CSR_CsrRamPlugin_csrMapper_selFilter);
  always @(*) begin
    CsrAccessPlugin_logic_fsm_completion_valid = 1'b0;
    case(CsrAccessPlugin_logic_fsm_stateReg)
      CsrAccessPlugin_logic_fsm_enumDef_READ : begin
      end
      CsrAccessPlugin_logic_fsm_enumDef_WRITE : begin
      end
      CsrAccessPlugin_logic_fsm_enumDef_COMPLETION : begin
        if(toplevel_execute_ctrl2_down_isReady) begin
          CsrAccessPlugin_logic_fsm_completion_valid = 1'b1;
        end
      end
      default : begin
      end
    endcase
  end

  assign CsrAccessPlugin_logic_fsm_completion_payload_uopId = CsrAccessPlugin_logic_fsm_regs_uopId;
  assign CsrAccessPlugin_logic_fsm_completion_payload_trap = toplevel_execute_ctrl2_down_TRAP_lane0;
  assign CsrAccessPlugin_logic_fsm_completion_payload_commit = toplevel_execute_ctrl2_down_COMMIT_lane0;
  assign CsrAccessPlugin_logic_wbWi_valid = toplevel_execute_ctrl3_down_CsrAccessPlugin_SEL_lane0;
  assign CsrAccessPlugin_logic_wbWi_payload = CsrAccessPlugin_logic_fsm_regs_csrValue;
  always @(*) begin
    HistoryPlugin_logic_onFetch_valueNext = HistoryPlugin_logic_onFetch_value;
    if(HistoryPlugin_logic_onFetch_ports_0_valid) begin
      HistoryPlugin_logic_onFetch_valueNext = HistoryPlugin_logic_onFetch_ports_0_payload_history;
    end
    if(HistoryPlugin_logic_onFetch_ports_1_valid) begin
      HistoryPlugin_logic_onFetch_valueNext = HistoryPlugin_logic_onFetch_ports_1_payload_history;
    end
    if(HistoryPlugin_logic_onFetch_ports_2_valid) begin
      HistoryPlugin_logic_onFetch_valueNext = HistoryPlugin_logic_onFetch_ports_2_payload_history;
    end
    if(HistoryPlugin_logic_onFetch_ports_3_valid) begin
      HistoryPlugin_logic_onFetch_valueNext = HistoryPlugin_logic_onFetch_ports_3_payload_history;
    end
  end

  assign HistoryPlugin_logic_onFetch_ports_0_valid = (|BtbPlugin_logic_historyPort_valid);
  assign HistoryPlugin_logic_onFetch_ports_0_payload_history = BtbPlugin_logic_historyPort_payload_history;
  assign HistoryPlugin_logic_onFetch_ports_1_valid = (|{early1_BranchPlugin_logic_historyPort_valid,early0_BranchPlugin_logic_historyPort_valid});
  assign _zz_HistoryPlugin_logic_onFetch_ports_1_payload_history = (((early0_BranchPlugin_logic_historyPort_valid && (&(! (early1_BranchPlugin_logic_historyPort_valid && (early1_BranchPlugin_logic_historyPort_payload_age < early0_BranchPlugin_logic_historyPort_payload_age))))) ? {early0_BranchPlugin_logic_historyPort_payload_age,early0_BranchPlugin_logic_historyPort_payload_history} : 13'h0) | ((early1_BranchPlugin_logic_historyPort_valid && (&(! (early0_BranchPlugin_logic_historyPort_valid && (early0_BranchPlugin_logic_historyPort_payload_age < early1_BranchPlugin_logic_historyPort_payload_age))))) ? {early1_BranchPlugin_logic_historyPort_payload_age,early1_BranchPlugin_logic_historyPort_payload_history} : 13'h0));
  assign HistoryPlugin_logic_onFetch_ports_1_payload_history = _zz_HistoryPlugin_logic_onFetch_ports_1_payload_history[11 : 0];
  assign HistoryPlugin_logic_onFetch_ports_1_payload_age = _zz_HistoryPlugin_logic_onFetch_ports_1_payload_history[12 : 12];
  assign HistoryPlugin_logic_onFetch_ports_2_valid = (|{late1_BranchPlugin_logic_historyPort_valid,late0_BranchPlugin_logic_historyPort_valid});
  assign _zz_HistoryPlugin_logic_onFetch_ports_2_payload_history = (((late0_BranchPlugin_logic_historyPort_valid && (&(! (late1_BranchPlugin_logic_historyPort_valid && (late1_BranchPlugin_logic_historyPort_payload_age < late0_BranchPlugin_logic_historyPort_payload_age))))) ? {late0_BranchPlugin_logic_historyPort_payload_age,late0_BranchPlugin_logic_historyPort_payload_history} : 13'h0) | ((late1_BranchPlugin_logic_historyPort_valid && (&(! (late0_BranchPlugin_logic_historyPort_valid && (late0_BranchPlugin_logic_historyPort_payload_age < late1_BranchPlugin_logic_historyPort_payload_age))))) ? {late1_BranchPlugin_logic_historyPort_payload_age,late1_BranchPlugin_logic_historyPort_payload_history} : 13'h0));
  assign HistoryPlugin_logic_onFetch_ports_2_payload_history = _zz_HistoryPlugin_logic_onFetch_ports_2_payload_history[11 : 0];
  assign HistoryPlugin_logic_onFetch_ports_2_payload_age = _zz_HistoryPlugin_logic_onFetch_ports_2_payload_history[12 : 12];
  assign HistoryPlugin_logic_onFetch_ports_3_valid = (|TrapPlugin_logic_harts_0_trap_historyPort_valid);
  assign HistoryPlugin_logic_onFetch_ports_3_payload_history = TrapPlugin_logic_harts_0_trap_historyPort_payload_history;
  assign fetch_logic_ctrls_0_down_Prediction_BRANCH_HISTORY = HistoryPlugin_logic_onFetch_valueNext;
  assign CsrRamPlugin_logic_writeLogic_hits = {CsrRamPlugin_setup_initPort_valid,{CsrRamPlugin_csrMapper_write_valid,TrapPlugin_logic_harts_0_crsPorts_write_valid}};
  assign CsrRamPlugin_logic_writeLogic_hit = (|CsrRamPlugin_logic_writeLogic_hits);
  assign CsrRamPlugin_logic_writeLogic_hits_ohFirst_input = CsrRamPlugin_logic_writeLogic_hits;
  assign CsrRamPlugin_logic_writeLogic_hits_ohFirst_masked = (CsrRamPlugin_logic_writeLogic_hits_ohFirst_input & (~ _zz_CsrRamPlugin_logic_writeLogic_hits_ohFirst_masked));
  assign CsrRamPlugin_logic_writeLogic_oh = CsrRamPlugin_logic_writeLogic_hits_ohFirst_masked;
  assign _zz_TrapPlugin_logic_harts_0_crsPorts_write_ready = CsrRamPlugin_logic_writeLogic_oh[0];
  assign _zz_CsrRamPlugin_csrMapper_write_ready = CsrRamPlugin_logic_writeLogic_oh[1];
  assign _zz_CsrRamPlugin_setup_initPort_ready = CsrRamPlugin_logic_writeLogic_oh[2];
  assign CsrRamPlugin_logic_writeLogic_port_valid = CsrRamPlugin_logic_writeLogic_hit;
  assign CsrRamPlugin_logic_writeLogic_port_payload_address = (((_zz_TrapPlugin_logic_harts_0_crsPorts_write_ready ? TrapPlugin_logic_harts_0_crsPorts_write_address : 3'b000) | (_zz_CsrRamPlugin_csrMapper_write_ready ? CsrRamPlugin_csrMapper_write_address : 3'b000)) | (_zz_CsrRamPlugin_setup_initPort_ready ? CsrRamPlugin_setup_initPort_address : 3'b000));
  assign CsrRamPlugin_logic_writeLogic_port_payload_data = (((_zz_TrapPlugin_logic_harts_0_crsPorts_write_ready ? TrapPlugin_logic_harts_0_crsPorts_write_data : 32'h0) | (_zz_CsrRamPlugin_csrMapper_write_ready ? CsrRamPlugin_csrMapper_write_data : 32'h0)) | (_zz_CsrRamPlugin_setup_initPort_ready ? CsrRamPlugin_setup_initPort_data : 32'h0));
  assign TrapPlugin_logic_harts_0_crsPorts_write_ready = _zz_TrapPlugin_logic_harts_0_crsPorts_write_ready;
  assign CsrRamPlugin_csrMapper_write_ready = _zz_CsrRamPlugin_csrMapper_write_ready;
  assign CsrRamPlugin_setup_initPort_ready = _zz_CsrRamPlugin_setup_initPort_ready;
  assign CsrRamPlugin_logic_readLogic_hits = {CsrRamPlugin_csrMapper_read_valid,TrapPlugin_logic_harts_0_crsPorts_read_valid};
  assign CsrRamPlugin_logic_readLogic_hit = (|CsrRamPlugin_logic_readLogic_hits);
  assign CsrRamPlugin_logic_readLogic_hits_ohFirst_input = CsrRamPlugin_logic_readLogic_hits;
  assign CsrRamPlugin_logic_readLogic_hits_ohFirst_masked = (CsrRamPlugin_logic_readLogic_hits_ohFirst_input & (~ _zz_CsrRamPlugin_logic_readLogic_hits_ohFirst_masked));
  assign CsrRamPlugin_logic_readLogic_oh = CsrRamPlugin_logic_readLogic_hits_ohFirst_masked;
  assign _zz_CsrRamPlugin_logic_readLogic_sel = CsrRamPlugin_logic_readLogic_oh[1];
  assign CsrRamPlugin_logic_readLogic_sel = _zz_CsrRamPlugin_logic_readLogic_sel;
  assign CsrRamPlugin_logic_readLogic_port_rsp = CsrRamPlugin_logic_mem_spinal_port1;
  assign CsrRamPlugin_logic_readLogic_port_cmd_valid = (((|CsrRamPlugin_logic_readLogic_oh) && (! CsrRamPlugin_logic_writeLogic_port_valid)) && (! CsrRamPlugin_logic_readLogic_busy));
  assign CsrRamPlugin_logic_readLogic_port_cmd_payload = _zz_CsrRamPlugin_logic_readLogic_port_cmd_payload;
  assign TrapPlugin_logic_harts_0_crsPorts_read_ready = CsrRamPlugin_logic_readLogic_ohReg[0];
  assign CsrRamPlugin_csrMapper_read_ready = CsrRamPlugin_logic_readLogic_ohReg[1];
  assign TrapPlugin_logic_harts_0_crsPorts_read_data = CsrRamPlugin_logic_readLogic_port_rsp;
  assign CsrRamPlugin_csrMapper_read_data = CsrRamPlugin_logic_readLogic_port_rsp;
  assign CsrRamPlugin_logic_flush_done = CsrRamPlugin_logic_flush_counter[3];
  assign CsrRamPlugin_setup_initPort_valid = (! CsrRamPlugin_logic_flush_done);
  assign CsrRamPlugin_setup_initPort_address = CsrRamPlugin_logic_flush_counter[2:0];
  assign CsrRamPlugin_setup_initPort_data = 32'h0;
  assign toplevel_execute_lane0_bypasser_integer_RS1_port_valid = (! execute_freeze_valid);
  assign toplevel_execute_lane0_bypasser_integer_RS1_port_address = toplevel_execute_ctrl0_down_RS1_PHYS_lane0;
  always @(*) begin
    toplevel_execute_lane0_bypasser_integer_RS1_bypassEnables[0] = (((toplevel_execute_ctrl2_up_LANE_SEL_lane0 && toplevel_execute_ctrl2_up_RD_ENABLE_lane0) && (toplevel_execute_ctrl2_down_RD_PHYS_lane0 == toplevel_execute_ctrl1_down_RS1_PHYS_lane0)) && 1'b1);
    toplevel_execute_lane0_bypasser_integer_RS1_bypassEnables[1] = (((toplevel_execute_ctrl2_up_LANE_SEL_lane1 && toplevel_execute_ctrl2_up_RD_ENABLE_lane1) && (toplevel_execute_ctrl2_down_RD_PHYS_lane1 == toplevel_execute_ctrl1_down_RS1_PHYS_lane0)) && 1'b1);
    toplevel_execute_lane0_bypasser_integer_RS1_bypassEnables[2] = (((toplevel_execute_ctrl3_up_LANE_SEL_lane0 && toplevel_execute_ctrl3_up_RD_ENABLE_lane0) && (toplevel_execute_ctrl3_down_RD_PHYS_lane0 == toplevel_execute_ctrl1_down_RS1_PHYS_lane0)) && 1'b1);
    toplevel_execute_lane0_bypasser_integer_RS1_bypassEnables[3] = (((toplevel_execute_ctrl3_up_LANE_SEL_lane1 && toplevel_execute_ctrl3_up_RD_ENABLE_lane1) && (toplevel_execute_ctrl3_down_RD_PHYS_lane1 == toplevel_execute_ctrl1_down_RS1_PHYS_lane0)) && 1'b1);
    toplevel_execute_lane0_bypasser_integer_RS1_bypassEnables[4] = (((toplevel_execute_ctrl4_up_LANE_SEL_lane0 && toplevel_execute_ctrl4_up_RD_ENABLE_lane0) && (toplevel_execute_ctrl4_down_RD_PHYS_lane0 == toplevel_execute_ctrl1_down_RS1_PHYS_lane0)) && 1'b1);
    toplevel_execute_lane0_bypasser_integer_RS1_bypassEnables[5] = (((toplevel_execute_ctrl4_up_LANE_SEL_lane1 && toplevel_execute_ctrl4_up_RD_ENABLE_lane1) && (toplevel_execute_ctrl4_down_RD_PHYS_lane1 == toplevel_execute_ctrl1_down_RS1_PHYS_lane0)) && 1'b1);
    toplevel_execute_lane0_bypasser_integer_RS1_bypassEnables[6] = (((toplevel_execute_ctrl5_up_LANE_SEL_lane0 && toplevel_execute_ctrl5_up_RD_ENABLE_lane0) && (toplevel_execute_ctrl5_down_RD_PHYS_lane0 == toplevel_execute_ctrl1_down_RS1_PHYS_lane0)) && 1'b1);
    toplevel_execute_lane0_bypasser_integer_RS1_bypassEnables[7] = (((toplevel_execute_ctrl5_up_LANE_SEL_lane1 && toplevel_execute_ctrl5_up_RD_ENABLE_lane1) && (toplevel_execute_ctrl5_down_RD_PHYS_lane1 == toplevel_execute_ctrl1_down_RS1_PHYS_lane0)) && 1'b1);
    toplevel_execute_lane0_bypasser_integer_RS1_bypassEnables[8] = 1'b1;
  end

  assign _zz_toplevel_execute_lane0_bypasser_integer_RS1_bypassEnables_bools_0 = toplevel_execute_lane0_bypasser_integer_RS1_bypassEnables;
  assign toplevel_execute_lane0_bypasser_integer_RS1_bypassEnables_bools_0 = _zz_toplevel_execute_lane0_bypasser_integer_RS1_bypassEnables_bools_0[0];
  assign toplevel_execute_lane0_bypasser_integer_RS1_bypassEnables_bools_1 = _zz_toplevel_execute_lane0_bypasser_integer_RS1_bypassEnables_bools_0[1];
  assign toplevel_execute_lane0_bypasser_integer_RS1_bypassEnables_bools_2 = _zz_toplevel_execute_lane0_bypasser_integer_RS1_bypassEnables_bools_0[2];
  assign toplevel_execute_lane0_bypasser_integer_RS1_bypassEnables_bools_3 = _zz_toplevel_execute_lane0_bypasser_integer_RS1_bypassEnables_bools_0[3];
  assign toplevel_execute_lane0_bypasser_integer_RS1_bypassEnables_bools_4 = _zz_toplevel_execute_lane0_bypasser_integer_RS1_bypassEnables_bools_0[4];
  assign toplevel_execute_lane0_bypasser_integer_RS1_bypassEnables_bools_5 = _zz_toplevel_execute_lane0_bypasser_integer_RS1_bypassEnables_bools_0[5];
  assign toplevel_execute_lane0_bypasser_integer_RS1_bypassEnables_bools_6 = _zz_toplevel_execute_lane0_bypasser_integer_RS1_bypassEnables_bools_0[6];
  assign toplevel_execute_lane0_bypasser_integer_RS1_bypassEnables_bools_7 = _zz_toplevel_execute_lane0_bypasser_integer_RS1_bypassEnables_bools_0[7];
  assign toplevel_execute_lane0_bypasser_integer_RS1_bypassEnables_bools_8 = _zz_toplevel_execute_lane0_bypasser_integer_RS1_bypassEnables_bools_0[8];
  always @(*) begin
    _zz_toplevel_execute_lane0_bypasser_integer_RS1_sel[0] = (toplevel_execute_lane0_bypasser_integer_RS1_bypassEnables_bools_0 && (! 1'b0));
    _zz_toplevel_execute_lane0_bypasser_integer_RS1_sel[1] = (toplevel_execute_lane0_bypasser_integer_RS1_bypassEnables_bools_1 && (! toplevel_execute_lane0_bypasser_integer_RS1_bypassEnables_bools_0));
    _zz_toplevel_execute_lane0_bypasser_integer_RS1_sel[2] = (toplevel_execute_lane0_bypasser_integer_RS1_bypassEnables_bools_2 && (! toplevel_execute_lane0_bypasser_integer_RS1_bypassEnables_range_0_to_1));
    _zz_toplevel_execute_lane0_bypasser_integer_RS1_sel[3] = (toplevel_execute_lane0_bypasser_integer_RS1_bypassEnables_bools_3 && (! toplevel_execute_lane0_bypasser_integer_RS1_bypassEnables_range_0_to_2));
    _zz_toplevel_execute_lane0_bypasser_integer_RS1_sel[4] = (toplevel_execute_lane0_bypasser_integer_RS1_bypassEnables_bools_4 && (! toplevel_execute_lane0_bypasser_integer_RS1_bypassEnables_range_0_to_3));
    _zz_toplevel_execute_lane0_bypasser_integer_RS1_sel[5] = (toplevel_execute_lane0_bypasser_integer_RS1_bypassEnables_bools_5 && (! (toplevel_execute_lane0_bypasser_integer_RS1_bypassEnables_bools_4 || toplevel_execute_lane0_bypasser_integer_RS1_bypassEnables_range_0_to_3)));
    _zz_toplevel_execute_lane0_bypasser_integer_RS1_sel[6] = (toplevel_execute_lane0_bypasser_integer_RS1_bypassEnables_bools_6 && (! (toplevel_execute_lane0_bypasser_integer_RS1_bypassEnables_range_4_to_5 || toplevel_execute_lane0_bypasser_integer_RS1_bypassEnables_range_0_to_3)));
    _zz_toplevel_execute_lane0_bypasser_integer_RS1_sel[7] = (toplevel_execute_lane0_bypasser_integer_RS1_bypassEnables_bools_7 && (! (toplevel_execute_lane0_bypasser_integer_RS1_bypassEnables_range_4_to_6 || toplevel_execute_lane0_bypasser_integer_RS1_bypassEnables_range_0_to_3)));
    _zz_toplevel_execute_lane0_bypasser_integer_RS1_sel[8] = (toplevel_execute_lane0_bypasser_integer_RS1_bypassEnables_bools_8 && (! (toplevel_execute_lane0_bypasser_integer_RS1_bypassEnables_range_4_to_7 || toplevel_execute_lane0_bypasser_integer_RS1_bypassEnables_range_0_to_3)));
  end

  assign toplevel_execute_lane0_bypasser_integer_RS1_bypassEnables_range_0_to_1 = (|{toplevel_execute_lane0_bypasser_integer_RS1_bypassEnables_bools_1,toplevel_execute_lane0_bypasser_integer_RS1_bypassEnables_bools_0});
  assign toplevel_execute_lane0_bypasser_integer_RS1_bypassEnables_range_0_to_2 = (|{toplevel_execute_lane0_bypasser_integer_RS1_bypassEnables_bools_2,{toplevel_execute_lane0_bypasser_integer_RS1_bypassEnables_bools_1,toplevel_execute_lane0_bypasser_integer_RS1_bypassEnables_bools_0}});
  assign toplevel_execute_lane0_bypasser_integer_RS1_bypassEnables_range_0_to_3 = (|{toplevel_execute_lane0_bypasser_integer_RS1_bypassEnables_bools_3,{toplevel_execute_lane0_bypasser_integer_RS1_bypassEnables_bools_2,{toplevel_execute_lane0_bypasser_integer_RS1_bypassEnables_bools_1,toplevel_execute_lane0_bypasser_integer_RS1_bypassEnables_bools_0}}});
  assign toplevel_execute_lane0_bypasser_integer_RS1_bypassEnables_range_4_to_5 = (|{toplevel_execute_lane0_bypasser_integer_RS1_bypassEnables_bools_5,toplevel_execute_lane0_bypasser_integer_RS1_bypassEnables_bools_4});
  assign toplevel_execute_lane0_bypasser_integer_RS1_bypassEnables_range_4_to_6 = (|{toplevel_execute_lane0_bypasser_integer_RS1_bypassEnables_bools_6,{toplevel_execute_lane0_bypasser_integer_RS1_bypassEnables_bools_5,toplevel_execute_lane0_bypasser_integer_RS1_bypassEnables_bools_4}});
  assign toplevel_execute_lane0_bypasser_integer_RS1_bypassEnables_range_4_to_7 = (|{toplevel_execute_lane0_bypasser_integer_RS1_bypassEnables_bools_7,{toplevel_execute_lane0_bypasser_integer_RS1_bypassEnables_bools_6,{toplevel_execute_lane0_bypasser_integer_RS1_bypassEnables_bools_5,toplevel_execute_lane0_bypasser_integer_RS1_bypassEnables_bools_4}}});
  assign toplevel_execute_lane0_bypasser_integer_RS1_sel = _zz_toplevel_execute_lane0_bypasser_integer_RS1_sel;
  assign _zz_toplevel_execute_ctrl1_down_integer_RS1_lane0 = toplevel_execute_lane0_bypasser_integer_RS1_sel[8 : 1];
  always @(*) begin
    _zz_toplevel_execute_ctrl1_down_integer_RS1_lane0_1 = ((((_zz__zz_toplevel_execute_ctrl1_down_integer_RS1_lane0_1 ? toplevel_execute_ctrl2_down_lane1_integer_WriteBackPlugin_logic_DATA_lane1 : _zz__zz_toplevel_execute_ctrl1_down_integer_RS1_lane0_1_1) | (_zz__zz_toplevel_execute_ctrl1_down_integer_RS1_lane0_1_2 ? toplevel_execute_ctrl3_down_lane0_integer_WriteBackPlugin_logic_DATA_lane0 : _zz__zz_toplevel_execute_ctrl1_down_integer_RS1_lane0_1_3)) | ((_zz__zz_toplevel_execute_ctrl1_down_integer_RS1_lane0_1_4 ? toplevel_execute_ctrl3_down_lane1_integer_WriteBackPlugin_logic_DATA_lane1 : _zz__zz_toplevel_execute_ctrl1_down_integer_RS1_lane0_1_5) | (_zz__zz_toplevel_execute_ctrl1_down_integer_RS1_lane0_1_6 ? toplevel_execute_ctrl4_down_lane0_integer_WriteBackPlugin_logic_DATA_lane0 : _zz__zz_toplevel_execute_ctrl1_down_integer_RS1_lane0_1_7))) | (((_zz__zz_toplevel_execute_ctrl1_down_integer_RS1_lane0_1_8 ? toplevel_execute_ctrl4_down_lane1_integer_WriteBackPlugin_logic_DATA_lane1 : _zz__zz_toplevel_execute_ctrl1_down_integer_RS1_lane0_1_9) | (_zz__zz_toplevel_execute_ctrl1_down_integer_RS1_lane0_1_10 ? toplevel_execute_ctrl5_down_lane0_integer_WriteBackPlugin_logic_DATA_lane0 : _zz__zz_toplevel_execute_ctrl1_down_integer_RS1_lane0_1_11)) | ((_zz__zz_toplevel_execute_ctrl1_down_integer_RS1_lane0_1_12 ? toplevel_execute_ctrl5_down_lane1_integer_WriteBackPlugin_logic_DATA_lane1 : _zz__zz_toplevel_execute_ctrl1_down_integer_RS1_lane0_1_13) | (_zz__zz_toplevel_execute_ctrl1_down_integer_RS1_lane0_1_14 ? toplevel_execute_lane0_bypasser_integer_RS1_port_data : _zz__zz_toplevel_execute_ctrl1_down_integer_RS1_lane0_1_15))));
    if(when_ExecuteLanePlugin_l190) begin
      _zz_toplevel_execute_ctrl1_down_integer_RS1_lane0_1 = toplevel_execute_ctrl2_down_lane0_integer_WriteBackPlugin_logic_DATA_lane0;
    end
  end

  assign toplevel_execute_ctrl1_down_integer_RS1_lane0 = _zz_toplevel_execute_ctrl1_down_integer_RS1_lane0_1;
  assign when_ExecuteLanePlugin_l190 = toplevel_execute_lane0_bypasser_integer_RS1_sel[0];
  assign toplevel_execute_lane0_bypasser_integer_RS1_along_bypasses_0_checks_0_selfHit = (((toplevel_execute_ctrl3_up_LANE_SEL_lane0 && toplevel_execute_ctrl3_up_RD_ENABLE_lane0) && (toplevel_execute_ctrl3_down_RD_PHYS_lane0 == toplevel_execute_ctrl2_down_RS1_PHYS_lane0)) && 1'b1);
  assign toplevel_execute_lane0_bypasser_integer_RS1_along_bypasses_0_checks_0_hit = (toplevel_execute_lane0_bypasser_integer_RS1_along_bypasses_0_checks_0_selfHit && (! 1'b0));
  assign toplevel_execute_lane0_bypasser_integer_RS1_along_bypasses_0_checks_1_selfHit = (((toplevel_execute_ctrl4_up_LANE_SEL_lane0 && toplevel_execute_ctrl4_up_RD_ENABLE_lane0) && (toplevel_execute_ctrl4_down_RD_PHYS_lane0 == toplevel_execute_ctrl2_down_RS1_PHYS_lane0)) && 1'b1);
  assign toplevel_execute_lane0_bypasser_integer_RS1_along_bypasses_0_checks_1_youngerHits_0 = (((toplevel_execute_ctrl3_up_LANE_SEL_lane0 && toplevel_execute_ctrl3_up_RD_ENABLE_lane0) && (toplevel_execute_ctrl3_down_RD_PHYS_lane0 == toplevel_execute_ctrl2_down_RS1_PHYS_lane0)) && 1'b1);
  assign toplevel_execute_lane0_bypasser_integer_RS1_along_bypasses_0_checks_1_youngerHits_1 = (((toplevel_execute_ctrl3_up_LANE_SEL_lane1 && toplevel_execute_ctrl3_up_RD_ENABLE_lane1) && (toplevel_execute_ctrl3_down_RD_PHYS_lane1 == toplevel_execute_ctrl2_down_RS1_PHYS_lane0)) && 1'b1);
  assign toplevel_execute_lane0_bypasser_integer_RS1_along_bypasses_0_checks_1_hit = (toplevel_execute_lane0_bypasser_integer_RS1_along_bypasses_0_checks_1_selfHit && (! (|{toplevel_execute_lane0_bypasser_integer_RS1_along_bypasses_0_checks_1_youngerHits_1,toplevel_execute_lane0_bypasser_integer_RS1_along_bypasses_0_checks_1_youngerHits_0})));
  assign toplevel_execute_lane0_bypasser_integer_RS1_along_bypasses_0_checks_2_selfHit = (((toplevel_execute_ctrl3_up_LANE_SEL_lane1 && toplevel_execute_ctrl3_up_RD_ENABLE_lane1) && (toplevel_execute_ctrl3_down_RD_PHYS_lane1 == toplevel_execute_ctrl2_down_RS1_PHYS_lane0)) && 1'b1);
  assign toplevel_execute_lane0_bypasser_integer_RS1_along_bypasses_0_checks_2_hit = (toplevel_execute_lane0_bypasser_integer_RS1_along_bypasses_0_checks_2_selfHit && (! 1'b0));
  assign toplevel_execute_lane0_bypasser_integer_RS1_along_bypasses_0_checks_3_selfHit = (((toplevel_execute_ctrl4_up_LANE_SEL_lane1 && toplevel_execute_ctrl4_up_RD_ENABLE_lane1) && (toplevel_execute_ctrl4_down_RD_PHYS_lane1 == toplevel_execute_ctrl2_down_RS1_PHYS_lane0)) && 1'b1);
  assign toplevel_execute_lane0_bypasser_integer_RS1_along_bypasses_0_checks_3_youngerHits_0 = (((toplevel_execute_ctrl3_up_LANE_SEL_lane0 && toplevel_execute_ctrl3_up_RD_ENABLE_lane0) && (toplevel_execute_ctrl3_down_RD_PHYS_lane0 == toplevel_execute_ctrl2_down_RS1_PHYS_lane0)) && 1'b1);
  assign toplevel_execute_lane0_bypasser_integer_RS1_along_bypasses_0_checks_3_youngerHits_1 = (((toplevel_execute_ctrl3_up_LANE_SEL_lane1 && toplevel_execute_ctrl3_up_RD_ENABLE_lane1) && (toplevel_execute_ctrl3_down_RD_PHYS_lane1 == toplevel_execute_ctrl2_down_RS1_PHYS_lane0)) && 1'b1);
  assign toplevel_execute_lane0_bypasser_integer_RS1_along_bypasses_0_checks_3_hit = (toplevel_execute_lane0_bypasser_integer_RS1_along_bypasses_0_checks_3_selfHit && (! (|{toplevel_execute_lane0_bypasser_integer_RS1_along_bypasses_0_checks_3_youngerHits_1,toplevel_execute_lane0_bypasser_integer_RS1_along_bypasses_0_checks_3_youngerHits_0})));
  assign toplevel_execute_lane0_bypasser_integer_RS1_along_bypasses_0_hits = {toplevel_execute_lane0_bypasser_integer_RS1_along_bypasses_0_checks_3_hit,{toplevel_execute_lane0_bypasser_integer_RS1_along_bypasses_0_checks_2_hit,{toplevel_execute_lane0_bypasser_integer_RS1_along_bypasses_0_checks_1_hit,toplevel_execute_lane0_bypasser_integer_RS1_along_bypasses_0_checks_0_hit}}};
  assign _zz_toplevel_execute_ctrl2_integer_RS1_lane0_bypass = {toplevel_execute_lane0_bypasser_integer_RS1_along_bypasses_0_hits,(! (|toplevel_execute_lane0_bypasser_integer_RS1_along_bypasses_0_hits))};
  assign toplevel_execute_ctrl2_integer_RS1_lane0_bypass = ((((_zz_toplevel_execute_ctrl2_integer_RS1_lane0_bypass[0] ? toplevel_execute_ctrl2_up_integer_RS1_lane0 : 32'h0) | (_zz_toplevel_execute_ctrl2_integer_RS1_lane0_bypass[1] ? toplevel_execute_ctrl3_down_lane0_integer_WriteBackPlugin_logic_DATA_lane0 : 32'h0)) | ((_zz_toplevel_execute_ctrl2_integer_RS1_lane0_bypass[2] ? toplevel_execute_ctrl4_down_lane0_integer_WriteBackPlugin_logic_DATA_lane0 : 32'h0) | (_zz_toplevel_execute_ctrl2_integer_RS1_lane0_bypass[3] ? toplevel_execute_ctrl3_down_lane1_integer_WriteBackPlugin_logic_DATA_lane1 : 32'h0))) | (_zz_toplevel_execute_ctrl2_integer_RS1_lane0_bypass[4] ? toplevel_execute_ctrl4_down_lane1_integer_WriteBackPlugin_logic_DATA_lane1 : 32'h0));
  assign toplevel_execute_lane0_bypasser_integer_RS1_along_bypasses_1_checks_0_selfHit = (((toplevel_execute_ctrl4_up_LANE_SEL_lane0 && toplevel_execute_ctrl4_up_RD_ENABLE_lane0) && (toplevel_execute_ctrl4_down_RD_PHYS_lane0 == toplevel_execute_ctrl3_down_RS1_PHYS_lane0)) && 1'b1);
  assign toplevel_execute_lane0_bypasser_integer_RS1_along_bypasses_1_checks_0_hit = (toplevel_execute_lane0_bypasser_integer_RS1_along_bypasses_1_checks_0_selfHit && (! 1'b0));
  assign toplevel_execute_lane0_bypasser_integer_RS1_along_bypasses_1_checks_1_selfHit = (((toplevel_execute_ctrl4_up_LANE_SEL_lane1 && toplevel_execute_ctrl4_up_RD_ENABLE_lane1) && (toplevel_execute_ctrl4_down_RD_PHYS_lane1 == toplevel_execute_ctrl3_down_RS1_PHYS_lane0)) && 1'b1);
  assign toplevel_execute_lane0_bypasser_integer_RS1_along_bypasses_1_checks_1_hit = (toplevel_execute_lane0_bypasser_integer_RS1_along_bypasses_1_checks_1_selfHit && (! 1'b0));
  assign toplevel_execute_lane0_bypasser_integer_RS1_along_bypasses_1_hits = {toplevel_execute_lane0_bypasser_integer_RS1_along_bypasses_1_checks_1_hit,toplevel_execute_lane0_bypasser_integer_RS1_along_bypasses_1_checks_0_hit};
  assign _zz_toplevel_execute_ctrl3_integer_RS1_lane0_bypass = {toplevel_execute_lane0_bypasser_integer_RS1_along_bypasses_1_hits,(! (|toplevel_execute_lane0_bypasser_integer_RS1_along_bypasses_1_hits))};
  assign toplevel_execute_ctrl3_integer_RS1_lane0_bypass = (((_zz_toplevel_execute_ctrl3_integer_RS1_lane0_bypass[0] ? toplevel_execute_ctrl3_up_integer_RS1_lane0 : 32'h0) | (_zz_toplevel_execute_ctrl3_integer_RS1_lane0_bypass[1] ? toplevel_execute_ctrl4_down_lane0_integer_WriteBackPlugin_logic_DATA_lane0 : 32'h0)) | (_zz_toplevel_execute_ctrl3_integer_RS1_lane0_bypass[2] ? toplevel_execute_ctrl4_down_lane1_integer_WriteBackPlugin_logic_DATA_lane1 : 32'h0));
  assign toplevel_execute_lane0_bypasser_integer_RS2_port_valid = (! execute_freeze_valid);
  assign toplevel_execute_lane0_bypasser_integer_RS2_port_address = toplevel_execute_ctrl0_down_RS2_PHYS_lane0;
  always @(*) begin
    toplevel_execute_lane0_bypasser_integer_RS2_bypassEnables[0] = (((toplevel_execute_ctrl2_up_LANE_SEL_lane0 && toplevel_execute_ctrl2_up_RD_ENABLE_lane0) && (toplevel_execute_ctrl2_down_RD_PHYS_lane0 == toplevel_execute_ctrl1_down_RS2_PHYS_lane0)) && 1'b1);
    toplevel_execute_lane0_bypasser_integer_RS2_bypassEnables[1] = (((toplevel_execute_ctrl2_up_LANE_SEL_lane1 && toplevel_execute_ctrl2_up_RD_ENABLE_lane1) && (toplevel_execute_ctrl2_down_RD_PHYS_lane1 == toplevel_execute_ctrl1_down_RS2_PHYS_lane0)) && 1'b1);
    toplevel_execute_lane0_bypasser_integer_RS2_bypassEnables[2] = (((toplevel_execute_ctrl3_up_LANE_SEL_lane0 && toplevel_execute_ctrl3_up_RD_ENABLE_lane0) && (toplevel_execute_ctrl3_down_RD_PHYS_lane0 == toplevel_execute_ctrl1_down_RS2_PHYS_lane0)) && 1'b1);
    toplevel_execute_lane0_bypasser_integer_RS2_bypassEnables[3] = (((toplevel_execute_ctrl3_up_LANE_SEL_lane1 && toplevel_execute_ctrl3_up_RD_ENABLE_lane1) && (toplevel_execute_ctrl3_down_RD_PHYS_lane1 == toplevel_execute_ctrl1_down_RS2_PHYS_lane0)) && 1'b1);
    toplevel_execute_lane0_bypasser_integer_RS2_bypassEnables[4] = (((toplevel_execute_ctrl4_up_LANE_SEL_lane0 && toplevel_execute_ctrl4_up_RD_ENABLE_lane0) && (toplevel_execute_ctrl4_down_RD_PHYS_lane0 == toplevel_execute_ctrl1_down_RS2_PHYS_lane0)) && 1'b1);
    toplevel_execute_lane0_bypasser_integer_RS2_bypassEnables[5] = (((toplevel_execute_ctrl4_up_LANE_SEL_lane1 && toplevel_execute_ctrl4_up_RD_ENABLE_lane1) && (toplevel_execute_ctrl4_down_RD_PHYS_lane1 == toplevel_execute_ctrl1_down_RS2_PHYS_lane0)) && 1'b1);
    toplevel_execute_lane0_bypasser_integer_RS2_bypassEnables[6] = (((toplevel_execute_ctrl5_up_LANE_SEL_lane0 && toplevel_execute_ctrl5_up_RD_ENABLE_lane0) && (toplevel_execute_ctrl5_down_RD_PHYS_lane0 == toplevel_execute_ctrl1_down_RS2_PHYS_lane0)) && 1'b1);
    toplevel_execute_lane0_bypasser_integer_RS2_bypassEnables[7] = (((toplevel_execute_ctrl5_up_LANE_SEL_lane1 && toplevel_execute_ctrl5_up_RD_ENABLE_lane1) && (toplevel_execute_ctrl5_down_RD_PHYS_lane1 == toplevel_execute_ctrl1_down_RS2_PHYS_lane0)) && 1'b1);
    toplevel_execute_lane0_bypasser_integer_RS2_bypassEnables[8] = 1'b1;
  end

  assign _zz_toplevel_execute_lane0_bypasser_integer_RS2_bypassEnables_bools_0 = toplevel_execute_lane0_bypasser_integer_RS2_bypassEnables;
  assign toplevel_execute_lane0_bypasser_integer_RS2_bypassEnables_bools_0 = _zz_toplevel_execute_lane0_bypasser_integer_RS2_bypassEnables_bools_0[0];
  assign toplevel_execute_lane0_bypasser_integer_RS2_bypassEnables_bools_1 = _zz_toplevel_execute_lane0_bypasser_integer_RS2_bypassEnables_bools_0[1];
  assign toplevel_execute_lane0_bypasser_integer_RS2_bypassEnables_bools_2 = _zz_toplevel_execute_lane0_bypasser_integer_RS2_bypassEnables_bools_0[2];
  assign toplevel_execute_lane0_bypasser_integer_RS2_bypassEnables_bools_3 = _zz_toplevel_execute_lane0_bypasser_integer_RS2_bypassEnables_bools_0[3];
  assign toplevel_execute_lane0_bypasser_integer_RS2_bypassEnables_bools_4 = _zz_toplevel_execute_lane0_bypasser_integer_RS2_bypassEnables_bools_0[4];
  assign toplevel_execute_lane0_bypasser_integer_RS2_bypassEnables_bools_5 = _zz_toplevel_execute_lane0_bypasser_integer_RS2_bypassEnables_bools_0[5];
  assign toplevel_execute_lane0_bypasser_integer_RS2_bypassEnables_bools_6 = _zz_toplevel_execute_lane0_bypasser_integer_RS2_bypassEnables_bools_0[6];
  assign toplevel_execute_lane0_bypasser_integer_RS2_bypassEnables_bools_7 = _zz_toplevel_execute_lane0_bypasser_integer_RS2_bypassEnables_bools_0[7];
  assign toplevel_execute_lane0_bypasser_integer_RS2_bypassEnables_bools_8 = _zz_toplevel_execute_lane0_bypasser_integer_RS2_bypassEnables_bools_0[8];
  always @(*) begin
    _zz_toplevel_execute_lane0_bypasser_integer_RS2_sel[0] = (toplevel_execute_lane0_bypasser_integer_RS2_bypassEnables_bools_0 && (! 1'b0));
    _zz_toplevel_execute_lane0_bypasser_integer_RS2_sel[1] = (toplevel_execute_lane0_bypasser_integer_RS2_bypassEnables_bools_1 && (! toplevel_execute_lane0_bypasser_integer_RS2_bypassEnables_bools_0));
    _zz_toplevel_execute_lane0_bypasser_integer_RS2_sel[2] = (toplevel_execute_lane0_bypasser_integer_RS2_bypassEnables_bools_2 && (! toplevel_execute_lane0_bypasser_integer_RS2_bypassEnables_range_0_to_1));
    _zz_toplevel_execute_lane0_bypasser_integer_RS2_sel[3] = (toplevel_execute_lane0_bypasser_integer_RS2_bypassEnables_bools_3 && (! toplevel_execute_lane0_bypasser_integer_RS2_bypassEnables_range_0_to_2));
    _zz_toplevel_execute_lane0_bypasser_integer_RS2_sel[4] = (toplevel_execute_lane0_bypasser_integer_RS2_bypassEnables_bools_4 && (! toplevel_execute_lane0_bypasser_integer_RS2_bypassEnables_range_0_to_3));
    _zz_toplevel_execute_lane0_bypasser_integer_RS2_sel[5] = (toplevel_execute_lane0_bypasser_integer_RS2_bypassEnables_bools_5 && (! (toplevel_execute_lane0_bypasser_integer_RS2_bypassEnables_bools_4 || toplevel_execute_lane0_bypasser_integer_RS2_bypassEnables_range_0_to_3)));
    _zz_toplevel_execute_lane0_bypasser_integer_RS2_sel[6] = (toplevel_execute_lane0_bypasser_integer_RS2_bypassEnables_bools_6 && (! (toplevel_execute_lane0_bypasser_integer_RS2_bypassEnables_range_4_to_5 || toplevel_execute_lane0_bypasser_integer_RS2_bypassEnables_range_0_to_3)));
    _zz_toplevel_execute_lane0_bypasser_integer_RS2_sel[7] = (toplevel_execute_lane0_bypasser_integer_RS2_bypassEnables_bools_7 && (! (toplevel_execute_lane0_bypasser_integer_RS2_bypassEnables_range_4_to_6 || toplevel_execute_lane0_bypasser_integer_RS2_bypassEnables_range_0_to_3)));
    _zz_toplevel_execute_lane0_bypasser_integer_RS2_sel[8] = (toplevel_execute_lane0_bypasser_integer_RS2_bypassEnables_bools_8 && (! (toplevel_execute_lane0_bypasser_integer_RS2_bypassEnables_range_4_to_7 || toplevel_execute_lane0_bypasser_integer_RS2_bypassEnables_range_0_to_3)));
  end

  assign toplevel_execute_lane0_bypasser_integer_RS2_bypassEnables_range_0_to_1 = (|{toplevel_execute_lane0_bypasser_integer_RS2_bypassEnables_bools_1,toplevel_execute_lane0_bypasser_integer_RS2_bypassEnables_bools_0});
  assign toplevel_execute_lane0_bypasser_integer_RS2_bypassEnables_range_0_to_2 = (|{toplevel_execute_lane0_bypasser_integer_RS2_bypassEnables_bools_2,{toplevel_execute_lane0_bypasser_integer_RS2_bypassEnables_bools_1,toplevel_execute_lane0_bypasser_integer_RS2_bypassEnables_bools_0}});
  assign toplevel_execute_lane0_bypasser_integer_RS2_bypassEnables_range_0_to_3 = (|{toplevel_execute_lane0_bypasser_integer_RS2_bypassEnables_bools_3,{toplevel_execute_lane0_bypasser_integer_RS2_bypassEnables_bools_2,{toplevel_execute_lane0_bypasser_integer_RS2_bypassEnables_bools_1,toplevel_execute_lane0_bypasser_integer_RS2_bypassEnables_bools_0}}});
  assign toplevel_execute_lane0_bypasser_integer_RS2_bypassEnables_range_4_to_5 = (|{toplevel_execute_lane0_bypasser_integer_RS2_bypassEnables_bools_5,toplevel_execute_lane0_bypasser_integer_RS2_bypassEnables_bools_4});
  assign toplevel_execute_lane0_bypasser_integer_RS2_bypassEnables_range_4_to_6 = (|{toplevel_execute_lane0_bypasser_integer_RS2_bypassEnables_bools_6,{toplevel_execute_lane0_bypasser_integer_RS2_bypassEnables_bools_5,toplevel_execute_lane0_bypasser_integer_RS2_bypassEnables_bools_4}});
  assign toplevel_execute_lane0_bypasser_integer_RS2_bypassEnables_range_4_to_7 = (|{toplevel_execute_lane0_bypasser_integer_RS2_bypassEnables_bools_7,{toplevel_execute_lane0_bypasser_integer_RS2_bypassEnables_bools_6,{toplevel_execute_lane0_bypasser_integer_RS2_bypassEnables_bools_5,toplevel_execute_lane0_bypasser_integer_RS2_bypassEnables_bools_4}}});
  assign toplevel_execute_lane0_bypasser_integer_RS2_sel = _zz_toplevel_execute_lane0_bypasser_integer_RS2_sel;
  assign _zz_toplevel_execute_ctrl1_down_integer_RS2_lane0 = toplevel_execute_lane0_bypasser_integer_RS2_sel[8 : 1];
  always @(*) begin
    _zz_toplevel_execute_ctrl1_down_integer_RS2_lane0_1 = ((((_zz__zz_toplevel_execute_ctrl1_down_integer_RS2_lane0_1 ? toplevel_execute_ctrl2_down_lane1_integer_WriteBackPlugin_logic_DATA_lane1 : _zz__zz_toplevel_execute_ctrl1_down_integer_RS2_lane0_1_1) | (_zz__zz_toplevel_execute_ctrl1_down_integer_RS2_lane0_1_2 ? toplevel_execute_ctrl3_down_lane0_integer_WriteBackPlugin_logic_DATA_lane0 : _zz__zz_toplevel_execute_ctrl1_down_integer_RS2_lane0_1_3)) | ((_zz__zz_toplevel_execute_ctrl1_down_integer_RS2_lane0_1_4 ? toplevel_execute_ctrl3_down_lane1_integer_WriteBackPlugin_logic_DATA_lane1 : _zz__zz_toplevel_execute_ctrl1_down_integer_RS2_lane0_1_5) | (_zz__zz_toplevel_execute_ctrl1_down_integer_RS2_lane0_1_6 ? toplevel_execute_ctrl4_down_lane0_integer_WriteBackPlugin_logic_DATA_lane0 : _zz__zz_toplevel_execute_ctrl1_down_integer_RS2_lane0_1_7))) | (((_zz__zz_toplevel_execute_ctrl1_down_integer_RS2_lane0_1_8 ? toplevel_execute_ctrl4_down_lane1_integer_WriteBackPlugin_logic_DATA_lane1 : _zz__zz_toplevel_execute_ctrl1_down_integer_RS2_lane0_1_9) | (_zz__zz_toplevel_execute_ctrl1_down_integer_RS2_lane0_1_10 ? toplevel_execute_ctrl5_down_lane0_integer_WriteBackPlugin_logic_DATA_lane0 : _zz__zz_toplevel_execute_ctrl1_down_integer_RS2_lane0_1_11)) | ((_zz__zz_toplevel_execute_ctrl1_down_integer_RS2_lane0_1_12 ? toplevel_execute_ctrl5_down_lane1_integer_WriteBackPlugin_logic_DATA_lane1 : _zz__zz_toplevel_execute_ctrl1_down_integer_RS2_lane0_1_13) | (_zz__zz_toplevel_execute_ctrl1_down_integer_RS2_lane0_1_14 ? toplevel_execute_lane0_bypasser_integer_RS2_port_data : _zz__zz_toplevel_execute_ctrl1_down_integer_RS2_lane0_1_15))));
    if(when_ExecuteLanePlugin_l190_1) begin
      _zz_toplevel_execute_ctrl1_down_integer_RS2_lane0_1 = toplevel_execute_ctrl2_down_lane0_integer_WriteBackPlugin_logic_DATA_lane0;
    end
  end

  assign toplevel_execute_ctrl1_down_integer_RS2_lane0 = _zz_toplevel_execute_ctrl1_down_integer_RS2_lane0_1;
  assign when_ExecuteLanePlugin_l190_1 = toplevel_execute_lane0_bypasser_integer_RS2_sel[0];
  assign toplevel_execute_lane0_bypasser_integer_RS2_along_bypasses_0_checks_0_selfHit = (((toplevel_execute_ctrl3_up_LANE_SEL_lane0 && toplevel_execute_ctrl3_up_RD_ENABLE_lane0) && (toplevel_execute_ctrl3_down_RD_PHYS_lane0 == toplevel_execute_ctrl2_down_RS2_PHYS_lane0)) && 1'b1);
  assign toplevel_execute_lane0_bypasser_integer_RS2_along_bypasses_0_checks_0_hit = (toplevel_execute_lane0_bypasser_integer_RS2_along_bypasses_0_checks_0_selfHit && (! 1'b0));
  assign toplevel_execute_lane0_bypasser_integer_RS2_along_bypasses_0_checks_1_selfHit = (((toplevel_execute_ctrl4_up_LANE_SEL_lane0 && toplevel_execute_ctrl4_up_RD_ENABLE_lane0) && (toplevel_execute_ctrl4_down_RD_PHYS_lane0 == toplevel_execute_ctrl2_down_RS2_PHYS_lane0)) && 1'b1);
  assign toplevel_execute_lane0_bypasser_integer_RS2_along_bypasses_0_checks_1_youngerHits_0 = (((toplevel_execute_ctrl3_up_LANE_SEL_lane0 && toplevel_execute_ctrl3_up_RD_ENABLE_lane0) && (toplevel_execute_ctrl3_down_RD_PHYS_lane0 == toplevel_execute_ctrl2_down_RS2_PHYS_lane0)) && 1'b1);
  assign toplevel_execute_lane0_bypasser_integer_RS2_along_bypasses_0_checks_1_youngerHits_1 = (((toplevel_execute_ctrl3_up_LANE_SEL_lane1 && toplevel_execute_ctrl3_up_RD_ENABLE_lane1) && (toplevel_execute_ctrl3_down_RD_PHYS_lane1 == toplevel_execute_ctrl2_down_RS2_PHYS_lane0)) && 1'b1);
  assign toplevel_execute_lane0_bypasser_integer_RS2_along_bypasses_0_checks_1_hit = (toplevel_execute_lane0_bypasser_integer_RS2_along_bypasses_0_checks_1_selfHit && (! (|{toplevel_execute_lane0_bypasser_integer_RS2_along_bypasses_0_checks_1_youngerHits_1,toplevel_execute_lane0_bypasser_integer_RS2_along_bypasses_0_checks_1_youngerHits_0})));
  assign toplevel_execute_lane0_bypasser_integer_RS2_along_bypasses_0_checks_2_selfHit = (((toplevel_execute_ctrl3_up_LANE_SEL_lane1 && toplevel_execute_ctrl3_up_RD_ENABLE_lane1) && (toplevel_execute_ctrl3_down_RD_PHYS_lane1 == toplevel_execute_ctrl2_down_RS2_PHYS_lane0)) && 1'b1);
  assign toplevel_execute_lane0_bypasser_integer_RS2_along_bypasses_0_checks_2_hit = (toplevel_execute_lane0_bypasser_integer_RS2_along_bypasses_0_checks_2_selfHit && (! 1'b0));
  assign toplevel_execute_lane0_bypasser_integer_RS2_along_bypasses_0_checks_3_selfHit = (((toplevel_execute_ctrl4_up_LANE_SEL_lane1 && toplevel_execute_ctrl4_up_RD_ENABLE_lane1) && (toplevel_execute_ctrl4_down_RD_PHYS_lane1 == toplevel_execute_ctrl2_down_RS2_PHYS_lane0)) && 1'b1);
  assign toplevel_execute_lane0_bypasser_integer_RS2_along_bypasses_0_checks_3_youngerHits_0 = (((toplevel_execute_ctrl3_up_LANE_SEL_lane0 && toplevel_execute_ctrl3_up_RD_ENABLE_lane0) && (toplevel_execute_ctrl3_down_RD_PHYS_lane0 == toplevel_execute_ctrl2_down_RS2_PHYS_lane0)) && 1'b1);
  assign toplevel_execute_lane0_bypasser_integer_RS2_along_bypasses_0_checks_3_youngerHits_1 = (((toplevel_execute_ctrl3_up_LANE_SEL_lane1 && toplevel_execute_ctrl3_up_RD_ENABLE_lane1) && (toplevel_execute_ctrl3_down_RD_PHYS_lane1 == toplevel_execute_ctrl2_down_RS2_PHYS_lane0)) && 1'b1);
  assign toplevel_execute_lane0_bypasser_integer_RS2_along_bypasses_0_checks_3_hit = (toplevel_execute_lane0_bypasser_integer_RS2_along_bypasses_0_checks_3_selfHit && (! (|{toplevel_execute_lane0_bypasser_integer_RS2_along_bypasses_0_checks_3_youngerHits_1,toplevel_execute_lane0_bypasser_integer_RS2_along_bypasses_0_checks_3_youngerHits_0})));
  assign toplevel_execute_lane0_bypasser_integer_RS2_along_bypasses_0_hits = {toplevel_execute_lane0_bypasser_integer_RS2_along_bypasses_0_checks_3_hit,{toplevel_execute_lane0_bypasser_integer_RS2_along_bypasses_0_checks_2_hit,{toplevel_execute_lane0_bypasser_integer_RS2_along_bypasses_0_checks_1_hit,toplevel_execute_lane0_bypasser_integer_RS2_along_bypasses_0_checks_0_hit}}};
  assign _zz_toplevel_execute_ctrl2_integer_RS2_lane0_bypass = {toplevel_execute_lane0_bypasser_integer_RS2_along_bypasses_0_hits,(! (|toplevel_execute_lane0_bypasser_integer_RS2_along_bypasses_0_hits))};
  assign toplevel_execute_ctrl2_integer_RS2_lane0_bypass = ((((_zz_toplevel_execute_ctrl2_integer_RS2_lane0_bypass[0] ? toplevel_execute_ctrl2_up_integer_RS2_lane0 : 32'h0) | (_zz_toplevel_execute_ctrl2_integer_RS2_lane0_bypass[1] ? toplevel_execute_ctrl3_down_lane0_integer_WriteBackPlugin_logic_DATA_lane0 : 32'h0)) | ((_zz_toplevel_execute_ctrl2_integer_RS2_lane0_bypass[2] ? toplevel_execute_ctrl4_down_lane0_integer_WriteBackPlugin_logic_DATA_lane0 : 32'h0) | (_zz_toplevel_execute_ctrl2_integer_RS2_lane0_bypass[3] ? toplevel_execute_ctrl3_down_lane1_integer_WriteBackPlugin_logic_DATA_lane1 : 32'h0))) | (_zz_toplevel_execute_ctrl2_integer_RS2_lane0_bypass[4] ? toplevel_execute_ctrl4_down_lane1_integer_WriteBackPlugin_logic_DATA_lane1 : 32'h0));
  assign toplevel_execute_lane0_bypasser_integer_RS2_along_bypasses_1_checks_0_selfHit = (((toplevel_execute_ctrl4_up_LANE_SEL_lane0 && toplevel_execute_ctrl4_up_RD_ENABLE_lane0) && (toplevel_execute_ctrl4_down_RD_PHYS_lane0 == toplevel_execute_ctrl3_down_RS2_PHYS_lane0)) && 1'b1);
  assign toplevel_execute_lane0_bypasser_integer_RS2_along_bypasses_1_checks_0_hit = (toplevel_execute_lane0_bypasser_integer_RS2_along_bypasses_1_checks_0_selfHit && (! 1'b0));
  assign toplevel_execute_lane0_bypasser_integer_RS2_along_bypasses_1_checks_1_selfHit = (((toplevel_execute_ctrl4_up_LANE_SEL_lane1 && toplevel_execute_ctrl4_up_RD_ENABLE_lane1) && (toplevel_execute_ctrl4_down_RD_PHYS_lane1 == toplevel_execute_ctrl3_down_RS2_PHYS_lane0)) && 1'b1);
  assign toplevel_execute_lane0_bypasser_integer_RS2_along_bypasses_1_checks_1_hit = (toplevel_execute_lane0_bypasser_integer_RS2_along_bypasses_1_checks_1_selfHit && (! 1'b0));
  assign toplevel_execute_lane0_bypasser_integer_RS2_along_bypasses_1_hits = {toplevel_execute_lane0_bypasser_integer_RS2_along_bypasses_1_checks_1_hit,toplevel_execute_lane0_bypasser_integer_RS2_along_bypasses_1_checks_0_hit};
  assign _zz_toplevel_execute_ctrl3_integer_RS2_lane0_bypass = {toplevel_execute_lane0_bypasser_integer_RS2_along_bypasses_1_hits,(! (|toplevel_execute_lane0_bypasser_integer_RS2_along_bypasses_1_hits))};
  assign toplevel_execute_ctrl3_integer_RS2_lane0_bypass = (((_zz_toplevel_execute_ctrl3_integer_RS2_lane0_bypass[0] ? toplevel_execute_ctrl3_up_integer_RS2_lane0 : 32'h0) | (_zz_toplevel_execute_ctrl3_integer_RS2_lane0_bypass[1] ? toplevel_execute_ctrl4_down_lane0_integer_WriteBackPlugin_logic_DATA_lane0 : 32'h0)) | (_zz_toplevel_execute_ctrl3_integer_RS2_lane0_bypass[2] ? toplevel_execute_ctrl4_down_lane1_integer_WriteBackPlugin_logic_DATA_lane1 : 32'h0));
  assign execute_lane0_logic_completions_onCtrl_0_port_valid = (((toplevel_execute_ctrl2_down_LANE_SEL_lane0 && toplevel_execute_ctrl2_down_isReady) && (! toplevel_execute_lane0_ctrls_2_downIsCancel)) && toplevel_execute_ctrl2_down_execute_lane0_logic_completions_onCtrl_0_ENABLE_lane0);
  assign execute_lane0_logic_completions_onCtrl_0_port_payload_uopId = toplevel_execute_ctrl2_down_Decode_UOP_ID_lane0;
  assign execute_lane0_logic_completions_onCtrl_0_port_payload_trap = toplevel_execute_ctrl2_down_TRAP_lane0;
  assign execute_lane0_logic_completions_onCtrl_0_port_payload_commit = toplevel_execute_ctrl2_down_COMMIT_lane0;
  assign execute_lane0_logic_completions_onCtrl_1_port_valid = (((toplevel_execute_ctrl3_down_LANE_SEL_lane0 && toplevel_execute_ctrl3_down_isReady) && (! toplevel_execute_lane0_ctrls_3_downIsCancel)) && toplevel_execute_ctrl3_down_execute_lane0_logic_completions_onCtrl_1_ENABLE_lane0);
  assign execute_lane0_logic_completions_onCtrl_1_port_payload_uopId = toplevel_execute_ctrl3_down_Decode_UOP_ID_lane0;
  assign execute_lane0_logic_completions_onCtrl_1_port_payload_trap = toplevel_execute_ctrl3_down_TRAP_lane0;
  assign execute_lane0_logic_completions_onCtrl_1_port_payload_commit = toplevel_execute_ctrl3_down_COMMIT_lane0;
  assign execute_lane0_logic_completions_onCtrl_2_port_valid = (((toplevel_execute_ctrl4_down_LANE_SEL_lane0 && toplevel_execute_ctrl4_down_isReady) && (! toplevel_execute_lane0_ctrls_4_downIsCancel)) && toplevel_execute_ctrl4_down_execute_lane0_logic_completions_onCtrl_2_ENABLE_lane0);
  assign execute_lane0_logic_completions_onCtrl_2_port_payload_uopId = toplevel_execute_ctrl4_down_Decode_UOP_ID_lane0;
  assign execute_lane0_logic_completions_onCtrl_2_port_payload_trap = toplevel_execute_ctrl4_down_TRAP_lane0;
  assign execute_lane0_logic_completions_onCtrl_2_port_payload_commit = toplevel_execute_ctrl4_down_COMMIT_lane0;
  assign execute_lane0_logic_decoding_decodingBits = {toplevel_execute_ctrl1_down_execute_lane0_LAYER_SEL_lane0,toplevel_execute_ctrl1_down_Decode_UOP_lane0};
  assign _zz_toplevel_execute_ctrl1_down_execute_lane0_logic_completions_onCtrl_0_ENABLE_lane0 = ((execute_lane0_logic_decoding_decodingBits & 33'h102002050) == 33'h100002010);
  assign _zz_toplevel_execute_ctrl1_down_execute_lane0_logic_completions_onCtrl_0_ENABLE_lane0_1 = ((execute_lane0_logic_decoding_decodingBits & 33'h100001030) == 33'h100000010);
  assign _zz_toplevel_execute_ctrl1_down_execute_lane0_logic_completions_onCtrl_0_ENABLE_lane0_2 = ((execute_lane0_logic_decoding_decodingBits & 33'h10000004c) == 33'h100000004);
  assign _zz_toplevel_execute_ctrl1_down_execute_lane0_logic_completions_onCtrl_0_ENABLE_lane0_3 = ((execute_lane0_logic_decoding_decodingBits & 33'h100002030) == 33'h100002010);
  always @(*) begin
    toplevel_execute_ctrl1_down_early0_IntAluPlugin_SEL_lane0 = _zz_toplevel_execute_ctrl1_down_early0_IntAluPlugin_SEL_lane0[0];
    if(toplevel_execute_ctrl1_down_TRAP_lane0) begin
      toplevel_execute_ctrl1_down_early0_IntAluPlugin_SEL_lane0 = 1'b0;
    end
  end

  assign _zz_toplevel_execute_ctrl1_down_execute_lane0_logic_completions_onCtrl_1_ENABLE_lane0 = ((execute_lane0_logic_decoding_decodingBits & 33'h100003034) == 33'h100001010);
  always @(*) begin
    toplevel_execute_ctrl1_down_early0_BarrelShifterPlugin_SEL_lane0 = _zz_toplevel_execute_ctrl1_down_early0_BarrelShifterPlugin_SEL_lane0[0];
    if(toplevel_execute_ctrl1_down_TRAP_lane0) begin
      toplevel_execute_ctrl1_down_early0_BarrelShifterPlugin_SEL_lane0 = 1'b0;
    end
  end

  assign _zz_toplevel_execute_ctrl1_down_execute_lane0_logic_completions_onCtrl_1_ENABLE_lane0_1 = ((execute_lane0_logic_decoding_decodingBits & 33'h100000050) == 33'h100000040);
  always @(*) begin
    toplevel_execute_ctrl1_down_early0_BranchPlugin_SEL_lane0 = _zz_toplevel_execute_ctrl1_down_early0_BranchPlugin_SEL_lane0[0];
    if(toplevel_execute_ctrl1_down_TRAP_lane0) begin
      toplevel_execute_ctrl1_down_early0_BranchPlugin_SEL_lane0 = 1'b0;
    end
  end

  always @(*) begin
    toplevel_execute_ctrl1_down_early0_MulPlugin_SEL_lane0 = _zz_toplevel_execute_ctrl1_down_early0_MulPlugin_SEL_lane0[0];
    if(toplevel_execute_ctrl1_down_TRAP_lane0) begin
      toplevel_execute_ctrl1_down_early0_MulPlugin_SEL_lane0 = 1'b0;
    end
  end

  assign _zz_toplevel_execute_ctrl1_down_execute_lane0_logic_completions_onCtrl_1_ENABLE_lane0_2 = ((execute_lane0_logic_decoding_decodingBits & 33'h002004064) == 33'h002004020);
  always @(*) begin
    toplevel_execute_ctrl1_down_early0_DivPlugin_SEL_lane0 = _zz_toplevel_execute_ctrl1_down_early0_DivPlugin_SEL_lane0[0];
    if(toplevel_execute_ctrl1_down_TRAP_lane0) begin
      toplevel_execute_ctrl1_down_early0_DivPlugin_SEL_lane0 = 1'b0;
    end
  end

  assign _zz_toplevel_execute_ctrl1_down_execute_lane0_logic_completions_onCtrl_0_ENABLE_lane0_4 = ((execute_lane0_logic_decoding_decodingBits & 33'h000001048) == 33'h000001008);
  always @(*) begin
    toplevel_execute_ctrl1_down_early0_EnvPlugin_SEL_lane0 = _zz_toplevel_execute_ctrl1_down_early0_EnvPlugin_SEL_lane0[0];
    if(toplevel_execute_ctrl1_down_TRAP_lane0) begin
      toplevel_execute_ctrl1_down_early0_EnvPlugin_SEL_lane0 = 1'b0;
    end
  end

  always @(*) begin
    toplevel_execute_ctrl1_down_late0_IntAluPlugin_SEL_lane0 = _zz_toplevel_execute_ctrl1_down_late0_IntAluPlugin_SEL_lane0[0];
    if(toplevel_execute_ctrl1_down_TRAP_lane0) begin
      toplevel_execute_ctrl1_down_late0_IntAluPlugin_SEL_lane0 = 1'b0;
    end
  end

  always @(*) begin
    toplevel_execute_ctrl1_down_late0_BarrelShifterPlugin_SEL_lane0 = _zz_toplevel_execute_ctrl1_down_late0_BarrelShifterPlugin_SEL_lane0[0];
    if(toplevel_execute_ctrl1_down_TRAP_lane0) begin
      toplevel_execute_ctrl1_down_late0_BarrelShifterPlugin_SEL_lane0 = 1'b0;
    end
  end

  assign _zz_toplevel_execute_ctrl1_down_late0_BranchPlugin_SEL_lane0 = ((execute_lane0_logic_decoding_decodingBits & 33'h100000010) == 33'h0);
  always @(*) begin
    toplevel_execute_ctrl1_down_late0_BranchPlugin_SEL_lane0 = _zz_toplevel_execute_ctrl1_down_late0_BranchPlugin_SEL_lane0_1[0];
    if(toplevel_execute_ctrl1_down_TRAP_lane0) begin
      toplevel_execute_ctrl1_down_late0_BranchPlugin_SEL_lane0 = 1'b0;
    end
  end

  always @(*) begin
    toplevel_execute_ctrl1_down_MulPlugin_HIGH_lane0 = _zz_toplevel_execute_ctrl1_down_MulPlugin_HIGH_lane0[0];
    if(toplevel_execute_ctrl1_down_TRAP_lane0) begin
      toplevel_execute_ctrl1_down_MulPlugin_HIGH_lane0 = 1'b0;
    end
  end

  always @(*) begin
    toplevel_execute_ctrl1_down_CsrAccessPlugin_SEL_lane0 = _zz_toplevel_execute_ctrl1_down_CsrAccessPlugin_SEL_lane0[0];
    if(toplevel_execute_ctrl1_down_TRAP_lane0) begin
      toplevel_execute_ctrl1_down_CsrAccessPlugin_SEL_lane0 = 1'b0;
    end
  end

  assign _zz_toplevel_execute_ctrl1_down_execute_lane0_logic_completions_onCtrl_2_ENABLE_lane0 = ((execute_lane0_logic_decoding_decodingBits & 33'h000000058) == 33'h0);
  assign _zz_toplevel_execute_ctrl1_down_execute_lane0_logic_completions_onCtrl_2_ENABLE_lane0_1 = ((execute_lane0_logic_decoding_decodingBits & 33'h000001050) == 33'h0);
  always @(*) begin
    toplevel_execute_ctrl1_down_AguPlugin_SEL_lane0 = _zz_toplevel_execute_ctrl1_down_AguPlugin_SEL_lane0[0];
    if(toplevel_execute_ctrl1_down_TRAP_lane0) begin
      toplevel_execute_ctrl1_down_AguPlugin_SEL_lane0 = 1'b0;
    end
  end

  always @(*) begin
    toplevel_execute_ctrl1_down_LsuPlugin_logic_FENCE_lane0 = _zz_toplevel_execute_ctrl1_down_LsuPlugin_logic_FENCE_lane0[0];
    if(toplevel_execute_ctrl1_down_TRAP_lane0) begin
      toplevel_execute_ctrl1_down_LsuPlugin_logic_FENCE_lane0 = 1'b0;
    end
  end

  assign _zz_toplevel_execute_ctrl1_down_AguPlugin_LOAD_lane0 = ((execute_lane0_logic_decoding_decodingBits & 33'h000000028) == 33'h0);
  assign _zz_toplevel_execute_ctrl1_down_lane0_integer_WriteBackPlugin_SEL_lane0 = ((execute_lane0_logic_decoding_decodingBits & 33'h00000000c) == 33'h000000004);
  assign _zz_toplevel_execute_ctrl1_down_AguPlugin_ATOMIC_lane0 = ((execute_lane0_logic_decoding_decodingBits & 33'h000002008) == 33'h000002008);
  always @(*) begin
    toplevel_execute_ctrl1_down_lane0_integer_WriteBackPlugin_SEL_lane0 = _zz_toplevel_execute_ctrl1_down_lane0_integer_WriteBackPlugin_SEL_lane0_1[0];
    if(toplevel_execute_ctrl1_down_TRAP_lane0) begin
      toplevel_execute_ctrl1_down_lane0_integer_WriteBackPlugin_SEL_lane0 = 1'b0;
    end
  end

  assign _zz_toplevel_execute_ctrl1_down_execute_lane0_logic_completions_onCtrl_0_ENABLE_lane0_5 = ((execute_lane0_logic_decoding_decodingBits & 33'h102003010) == 33'h100000010);
  assign _zz_toplevel_execute_ctrl1_down_execute_lane0_logic_completions_onCtrl_0_ENABLE_lane0_6 = ((execute_lane0_logic_decoding_decodingBits & 33'h110003010) == 33'h110000010);
  always @(*) begin
    toplevel_execute_ctrl1_down_COMPLETION_AT_2_lane0 = _zz_toplevel_execute_ctrl1_down_COMPLETION_AT_2_lane0[0];
    if(toplevel_execute_ctrl1_down_TRAP_lane0) begin
      toplevel_execute_ctrl1_down_COMPLETION_AT_2_lane0 = 1'b0;
    end
  end

  assign _zz_toplevel_execute_ctrl1_down_execute_lane0_logic_completions_onCtrl_1_ENABLE_lane0_3 = ((execute_lane0_logic_decoding_decodingBits & 33'h102003014) == 33'h100001010);
  assign _zz_toplevel_execute_ctrl1_down_execute_lane0_logic_completions_onCtrl_1_ENABLE_lane0_4 = ((execute_lane0_logic_decoding_decodingBits & 33'h100001040) == 33'h100001040);
  assign _zz_toplevel_execute_ctrl1_down_execute_lane0_logic_completions_onCtrl_1_ENABLE_lane0_5 = ((execute_lane0_logic_decoding_decodingBits & 33'h100002040) == 33'h100002040);
  always @(*) begin
    toplevel_execute_ctrl1_down_COMPLETION_AT_3_lane0 = _zz_toplevel_execute_ctrl1_down_COMPLETION_AT_3_lane0[0];
    if(toplevel_execute_ctrl1_down_TRAP_lane0) begin
      toplevel_execute_ctrl1_down_COMPLETION_AT_3_lane0 = 1'b0;
    end
  end

  assign _zz_toplevel_execute_ctrl1_down_execute_lane0_logic_completions_onCtrl_2_ENABLE_lane0_2 = ((execute_lane0_logic_decoding_decodingBits & 33'h002004064) == 33'h002000020);
  assign _zz_toplevel_execute_ctrl1_down_execute_lane0_logic_completions_onCtrl_2_ENABLE_lane0_3 = ((execute_lane0_logic_decoding_decodingBits & 33'h100000000) == 33'h0);
  always @(*) begin
    toplevel_execute_ctrl1_down_COMPLETION_AT_4_lane0 = _zz_toplevel_execute_ctrl1_down_COMPLETION_AT_4_lane0[0];
    if(toplevel_execute_ctrl1_down_TRAP_lane0) begin
      toplevel_execute_ctrl1_down_COMPLETION_AT_4_lane0 = 1'b0;
    end
  end

  always @(*) begin
    toplevel_execute_ctrl1_down_execute_lane0_logic_completions_onCtrl_0_ENABLE_lane0 = _zz_toplevel_execute_ctrl1_down_execute_lane0_logic_completions_onCtrl_0_ENABLE_lane0_7[0];
    if(toplevel_execute_ctrl1_down_TRAP_lane0) begin
      toplevel_execute_ctrl1_down_execute_lane0_logic_completions_onCtrl_0_ENABLE_lane0 = 1'b0;
    end
  end

  always @(*) begin
    toplevel_execute_ctrl1_down_execute_lane0_logic_completions_onCtrl_1_ENABLE_lane0 = _zz_toplevel_execute_ctrl1_down_execute_lane0_logic_completions_onCtrl_1_ENABLE_lane0_6[0];
    if(toplevel_execute_ctrl1_down_TRAP_lane0) begin
      toplevel_execute_ctrl1_down_execute_lane0_logic_completions_onCtrl_1_ENABLE_lane0 = 1'b0;
    end
  end

  always @(*) begin
    toplevel_execute_ctrl1_down_execute_lane0_logic_completions_onCtrl_2_ENABLE_lane0 = _zz_toplevel_execute_ctrl1_down_execute_lane0_logic_completions_onCtrl_2_ENABLE_lane0_4[0];
    if(toplevel_execute_ctrl1_down_TRAP_lane0) begin
      toplevel_execute_ctrl1_down_execute_lane0_logic_completions_onCtrl_2_ENABLE_lane0 = 1'b0;
    end
  end

  assign _zz_toplevel_execute_ctrl1_down_late0_IntAluPlugin_ALU_ADD_SUB_lane0 = ((execute_lane0_logic_decoding_decodingBits & 33'h000006000) == 33'h0);
  assign _zz_toplevel_execute_ctrl1_down_late0_SrcPlugin_logic_SRC2_CTRL_lane0 = ((execute_lane0_logic_decoding_decodingBits & 33'h000000004) == 33'h000000004);
  assign toplevel_execute_ctrl1_down_early0_IntAluPlugin_ALU_ADD_SUB_lane0 = _zz_toplevel_execute_ctrl1_down_early0_IntAluPlugin_ALU_ADD_SUB_lane0[0];
  assign _zz_toplevel_execute_ctrl1_down_late0_IntAluPlugin_ALU_SLTX_lane0 = ((execute_lane0_logic_decoding_decodingBits & 33'h000006004) == 33'h000002000);
  assign toplevel_execute_ctrl1_down_early0_IntAluPlugin_ALU_SLTX_lane0 = _zz_toplevel_execute_ctrl1_down_early0_IntAluPlugin_ALU_SLTX_lane0[0];
  assign _zz_toplevel_execute_ctrl1_down_late0_IntAluPlugin_ALU_BITWISE_CTRL_lane0 = ((execute_lane0_logic_decoding_decodingBits & 33'h000003000) == 33'h000002000);
  assign _zz_toplevel_execute_ctrl1_down_BarrelShifterPlugin_LEFT_lane0 = ((execute_lane0_logic_decoding_decodingBits & 33'h000004000) == 33'h0);
  assign _zz_toplevel_execute_ctrl1_down_CsrAccessPlugin_CSR_CLEAR_lane0 = ((execute_lane0_logic_decoding_decodingBits & 33'h000001000) == 33'h000001000);
  assign _zz_toplevel_execute_ctrl1_down_early0_IntAluPlugin_ALU_BITWISE_CTRL_lane0_1 = {(|{_zz_toplevel_execute_ctrl1_down_CsrAccessPlugin_CSR_CLEAR_lane0,{_zz_toplevel_execute_ctrl1_down_late0_SrcPlugin_logic_SRC2_CTRL_lane0,_zz_toplevel_execute_ctrl1_down_BarrelShifterPlugin_LEFT_lane0}}),(|{_zz_toplevel_execute_ctrl1_down_late0_SrcPlugin_logic_SRC2_CTRL_lane0,{_zz_toplevel_execute_ctrl1_down_BarrelShifterPlugin_LEFT_lane0,_zz_toplevel_execute_ctrl1_down_late0_IntAluPlugin_ALU_BITWISE_CTRL_lane0}})};
  assign _zz_toplevel_execute_ctrl1_down_early0_IntAluPlugin_ALU_BITWISE_CTRL_lane0 = _zz_toplevel_execute_ctrl1_down_early0_IntAluPlugin_ALU_BITWISE_CTRL_lane0_1;
  assign _zz_toplevel_execute_ctrl1_down_early0_IntAluPlugin_ALU_BITWISE_CTRL_lane0_2 = _zz_toplevel_execute_ctrl1_down_early0_IntAluPlugin_ALU_BITWISE_CTRL_lane0;
  assign toplevel_execute_ctrl1_down_early0_IntAluPlugin_ALU_BITWISE_CTRL_lane0 = _zz_toplevel_execute_ctrl1_down_early0_IntAluPlugin_ALU_BITWISE_CTRL_lane0_2;
  assign toplevel_execute_ctrl1_down_SrcStageables_REVERT_lane0 = _zz_toplevel_execute_ctrl1_down_SrcStageables_REVERT_lane0[0];
  assign toplevel_execute_ctrl1_down_SrcStageables_ZERO_lane0 = _zz_toplevel_execute_ctrl1_down_SrcStageables_ZERO_lane0[0];
  assign toplevel_execute_ctrl1_down_early0_SrcPlugin_logic_SRC1_CTRL_lane0 = (|((execute_lane0_logic_decoding_decodingBits & 33'h00000004c) == 33'h000000004));
  assign _zz_toplevel_execute_ctrl1_down_late0_SrcPlugin_logic_SRC2_CTRL_lane0_1 = ((execute_lane0_logic_decoding_decodingBits & 33'h000000024) == 33'h0);
  assign toplevel_execute_ctrl1_down_early0_SrcPlugin_logic_SRC2_CTRL_lane0 = {(|{_zz_toplevel_execute_ctrl1_down_late0_SrcPlugin_logic_SRC2_CTRL_lane0,((execute_lane0_logic_decoding_decodingBits & 33'h000000070) == 33'h000000020)}),(|{((execute_lane0_logic_decoding_decodingBits & 33'h000000050) == 33'h0),_zz_toplevel_execute_ctrl1_down_late0_SrcPlugin_logic_SRC2_CTRL_lane0_1})};
  assign toplevel_execute_ctrl1_down_lane0_IntFormatPlugin_logic_SIGNED_lane0 = _zz_toplevel_execute_ctrl1_down_lane0_IntFormatPlugin_logic_SIGNED_lane0[0];
  assign _zz_toplevel_execute_ctrl1_down_AguPlugin_STORE_lane0 = ((execute_lane0_logic_decoding_decodingBits & 33'h010000020) == 33'h000000020);
  assign toplevel_execute_ctrl1_down_lane0_IntFormatPlugin_logic_WIDTH_ID_lane0 = {(|{((execute_lane0_logic_decoding_decodingBits & 33'h000000010) == 33'h000000010),{((execute_lane0_logic_decoding_decodingBits & _zz_toplevel_execute_ctrl1_down_lane0_IntFormatPlugin_logic_WIDTH_ID_lane0) == 33'h000002000),{_zz_toplevel_execute_ctrl1_down_AguPlugin_STORE_lane0,(_zz_toplevel_execute_ctrl1_down_lane0_IntFormatPlugin_logic_WIDTH_ID_lane0_1 == _zz_toplevel_execute_ctrl1_down_lane0_IntFormatPlugin_logic_WIDTH_ID_lane0_2)}}}),(|((execute_lane0_logic_decoding_decodingBits & 33'h000001010) == 33'h000001000))};
  assign _zz_toplevel_execute_ctrl1_down_BYPASSED_AT_3_lane0 = ((execute_lane0_logic_decoding_decodingBits & 33'h10000000c) == 33'h100000004);
  assign toplevel_execute_ctrl1_down_BYPASSED_AT_2_lane0 = _zz_toplevel_execute_ctrl1_down_BYPASSED_AT_2_lane0[0];
  assign toplevel_execute_ctrl1_down_BYPASSED_AT_3_lane0 = _zz_toplevel_execute_ctrl1_down_BYPASSED_AT_3_lane0_1[0];
  assign _zz_toplevel_execute_ctrl1_down_SrcStageables_UNSIGNED_lane0 = ((execute_lane0_logic_decoding_decodingBits & 33'h000002010) == 33'h000002000);
  assign toplevel_execute_ctrl1_down_MAY_FLUSH_PRECISE_3_lane0 = _zz_toplevel_execute_ctrl1_down_MAY_FLUSH_PRECISE_3_lane0[0];
  assign toplevel_execute_ctrl1_down_MAY_FLUSH_PRECISE_4_lane0 = _zz_toplevel_execute_ctrl1_down_MAY_FLUSH_PRECISE_4_lane0[0];
  assign toplevel_execute_ctrl1_down_SrcStageables_UNSIGNED_lane0 = _zz_toplevel_execute_ctrl1_down_SrcStageables_UNSIGNED_lane0_1[0];
  assign toplevel_execute_ctrl1_down_BarrelShifterPlugin_LEFT_lane0 = _zz_toplevel_execute_ctrl1_down_BarrelShifterPlugin_LEFT_lane0_1[0];
  assign toplevel_execute_ctrl1_down_BarrelShifterPlugin_SIGNED_lane0 = _zz_toplevel_execute_ctrl1_down_BarrelShifterPlugin_SIGNED_lane0[0];
  assign _zz_toplevel_execute_ctrl1_down_BranchPlugin_BRANCH_CTRL_lane0_1 = {(|_zz_toplevel_execute_ctrl1_down_lane0_integer_WriteBackPlugin_SEL_lane0),(|((execute_lane0_logic_decoding_decodingBits & 33'h000000008) == 33'h000000008))};
  assign _zz_toplevel_execute_ctrl1_down_BranchPlugin_BRANCH_CTRL_lane0 = _zz_toplevel_execute_ctrl1_down_BranchPlugin_BRANCH_CTRL_lane0_1;
  assign _zz_toplevel_execute_ctrl1_down_BranchPlugin_BRANCH_CTRL_lane0_2 = _zz_toplevel_execute_ctrl1_down_BranchPlugin_BRANCH_CTRL_lane0;
  assign toplevel_execute_ctrl1_down_BranchPlugin_BRANCH_CTRL_lane0 = _zz_toplevel_execute_ctrl1_down_BranchPlugin_BRANCH_CTRL_lane0_2;
  assign toplevel_execute_ctrl1_down_RsUnsignedPlugin_RS1_SIGNED_lane0 = _zz_toplevel_execute_ctrl1_down_RsUnsignedPlugin_RS1_SIGNED_lane0[0];
  assign toplevel_execute_ctrl1_down_RsUnsignedPlugin_RS2_SIGNED_lane0 = _zz_toplevel_execute_ctrl1_down_RsUnsignedPlugin_RS2_SIGNED_lane0[0];
  assign _zz_toplevel_execute_ctrl1_down_CsrAccessPlugin_CSR_MASK_lane0 = ((execute_lane0_logic_decoding_decodingBits & 33'h000002000) == 33'h000002000);
  assign toplevel_execute_ctrl1_down_DivPlugin_REM_lane0 = _zz_toplevel_execute_ctrl1_down_DivPlugin_REM_lane0[0];
  assign toplevel_execute_ctrl1_down_CsrAccessPlugin_CSR_IMM_lane0 = _zz_toplevel_execute_ctrl1_down_CsrAccessPlugin_CSR_IMM_lane0[0];
  assign toplevel_execute_ctrl1_down_CsrAccessPlugin_CSR_MASK_lane0 = _zz_toplevel_execute_ctrl1_down_CsrAccessPlugin_CSR_MASK_lane0_1[0];
  assign toplevel_execute_ctrl1_down_CsrAccessPlugin_CSR_CLEAR_lane0 = _zz_toplevel_execute_ctrl1_down_CsrAccessPlugin_CSR_CLEAR_lane0_1[0];
  assign toplevel_execute_ctrl1_down_AguPlugin_LOAD_lane0 = _zz_toplevel_execute_ctrl1_down_AguPlugin_LOAD_lane0_1[0];
  assign toplevel_execute_ctrl1_down_AguPlugin_STORE_lane0 = _zz_toplevel_execute_ctrl1_down_AguPlugin_STORE_lane0_1[0];
  assign toplevel_execute_ctrl1_down_AguPlugin_ATOMIC_lane0 = _zz_toplevel_execute_ctrl1_down_AguPlugin_ATOMIC_lane0_1[0];
  assign toplevel_execute_ctrl1_down_AguPlugin_FLOAT_lane0 = _zz_toplevel_execute_ctrl1_down_AguPlugin_FLOAT_lane0[0];
  assign toplevel_execute_ctrl1_down_LsuPlugin_logic_LSU_PREFETCH_lane0 = _zz_toplevel_execute_ctrl1_down_LsuPlugin_logic_LSU_PREFETCH_lane0[0];
  assign _zz_toplevel_execute_ctrl1_down_early0_EnvPlugin_OP_lane0 = ((execute_lane0_logic_decoding_decodingBits & 33'h000000040) == 33'h0);
  assign _zz_toplevel_execute_ctrl1_down_early0_EnvPlugin_OP_lane0_2 = {(|{((execute_lane0_logic_decoding_decodingBits & _zz__zz_toplevel_execute_ctrl1_down_early0_EnvPlugin_OP_lane0_2) == 33'h002000000),((execute_lane0_logic_decoding_decodingBits & _zz__zz_toplevel_execute_ctrl1_down_early0_EnvPlugin_OP_lane0_2_1) == 33'h010000000)}),{(|{_zz_toplevel_execute_ctrl1_down_early0_EnvPlugin_OP_lane0,(_zz__zz_toplevel_execute_ctrl1_down_early0_EnvPlugin_OP_lane0_2_2 == _zz__zz_toplevel_execute_ctrl1_down_early0_EnvPlugin_OP_lane0_2_3)}),(|{_zz_toplevel_execute_ctrl1_down_early0_EnvPlugin_OP_lane0,{_zz__zz_toplevel_execute_ctrl1_down_early0_EnvPlugin_OP_lane0_2_4,_zz__zz_toplevel_execute_ctrl1_down_early0_EnvPlugin_OP_lane0_2_5}})}};
  assign _zz_toplevel_execute_ctrl1_down_early0_EnvPlugin_OP_lane0_1 = _zz_toplevel_execute_ctrl1_down_early0_EnvPlugin_OP_lane0_2;
  assign _zz_toplevel_execute_ctrl1_down_early0_EnvPlugin_OP_lane0_3 = _zz_toplevel_execute_ctrl1_down_early0_EnvPlugin_OP_lane0_1;
  assign toplevel_execute_ctrl1_down_early0_EnvPlugin_OP_lane0 = _zz_toplevel_execute_ctrl1_down_early0_EnvPlugin_OP_lane0_3;
  assign toplevel_execute_ctrl1_down_late0_IntAluPlugin_ALU_ADD_SUB_lane0 = _zz_toplevel_execute_ctrl1_down_late0_IntAluPlugin_ALU_ADD_SUB_lane0_1[0];
  assign toplevel_execute_ctrl1_down_late0_IntAluPlugin_ALU_SLTX_lane0 = _zz_toplevel_execute_ctrl1_down_late0_IntAluPlugin_ALU_SLTX_lane0_1[0];
  assign _zz_toplevel_execute_ctrl1_down_late0_IntAluPlugin_ALU_BITWISE_CTRL_lane0_2 = {(|{_zz_toplevel_execute_ctrl1_down_CsrAccessPlugin_CSR_CLEAR_lane0,{_zz_toplevel_execute_ctrl1_down_late0_SrcPlugin_logic_SRC2_CTRL_lane0,_zz_toplevel_execute_ctrl1_down_BarrelShifterPlugin_LEFT_lane0}}),(|{_zz_toplevel_execute_ctrl1_down_late0_SrcPlugin_logic_SRC2_CTRL_lane0,{_zz_toplevel_execute_ctrl1_down_BarrelShifterPlugin_LEFT_lane0,_zz_toplevel_execute_ctrl1_down_late0_IntAluPlugin_ALU_BITWISE_CTRL_lane0}})};
  assign _zz_toplevel_execute_ctrl1_down_late0_IntAluPlugin_ALU_BITWISE_CTRL_lane0_1 = _zz_toplevel_execute_ctrl1_down_late0_IntAluPlugin_ALU_BITWISE_CTRL_lane0_2;
  assign _zz_toplevel_execute_ctrl1_down_late0_IntAluPlugin_ALU_BITWISE_CTRL_lane0_3 = _zz_toplevel_execute_ctrl1_down_late0_IntAluPlugin_ALU_BITWISE_CTRL_lane0_1;
  assign toplevel_execute_ctrl1_down_late0_IntAluPlugin_ALU_BITWISE_CTRL_lane0 = _zz_toplevel_execute_ctrl1_down_late0_IntAluPlugin_ALU_BITWISE_CTRL_lane0_3;
  assign toplevel_execute_ctrl1_down_late0_SrcPlugin_logic_SRC1_CTRL_lane0 = (|_zz_toplevel_execute_ctrl1_down_late0_SrcPlugin_logic_SRC2_CTRL_lane0);
  assign toplevel_execute_ctrl1_down_late0_SrcPlugin_logic_SRC2_CTRL_lane0 = {(|_zz_toplevel_execute_ctrl1_down_late0_SrcPlugin_logic_SRC2_CTRL_lane0),(|_zz_toplevel_execute_ctrl1_down_late0_SrcPlugin_logic_SRC2_CTRL_lane0_1)};
  assign when_ExecuteLanePlugin_l300 = (|{(late1_BranchPlugin_logic_flushPort_valid && 1'b1),{(early1_BranchPlugin_logic_flushPort_valid && 1'b1),{(late0_BranchPlugin_logic_flushPort_valid && 1'b1),{(early0_EnvPlugin_logic_flushPort_valid && 1'b1),{(CsrAccessPlugin_logic_flushPort_valid && 1'b1),{(early0_BranchPlugin_logic_flushPort_valid && 1'b1),(LsuPlugin_logic_flushPort_valid && 1'b1)}}}}}});
  assign toplevel_execute_lane0_ctrls_0_downIsCancel = 1'b0;
  assign toplevel_execute_lane0_ctrls_0_upIsCancel = when_ExecuteLanePlugin_l300;
  assign when_ExecuteLanePlugin_l300_1 = (|{(late1_BranchPlugin_logic_flushPort_valid && 1'b1),{(early1_BranchPlugin_logic_flushPort_valid && 1'b1),{(late0_BranchPlugin_logic_flushPort_valid && 1'b1),{(early0_EnvPlugin_logic_flushPort_valid && 1'b1),{(CsrAccessPlugin_logic_flushPort_valid && 1'b1),{(early0_BranchPlugin_logic_flushPort_valid && 1'b1),(LsuPlugin_logic_flushPort_valid && 1'b1)}}}}}});
  assign toplevel_execute_lane0_ctrls_1_downIsCancel = 1'b0;
  assign toplevel_execute_lane0_ctrls_1_upIsCancel = when_ExecuteLanePlugin_l300_1;
  assign when_ExecuteLanePlugin_l300_2 = (|{(late1_BranchPlugin_logic_flushPort_valid && 1'b1),{(early1_BranchPlugin_logic_flushPort_valid && 1'b1),{(late0_BranchPlugin_logic_flushPort_valid && 1'b1),{((early0_EnvPlugin_logic_flushPort_valid && 1'b1) && ((early0_EnvPlugin_logic_flushPort_payload_laneAge < toplevel_execute_ctrl2_down_LANE_AGE_lane0) || (_zz_when_ExecuteLanePlugin_l300_2 && early0_EnvPlugin_logic_flushPort_payload_self))),{((CsrAccessPlugin_logic_flushPort_valid && _zz_when_ExecuteLanePlugin_l300_2_1) && (_zz_when_ExecuteLanePlugin_l300_2_2 || _zz_when_ExecuteLanePlugin_l300_2_3)),{(early0_BranchPlugin_logic_flushPort_valid && _zz_when_ExecuteLanePlugin_l300_2_4),(LsuPlugin_logic_flushPort_valid && _zz_when_ExecuteLanePlugin_l300_2_5)}}}}}});
  assign toplevel_execute_lane0_ctrls_2_downIsCancel = 1'b0;
  assign toplevel_execute_lane0_ctrls_2_upIsCancel = when_ExecuteLanePlugin_l300_2;
  assign when_ExecuteLanePlugin_l300_3 = (|{(late1_BranchPlugin_logic_flushPort_valid && 1'b1),{((early1_BranchPlugin_logic_flushPort_valid && 1'b1) && ((early1_BranchPlugin_logic_flushPort_payload_laneAge < toplevel_execute_ctrl3_down_LANE_AGE_lane0) || ((early1_BranchPlugin_logic_flushPort_payload_laneAge == toplevel_execute_ctrl3_down_LANE_AGE_lane0) && early1_BranchPlugin_logic_flushPort_payload_self))),{(late0_BranchPlugin_logic_flushPort_valid && 1'b1),{((early0_BranchPlugin_logic_flushPort_valid && _zz_when_ExecuteLanePlugin_l300_3) && (_zz_when_ExecuteLanePlugin_l300_3_1 || _zz_when_ExecuteLanePlugin_l300_3_2)),(LsuPlugin_logic_flushPort_valid && 1'b1)}}}});
  assign toplevel_execute_lane0_ctrls_3_downIsCancel = 1'b0;
  assign toplevel_execute_lane0_ctrls_3_upIsCancel = when_ExecuteLanePlugin_l300_3;
  assign when_ExecuteLanePlugin_l300_4 = (|{((late1_BranchPlugin_logic_flushPort_valid && 1'b1) && ((late1_BranchPlugin_logic_flushPort_payload_laneAge < toplevel_execute_ctrl4_down_LANE_AGE_lane0) || ((late1_BranchPlugin_logic_flushPort_payload_laneAge == toplevel_execute_ctrl4_down_LANE_AGE_lane0) && late1_BranchPlugin_logic_flushPort_payload_self))),{((late0_BranchPlugin_logic_flushPort_valid && 1'b1) && ((late0_BranchPlugin_logic_flushPort_payload_laneAge < toplevel_execute_ctrl4_down_LANE_AGE_lane0) || (_zz_when_ExecuteLanePlugin_l300_4 && late0_BranchPlugin_logic_flushPort_payload_self))),((LsuPlugin_logic_flushPort_valid && 1'b1) && ((LsuPlugin_logic_flushPort_payload_laneAge < toplevel_execute_ctrl4_down_LANE_AGE_lane0) || (_zz_when_ExecuteLanePlugin_l300_4_1 && LsuPlugin_logic_flushPort_payload_self)))}});
  assign toplevel_execute_lane0_ctrls_4_downIsCancel = 1'b0;
  assign toplevel_execute_lane0_ctrls_4_upIsCancel = when_ExecuteLanePlugin_l300_4;
  assign toplevel_execute_lane0_ctrls_5_downIsCancel = 1'b0;
  assign toplevel_execute_lane0_ctrls_5_upIsCancel = 1'b0;
  assign execute_lane0_logic_trapPending[0] = (|{((toplevel_execute_ctrl4_up_LANE_SEL_lane0 && 1'b1) && toplevel_execute_ctrl4_down_TRAP_lane0),{((toplevel_execute_ctrl3_up_LANE_SEL_lane0 && 1'b1) && toplevel_execute_ctrl3_down_TRAP_lane0),{((toplevel_execute_ctrl2_up_LANE_SEL_lane0 && 1'b1) && toplevel_execute_ctrl2_down_TRAP_lane0),((toplevel_execute_ctrl1_up_LANE_SEL_lane0 && 1'b1) && toplevel_execute_ctrl1_down_TRAP_lane0)}}});
  assign toplevel_execute_ctrl2_up_COMMIT_lane0 = (! toplevel_execute_ctrl2_up_TRAP_lane0);
  assign WhiteboxerPlugin_logic_csr_access_valid = CsrAccessPlugin_logic_fsm_regs_fire;
  assign WhiteboxerPlugin_logic_csr_access_payload_uopId = CsrAccessPlugin_logic_fsm_regs_uopId;
  assign WhiteboxerPlugin_logic_csr_access_payload_address = _zz_WhiteboxerPlugin_logic_csr_access_payload_address[31 : 20];
  assign WhiteboxerPlugin_logic_csr_access_payload_write = CsrAccessPlugin_logic_fsm_regs_onWriteBits;
  assign WhiteboxerPlugin_logic_csr_access_payload_read = CsrAccessPlugin_logic_fsm_regs_csrValue;
  assign WhiteboxerPlugin_logic_csr_access_payload_writeDone = CsrAccessPlugin_logic_fsm_regs_write;
  assign WhiteboxerPlugin_logic_csr_access_payload_readDone = CsrAccessPlugin_logic_fsm_regs_read;
  assign WhiteboxerPlugin_logic_csr_port_valid = WhiteboxerPlugin_logic_csr_access_valid;
  assign WhiteboxerPlugin_logic_csr_port_payload_uopId = WhiteboxerPlugin_logic_csr_access_payload_uopId;
  assign WhiteboxerPlugin_logic_csr_port_payload_address = WhiteboxerPlugin_logic_csr_access_payload_address;
  assign WhiteboxerPlugin_logic_csr_port_payload_write = WhiteboxerPlugin_logic_csr_access_payload_write;
  assign WhiteboxerPlugin_logic_csr_port_payload_read = WhiteboxerPlugin_logic_csr_access_payload_read;
  assign WhiteboxerPlugin_logic_csr_port_payload_writeDone = WhiteboxerPlugin_logic_csr_access_payload_writeDone;
  assign WhiteboxerPlugin_logic_csr_port_payload_readDone = WhiteboxerPlugin_logic_csr_access_payload_readDone;
  assign WhiteboxerPlugin_logic_rfWrites_ports_0_valid = lane0_integer_WriteBackPlugin_logic_stages_0_write_valid;
  assign WhiteboxerPlugin_logic_rfWrites_ports_0_payload_uopId = lane0_integer_WriteBackPlugin_logic_stages_0_write_payload_uopId;
  assign WhiteboxerPlugin_logic_rfWrites_ports_0_payload_data = lane0_integer_WriteBackPlugin_logic_stages_0_write_payload_data;
  assign WhiteboxerPlugin_logic_rfWrites_ports_1_valid = lane0_integer_WriteBackPlugin_logic_stages_1_write_valid;
  assign WhiteboxerPlugin_logic_rfWrites_ports_1_payload_uopId = lane0_integer_WriteBackPlugin_logic_stages_1_write_payload_uopId;
  assign WhiteboxerPlugin_logic_rfWrites_ports_1_payload_data = lane0_integer_WriteBackPlugin_logic_stages_1_write_payload_data;
  assign WhiteboxerPlugin_logic_rfWrites_ports_2_valid = lane0_integer_WriteBackPlugin_logic_stages_2_write_valid;
  assign WhiteboxerPlugin_logic_rfWrites_ports_2_payload_uopId = lane0_integer_WriteBackPlugin_logic_stages_2_write_payload_uopId;
  assign WhiteboxerPlugin_logic_rfWrites_ports_2_payload_data = lane0_integer_WriteBackPlugin_logic_stages_2_write_payload_data;
  assign WhiteboxerPlugin_logic_rfWrites_ports_3_valid = lane1_integer_WriteBackPlugin_logic_stages_0_write_valid;
  assign WhiteboxerPlugin_logic_rfWrites_ports_3_payload_uopId = lane1_integer_WriteBackPlugin_logic_stages_0_write_payload_uopId;
  assign WhiteboxerPlugin_logic_rfWrites_ports_3_payload_data = lane1_integer_WriteBackPlugin_logic_stages_0_write_payload_data;
  assign WhiteboxerPlugin_logic_rfWrites_ports_4_valid = lane1_integer_WriteBackPlugin_logic_stages_1_write_valid;
  assign WhiteboxerPlugin_logic_rfWrites_ports_4_payload_uopId = lane1_integer_WriteBackPlugin_logic_stages_1_write_payload_uopId;
  assign WhiteboxerPlugin_logic_rfWrites_ports_4_payload_data = lane1_integer_WriteBackPlugin_logic_stages_1_write_payload_data;
  assign WhiteboxerPlugin_logic_rfWrites_ports_5_valid = lane1_integer_WriteBackPlugin_logic_stages_2_write_valid;
  assign WhiteboxerPlugin_logic_rfWrites_ports_5_payload_uopId = lane1_integer_WriteBackPlugin_logic_stages_2_write_payload_uopId;
  assign WhiteboxerPlugin_logic_rfWrites_ports_5_payload_data = lane1_integer_WriteBackPlugin_logic_stages_2_write_payload_data;
  assign WhiteboxerPlugin_logic_completions_ports_0_valid = DecoderPlugin_logic_laneLogic_0_completionPort_valid;
  assign WhiteboxerPlugin_logic_completions_ports_0_payload_uopId = DecoderPlugin_logic_laneLogic_0_completionPort_payload_uopId;
  assign WhiteboxerPlugin_logic_completions_ports_0_payload_trap = DecoderPlugin_logic_laneLogic_0_completionPort_payload_trap;
  assign WhiteboxerPlugin_logic_completions_ports_0_payload_commit = DecoderPlugin_logic_laneLogic_0_completionPort_payload_commit;
  assign WhiteboxerPlugin_logic_completions_ports_1_valid = DecoderPlugin_logic_laneLogic_1_completionPort_valid;
  assign WhiteboxerPlugin_logic_completions_ports_1_payload_uopId = DecoderPlugin_logic_laneLogic_1_completionPort_payload_uopId;
  assign WhiteboxerPlugin_logic_completions_ports_1_payload_trap = DecoderPlugin_logic_laneLogic_1_completionPort_payload_trap;
  assign WhiteboxerPlugin_logic_completions_ports_1_payload_commit = DecoderPlugin_logic_laneLogic_1_completionPort_payload_commit;
  assign WhiteboxerPlugin_logic_completions_ports_2_valid = execute_lane0_logic_completions_onCtrl_0_port_valid;
  assign WhiteboxerPlugin_logic_completions_ports_2_payload_uopId = execute_lane0_logic_completions_onCtrl_0_port_payload_uopId;
  assign WhiteboxerPlugin_logic_completions_ports_2_payload_trap = execute_lane0_logic_completions_onCtrl_0_port_payload_trap;
  assign WhiteboxerPlugin_logic_completions_ports_2_payload_commit = execute_lane0_logic_completions_onCtrl_0_port_payload_commit;
  assign WhiteboxerPlugin_logic_completions_ports_3_valid = execute_lane0_logic_completions_onCtrl_1_port_valid;
  assign WhiteboxerPlugin_logic_completions_ports_3_payload_uopId = execute_lane0_logic_completions_onCtrl_1_port_payload_uopId;
  assign WhiteboxerPlugin_logic_completions_ports_3_payload_trap = execute_lane0_logic_completions_onCtrl_1_port_payload_trap;
  assign WhiteboxerPlugin_logic_completions_ports_3_payload_commit = execute_lane0_logic_completions_onCtrl_1_port_payload_commit;
  assign WhiteboxerPlugin_logic_completions_ports_4_valid = execute_lane0_logic_completions_onCtrl_2_port_valid;
  assign WhiteboxerPlugin_logic_completions_ports_4_payload_uopId = execute_lane0_logic_completions_onCtrl_2_port_payload_uopId;
  assign WhiteboxerPlugin_logic_completions_ports_4_payload_trap = execute_lane0_logic_completions_onCtrl_2_port_payload_trap;
  assign WhiteboxerPlugin_logic_completions_ports_4_payload_commit = execute_lane0_logic_completions_onCtrl_2_port_payload_commit;
  assign fetch_logic_flushes_0_doIt = (|{(DecoderPlugin_logic_laneLogic_1_flushPort_valid && 1'b1),{(DecoderPlugin_logic_laneLogic_0_flushPort_valid && 1'b1),{(late1_BranchPlugin_logic_flushPort_valid && 1'b1),{(early1_BranchPlugin_logic_flushPort_valid && 1'b1),{(late0_BranchPlugin_logic_flushPort_valid && 1'b1),{(early0_EnvPlugin_logic_flushPort_valid && _zz_fetch_logic_flushes_0_doIt),{_zz_fetch_logic_flushes_0_doIt_1,{_zz_fetch_logic_flushes_0_doIt_2,_zz_fetch_logic_flushes_0_doIt_3}}}}}}}});
  assign fetch_logic_ctrls_1_throwWhen_FetchPipelinePlugin_l44 = fetch_logic_flushes_0_doIt;
  assign fetch_logic_flushes_1_doIt = (|{(DecoderPlugin_logic_laneLogic_1_flushPort_valid && 1'b1),{(DecoderPlugin_logic_laneLogic_0_flushPort_valid && 1'b1),{(late1_BranchPlugin_logic_flushPort_valid && 1'b1),{(early1_BranchPlugin_logic_flushPort_valid && 1'b1),{(late0_BranchPlugin_logic_flushPort_valid && 1'b1),{(early0_EnvPlugin_logic_flushPort_valid && _zz_fetch_logic_flushes_1_doIt),{_zz_fetch_logic_flushes_1_doIt_1,{_zz_fetch_logic_flushes_1_doIt_2,_zz_fetch_logic_flushes_1_doIt_3}}}}}}}});
  assign fetch_logic_ctrls_2_forgetsSingleRequest_FetchPipelinePlugin_l46 = fetch_logic_flushes_1_doIt;
  always @(*) begin
    toplevel_execute_lane1_bypasser_integer_RS1_bypassEnables[0] = (((toplevel_execute_ctrl2_up_LANE_SEL_lane0 && toplevel_execute_ctrl2_up_RD_ENABLE_lane0) && (toplevel_execute_ctrl2_down_RD_PHYS_lane0 == toplevel_execute_ctrl1_down_RS1_PHYS_lane1)) && 1'b1);
    toplevel_execute_lane1_bypasser_integer_RS1_bypassEnables[1] = (((toplevel_execute_ctrl2_up_LANE_SEL_lane1 && toplevel_execute_ctrl2_up_RD_ENABLE_lane1) && (toplevel_execute_ctrl2_down_RD_PHYS_lane1 == toplevel_execute_ctrl1_down_RS1_PHYS_lane1)) && 1'b1);
    toplevel_execute_lane1_bypasser_integer_RS1_bypassEnables[2] = (((toplevel_execute_ctrl3_up_LANE_SEL_lane0 && toplevel_execute_ctrl3_up_RD_ENABLE_lane0) && (toplevel_execute_ctrl3_down_RD_PHYS_lane0 == toplevel_execute_ctrl1_down_RS1_PHYS_lane1)) && 1'b1);
    toplevel_execute_lane1_bypasser_integer_RS1_bypassEnables[3] = (((toplevel_execute_ctrl3_up_LANE_SEL_lane1 && toplevel_execute_ctrl3_up_RD_ENABLE_lane1) && (toplevel_execute_ctrl3_down_RD_PHYS_lane1 == toplevel_execute_ctrl1_down_RS1_PHYS_lane1)) && 1'b1);
    toplevel_execute_lane1_bypasser_integer_RS1_bypassEnables[4] = (((toplevel_execute_ctrl4_up_LANE_SEL_lane0 && toplevel_execute_ctrl4_up_RD_ENABLE_lane0) && (toplevel_execute_ctrl4_down_RD_PHYS_lane0 == toplevel_execute_ctrl1_down_RS1_PHYS_lane1)) && 1'b1);
    toplevel_execute_lane1_bypasser_integer_RS1_bypassEnables[5] = (((toplevel_execute_ctrl4_up_LANE_SEL_lane1 && toplevel_execute_ctrl4_up_RD_ENABLE_lane1) && (toplevel_execute_ctrl4_down_RD_PHYS_lane1 == toplevel_execute_ctrl1_down_RS1_PHYS_lane1)) && 1'b1);
    toplevel_execute_lane1_bypasser_integer_RS1_bypassEnables[6] = (((toplevel_execute_ctrl5_up_LANE_SEL_lane0 && toplevel_execute_ctrl5_up_RD_ENABLE_lane0) && (toplevel_execute_ctrl5_down_RD_PHYS_lane0 == toplevel_execute_ctrl1_down_RS1_PHYS_lane1)) && 1'b1);
    toplevel_execute_lane1_bypasser_integer_RS1_bypassEnables[7] = (((toplevel_execute_ctrl5_up_LANE_SEL_lane1 && toplevel_execute_ctrl5_up_RD_ENABLE_lane1) && (toplevel_execute_ctrl5_down_RD_PHYS_lane1 == toplevel_execute_ctrl1_down_RS1_PHYS_lane1)) && 1'b1);
    toplevel_execute_lane1_bypasser_integer_RS1_bypassEnables[8] = 1'b1;
  end

  assign _zz_toplevel_execute_lane1_bypasser_integer_RS1_bypassEnables_bools_0 = toplevel_execute_lane1_bypasser_integer_RS1_bypassEnables;
  assign toplevel_execute_lane1_bypasser_integer_RS1_bypassEnables_bools_0 = _zz_toplevel_execute_lane1_bypasser_integer_RS1_bypassEnables_bools_0[0];
  assign toplevel_execute_lane1_bypasser_integer_RS1_bypassEnables_bools_1 = _zz_toplevel_execute_lane1_bypasser_integer_RS1_bypassEnables_bools_0[1];
  assign toplevel_execute_lane1_bypasser_integer_RS1_bypassEnables_bools_2 = _zz_toplevel_execute_lane1_bypasser_integer_RS1_bypassEnables_bools_0[2];
  assign toplevel_execute_lane1_bypasser_integer_RS1_bypassEnables_bools_3 = _zz_toplevel_execute_lane1_bypasser_integer_RS1_bypassEnables_bools_0[3];
  assign toplevel_execute_lane1_bypasser_integer_RS1_bypassEnables_bools_4 = _zz_toplevel_execute_lane1_bypasser_integer_RS1_bypassEnables_bools_0[4];
  assign toplevel_execute_lane1_bypasser_integer_RS1_bypassEnables_bools_5 = _zz_toplevel_execute_lane1_bypasser_integer_RS1_bypassEnables_bools_0[5];
  assign toplevel_execute_lane1_bypasser_integer_RS1_bypassEnables_bools_6 = _zz_toplevel_execute_lane1_bypasser_integer_RS1_bypassEnables_bools_0[6];
  assign toplevel_execute_lane1_bypasser_integer_RS1_bypassEnables_bools_7 = _zz_toplevel_execute_lane1_bypasser_integer_RS1_bypassEnables_bools_0[7];
  assign toplevel_execute_lane1_bypasser_integer_RS1_bypassEnables_bools_8 = _zz_toplevel_execute_lane1_bypasser_integer_RS1_bypassEnables_bools_0[8];
  always @(*) begin
    _zz_toplevel_execute_lane1_bypasser_integer_RS1_sel[0] = (toplevel_execute_lane1_bypasser_integer_RS1_bypassEnables_bools_0 && (! 1'b0));
    _zz_toplevel_execute_lane1_bypasser_integer_RS1_sel[1] = (toplevel_execute_lane1_bypasser_integer_RS1_bypassEnables_bools_1 && (! toplevel_execute_lane1_bypasser_integer_RS1_bypassEnables_bools_0));
    _zz_toplevel_execute_lane1_bypasser_integer_RS1_sel[2] = (toplevel_execute_lane1_bypasser_integer_RS1_bypassEnables_bools_2 && (! toplevel_execute_lane1_bypasser_integer_RS1_bypassEnables_range_0_to_1));
    _zz_toplevel_execute_lane1_bypasser_integer_RS1_sel[3] = (toplevel_execute_lane1_bypasser_integer_RS1_bypassEnables_bools_3 && (! toplevel_execute_lane1_bypasser_integer_RS1_bypassEnables_range_0_to_2));
    _zz_toplevel_execute_lane1_bypasser_integer_RS1_sel[4] = (toplevel_execute_lane1_bypasser_integer_RS1_bypassEnables_bools_4 && (! toplevel_execute_lane1_bypasser_integer_RS1_bypassEnables_range_0_to_3));
    _zz_toplevel_execute_lane1_bypasser_integer_RS1_sel[5] = (toplevel_execute_lane1_bypasser_integer_RS1_bypassEnables_bools_5 && (! (toplevel_execute_lane1_bypasser_integer_RS1_bypassEnables_bools_4 || toplevel_execute_lane1_bypasser_integer_RS1_bypassEnables_range_0_to_3)));
    _zz_toplevel_execute_lane1_bypasser_integer_RS1_sel[6] = (toplevel_execute_lane1_bypasser_integer_RS1_bypassEnables_bools_6 && (! (toplevel_execute_lane1_bypasser_integer_RS1_bypassEnables_range_4_to_5 || toplevel_execute_lane1_bypasser_integer_RS1_bypassEnables_range_0_to_3)));
    _zz_toplevel_execute_lane1_bypasser_integer_RS1_sel[7] = (toplevel_execute_lane1_bypasser_integer_RS1_bypassEnables_bools_7 && (! (toplevel_execute_lane1_bypasser_integer_RS1_bypassEnables_range_4_to_6 || toplevel_execute_lane1_bypasser_integer_RS1_bypassEnables_range_0_to_3)));
    _zz_toplevel_execute_lane1_bypasser_integer_RS1_sel[8] = (toplevel_execute_lane1_bypasser_integer_RS1_bypassEnables_bools_8 && (! (toplevel_execute_lane1_bypasser_integer_RS1_bypassEnables_range_4_to_7 || toplevel_execute_lane1_bypasser_integer_RS1_bypassEnables_range_0_to_3)));
  end

  assign toplevel_execute_lane1_bypasser_integer_RS1_bypassEnables_range_0_to_1 = (|{toplevel_execute_lane1_bypasser_integer_RS1_bypassEnables_bools_1,toplevel_execute_lane1_bypasser_integer_RS1_bypassEnables_bools_0});
  assign toplevel_execute_lane1_bypasser_integer_RS1_bypassEnables_range_0_to_2 = (|{toplevel_execute_lane1_bypasser_integer_RS1_bypassEnables_bools_2,{toplevel_execute_lane1_bypasser_integer_RS1_bypassEnables_bools_1,toplevel_execute_lane1_bypasser_integer_RS1_bypassEnables_bools_0}});
  assign toplevel_execute_lane1_bypasser_integer_RS1_bypassEnables_range_0_to_3 = (|{toplevel_execute_lane1_bypasser_integer_RS1_bypassEnables_bools_3,{toplevel_execute_lane1_bypasser_integer_RS1_bypassEnables_bools_2,{toplevel_execute_lane1_bypasser_integer_RS1_bypassEnables_bools_1,toplevel_execute_lane1_bypasser_integer_RS1_bypassEnables_bools_0}}});
  assign toplevel_execute_lane1_bypasser_integer_RS1_bypassEnables_range_4_to_5 = (|{toplevel_execute_lane1_bypasser_integer_RS1_bypassEnables_bools_5,toplevel_execute_lane1_bypasser_integer_RS1_bypassEnables_bools_4});
  assign toplevel_execute_lane1_bypasser_integer_RS1_bypassEnables_range_4_to_6 = (|{toplevel_execute_lane1_bypasser_integer_RS1_bypassEnables_bools_6,{toplevel_execute_lane1_bypasser_integer_RS1_bypassEnables_bools_5,toplevel_execute_lane1_bypasser_integer_RS1_bypassEnables_bools_4}});
  assign toplevel_execute_lane1_bypasser_integer_RS1_bypassEnables_range_4_to_7 = (|{toplevel_execute_lane1_bypasser_integer_RS1_bypassEnables_bools_7,{toplevel_execute_lane1_bypasser_integer_RS1_bypassEnables_bools_6,{toplevel_execute_lane1_bypasser_integer_RS1_bypassEnables_bools_5,toplevel_execute_lane1_bypasser_integer_RS1_bypassEnables_bools_4}}});
  assign toplevel_execute_lane1_bypasser_integer_RS1_sel = _zz_toplevel_execute_lane1_bypasser_integer_RS1_sel;
  assign _zz_toplevel_execute_ctrl1_down_integer_RS1_lane1 = toplevel_execute_lane1_bypasser_integer_RS1_sel[8 : 1];
  always @(*) begin
    _zz_toplevel_execute_ctrl1_down_integer_RS1_lane1_1 = ((((_zz__zz_toplevel_execute_ctrl1_down_integer_RS1_lane1_1 ? toplevel_execute_ctrl2_down_lane1_integer_WriteBackPlugin_logic_DATA_lane1 : _zz__zz_toplevel_execute_ctrl1_down_integer_RS1_lane1_1_1) | (_zz__zz_toplevel_execute_ctrl1_down_integer_RS1_lane1_1_2 ? toplevel_execute_ctrl3_down_lane0_integer_WriteBackPlugin_logic_DATA_lane0 : _zz__zz_toplevel_execute_ctrl1_down_integer_RS1_lane1_1_3)) | ((_zz__zz_toplevel_execute_ctrl1_down_integer_RS1_lane1_1_4 ? toplevel_execute_ctrl3_down_lane1_integer_WriteBackPlugin_logic_DATA_lane1 : _zz__zz_toplevel_execute_ctrl1_down_integer_RS1_lane1_1_5) | (_zz__zz_toplevel_execute_ctrl1_down_integer_RS1_lane1_1_6 ? toplevel_execute_ctrl4_down_lane0_integer_WriteBackPlugin_logic_DATA_lane0 : _zz__zz_toplevel_execute_ctrl1_down_integer_RS1_lane1_1_7))) | (((_zz__zz_toplevel_execute_ctrl1_down_integer_RS1_lane1_1_8 ? toplevel_execute_ctrl4_down_lane1_integer_WriteBackPlugin_logic_DATA_lane1 : _zz__zz_toplevel_execute_ctrl1_down_integer_RS1_lane1_1_9) | (_zz__zz_toplevel_execute_ctrl1_down_integer_RS1_lane1_1_10 ? toplevel_execute_ctrl5_down_lane0_integer_WriteBackPlugin_logic_DATA_lane0 : _zz__zz_toplevel_execute_ctrl1_down_integer_RS1_lane1_1_11)) | ((_zz__zz_toplevel_execute_ctrl1_down_integer_RS1_lane1_1_12 ? toplevel_execute_ctrl5_down_lane1_integer_WriteBackPlugin_logic_DATA_lane1 : _zz__zz_toplevel_execute_ctrl1_down_integer_RS1_lane1_1_13) | (_zz__zz_toplevel_execute_ctrl1_down_integer_RS1_lane1_1_14 ? toplevel_execute_lane1_bypasser_integer_RS1_port_data : _zz__zz_toplevel_execute_ctrl1_down_integer_RS1_lane1_1_15))));
    if(when_ExecuteLanePlugin_l190_2) begin
      _zz_toplevel_execute_ctrl1_down_integer_RS1_lane1_1 = toplevel_execute_ctrl2_down_lane0_integer_WriteBackPlugin_logic_DATA_lane0;
    end
  end

  assign toplevel_execute_ctrl1_down_integer_RS1_lane1 = _zz_toplevel_execute_ctrl1_down_integer_RS1_lane1_1;
  assign when_ExecuteLanePlugin_l190_2 = toplevel_execute_lane1_bypasser_integer_RS1_sel[0];
  assign toplevel_execute_lane1_bypasser_integer_RS1_along_bypasses_0_checks_0_selfHit = (((toplevel_execute_ctrl3_up_LANE_SEL_lane0 && toplevel_execute_ctrl3_up_RD_ENABLE_lane0) && (toplevel_execute_ctrl3_down_RD_PHYS_lane0 == toplevel_execute_ctrl2_down_RS1_PHYS_lane1)) && 1'b1);
  assign toplevel_execute_lane1_bypasser_integer_RS1_along_bypasses_0_checks_0_hit = (toplevel_execute_lane1_bypasser_integer_RS1_along_bypasses_0_checks_0_selfHit && (! 1'b0));
  assign toplevel_execute_lane1_bypasser_integer_RS1_along_bypasses_0_checks_1_selfHit = (((toplevel_execute_ctrl4_up_LANE_SEL_lane0 && toplevel_execute_ctrl4_up_RD_ENABLE_lane0) && (toplevel_execute_ctrl4_down_RD_PHYS_lane0 == toplevel_execute_ctrl2_down_RS1_PHYS_lane1)) && 1'b1);
  assign toplevel_execute_lane1_bypasser_integer_RS1_along_bypasses_0_checks_1_youngerHits_0 = (((toplevel_execute_ctrl3_up_LANE_SEL_lane0 && toplevel_execute_ctrl3_up_RD_ENABLE_lane0) && (toplevel_execute_ctrl3_down_RD_PHYS_lane0 == toplevel_execute_ctrl2_down_RS1_PHYS_lane1)) && 1'b1);
  assign toplevel_execute_lane1_bypasser_integer_RS1_along_bypasses_0_checks_1_youngerHits_1 = (((toplevel_execute_ctrl3_up_LANE_SEL_lane1 && toplevel_execute_ctrl3_up_RD_ENABLE_lane1) && (toplevel_execute_ctrl3_down_RD_PHYS_lane1 == toplevel_execute_ctrl2_down_RS1_PHYS_lane1)) && 1'b1);
  assign toplevel_execute_lane1_bypasser_integer_RS1_along_bypasses_0_checks_1_hit = (toplevel_execute_lane1_bypasser_integer_RS1_along_bypasses_0_checks_1_selfHit && (! (|{toplevel_execute_lane1_bypasser_integer_RS1_along_bypasses_0_checks_1_youngerHits_1,toplevel_execute_lane1_bypasser_integer_RS1_along_bypasses_0_checks_1_youngerHits_0})));
  assign toplevel_execute_lane1_bypasser_integer_RS1_along_bypasses_0_checks_2_selfHit = (((toplevel_execute_ctrl3_up_LANE_SEL_lane1 && toplevel_execute_ctrl3_up_RD_ENABLE_lane1) && (toplevel_execute_ctrl3_down_RD_PHYS_lane1 == toplevel_execute_ctrl2_down_RS1_PHYS_lane1)) && 1'b1);
  assign toplevel_execute_lane1_bypasser_integer_RS1_along_bypasses_0_checks_2_hit = (toplevel_execute_lane1_bypasser_integer_RS1_along_bypasses_0_checks_2_selfHit && (! 1'b0));
  assign toplevel_execute_lane1_bypasser_integer_RS1_along_bypasses_0_checks_3_selfHit = (((toplevel_execute_ctrl4_up_LANE_SEL_lane1 && toplevel_execute_ctrl4_up_RD_ENABLE_lane1) && (toplevel_execute_ctrl4_down_RD_PHYS_lane1 == toplevel_execute_ctrl2_down_RS1_PHYS_lane1)) && 1'b1);
  assign toplevel_execute_lane1_bypasser_integer_RS1_along_bypasses_0_checks_3_youngerHits_0 = (((toplevel_execute_ctrl3_up_LANE_SEL_lane0 && toplevel_execute_ctrl3_up_RD_ENABLE_lane0) && (toplevel_execute_ctrl3_down_RD_PHYS_lane0 == toplevel_execute_ctrl2_down_RS1_PHYS_lane1)) && 1'b1);
  assign toplevel_execute_lane1_bypasser_integer_RS1_along_bypasses_0_checks_3_youngerHits_1 = (((toplevel_execute_ctrl3_up_LANE_SEL_lane1 && toplevel_execute_ctrl3_up_RD_ENABLE_lane1) && (toplevel_execute_ctrl3_down_RD_PHYS_lane1 == toplevel_execute_ctrl2_down_RS1_PHYS_lane1)) && 1'b1);
  assign toplevel_execute_lane1_bypasser_integer_RS1_along_bypasses_0_checks_3_hit = (toplevel_execute_lane1_bypasser_integer_RS1_along_bypasses_0_checks_3_selfHit && (! (|{toplevel_execute_lane1_bypasser_integer_RS1_along_bypasses_0_checks_3_youngerHits_1,toplevel_execute_lane1_bypasser_integer_RS1_along_bypasses_0_checks_3_youngerHits_0})));
  assign toplevel_execute_lane1_bypasser_integer_RS1_along_bypasses_0_hits = {toplevel_execute_lane1_bypasser_integer_RS1_along_bypasses_0_checks_3_hit,{toplevel_execute_lane1_bypasser_integer_RS1_along_bypasses_0_checks_2_hit,{toplevel_execute_lane1_bypasser_integer_RS1_along_bypasses_0_checks_1_hit,toplevel_execute_lane1_bypasser_integer_RS1_along_bypasses_0_checks_0_hit}}};
  assign _zz_toplevel_execute_ctrl2_integer_RS1_lane1_bypass = {toplevel_execute_lane1_bypasser_integer_RS1_along_bypasses_0_hits,(! (|toplevel_execute_lane1_bypasser_integer_RS1_along_bypasses_0_hits))};
  assign toplevel_execute_ctrl2_integer_RS1_lane1_bypass = ((((_zz_toplevel_execute_ctrl2_integer_RS1_lane1_bypass[0] ? toplevel_execute_ctrl2_up_integer_RS1_lane1 : 32'h0) | (_zz_toplevel_execute_ctrl2_integer_RS1_lane1_bypass[1] ? toplevel_execute_ctrl3_down_lane0_integer_WriteBackPlugin_logic_DATA_lane0 : 32'h0)) | ((_zz_toplevel_execute_ctrl2_integer_RS1_lane1_bypass[2] ? toplevel_execute_ctrl4_down_lane0_integer_WriteBackPlugin_logic_DATA_lane0 : 32'h0) | (_zz_toplevel_execute_ctrl2_integer_RS1_lane1_bypass[3] ? toplevel_execute_ctrl3_down_lane1_integer_WriteBackPlugin_logic_DATA_lane1 : 32'h0))) | (_zz_toplevel_execute_ctrl2_integer_RS1_lane1_bypass[4] ? toplevel_execute_ctrl4_down_lane1_integer_WriteBackPlugin_logic_DATA_lane1 : 32'h0));
  assign toplevel_execute_lane1_bypasser_integer_RS1_along_bypasses_1_checks_0_selfHit = (((toplevel_execute_ctrl4_up_LANE_SEL_lane0 && toplevel_execute_ctrl4_up_RD_ENABLE_lane0) && (toplevel_execute_ctrl4_down_RD_PHYS_lane0 == toplevel_execute_ctrl3_down_RS1_PHYS_lane1)) && 1'b1);
  assign toplevel_execute_lane1_bypasser_integer_RS1_along_bypasses_1_checks_0_hit = (toplevel_execute_lane1_bypasser_integer_RS1_along_bypasses_1_checks_0_selfHit && (! 1'b0));
  assign toplevel_execute_lane1_bypasser_integer_RS1_along_bypasses_1_checks_1_selfHit = (((toplevel_execute_ctrl4_up_LANE_SEL_lane1 && toplevel_execute_ctrl4_up_RD_ENABLE_lane1) && (toplevel_execute_ctrl4_down_RD_PHYS_lane1 == toplevel_execute_ctrl3_down_RS1_PHYS_lane1)) && 1'b1);
  assign toplevel_execute_lane1_bypasser_integer_RS1_along_bypasses_1_checks_1_hit = (toplevel_execute_lane1_bypasser_integer_RS1_along_bypasses_1_checks_1_selfHit && (! 1'b0));
  assign toplevel_execute_lane1_bypasser_integer_RS1_along_bypasses_1_hits = {toplevel_execute_lane1_bypasser_integer_RS1_along_bypasses_1_checks_1_hit,toplevel_execute_lane1_bypasser_integer_RS1_along_bypasses_1_checks_0_hit};
  assign _zz_toplevel_execute_ctrl3_integer_RS1_lane1_bypass = {toplevel_execute_lane1_bypasser_integer_RS1_along_bypasses_1_hits,(! (|toplevel_execute_lane1_bypasser_integer_RS1_along_bypasses_1_hits))};
  assign toplevel_execute_ctrl3_integer_RS1_lane1_bypass = (((_zz_toplevel_execute_ctrl3_integer_RS1_lane1_bypass[0] ? toplevel_execute_ctrl3_up_integer_RS1_lane1 : 32'h0) | (_zz_toplevel_execute_ctrl3_integer_RS1_lane1_bypass[1] ? toplevel_execute_ctrl4_down_lane0_integer_WriteBackPlugin_logic_DATA_lane0 : 32'h0)) | (_zz_toplevel_execute_ctrl3_integer_RS1_lane1_bypass[2] ? toplevel_execute_ctrl4_down_lane1_integer_WriteBackPlugin_logic_DATA_lane1 : 32'h0));
  assign toplevel_execute_lane1_bypasser_integer_RS2_port_valid = (! execute_freeze_valid);
  assign toplevel_execute_lane1_bypasser_integer_RS2_port_address = toplevel_execute_ctrl0_down_RS2_PHYS_lane1;
  always @(*) begin
    toplevel_execute_lane1_bypasser_integer_RS2_bypassEnables[0] = (((toplevel_execute_ctrl2_up_LANE_SEL_lane0 && toplevel_execute_ctrl2_up_RD_ENABLE_lane0) && (toplevel_execute_ctrl2_down_RD_PHYS_lane0 == toplevel_execute_ctrl1_down_RS2_PHYS_lane1)) && 1'b1);
    toplevel_execute_lane1_bypasser_integer_RS2_bypassEnables[1] = (((toplevel_execute_ctrl2_up_LANE_SEL_lane1 && toplevel_execute_ctrl2_up_RD_ENABLE_lane1) && (toplevel_execute_ctrl2_down_RD_PHYS_lane1 == toplevel_execute_ctrl1_down_RS2_PHYS_lane1)) && 1'b1);
    toplevel_execute_lane1_bypasser_integer_RS2_bypassEnables[2] = (((toplevel_execute_ctrl3_up_LANE_SEL_lane0 && toplevel_execute_ctrl3_up_RD_ENABLE_lane0) && (toplevel_execute_ctrl3_down_RD_PHYS_lane0 == toplevel_execute_ctrl1_down_RS2_PHYS_lane1)) && 1'b1);
    toplevel_execute_lane1_bypasser_integer_RS2_bypassEnables[3] = (((toplevel_execute_ctrl3_up_LANE_SEL_lane1 && toplevel_execute_ctrl3_up_RD_ENABLE_lane1) && (toplevel_execute_ctrl3_down_RD_PHYS_lane1 == toplevel_execute_ctrl1_down_RS2_PHYS_lane1)) && 1'b1);
    toplevel_execute_lane1_bypasser_integer_RS2_bypassEnables[4] = (((toplevel_execute_ctrl4_up_LANE_SEL_lane0 && toplevel_execute_ctrl4_up_RD_ENABLE_lane0) && (toplevel_execute_ctrl4_down_RD_PHYS_lane0 == toplevel_execute_ctrl1_down_RS2_PHYS_lane1)) && 1'b1);
    toplevel_execute_lane1_bypasser_integer_RS2_bypassEnables[5] = (((toplevel_execute_ctrl4_up_LANE_SEL_lane1 && toplevel_execute_ctrl4_up_RD_ENABLE_lane1) && (toplevel_execute_ctrl4_down_RD_PHYS_lane1 == toplevel_execute_ctrl1_down_RS2_PHYS_lane1)) && 1'b1);
    toplevel_execute_lane1_bypasser_integer_RS2_bypassEnables[6] = (((toplevel_execute_ctrl5_up_LANE_SEL_lane0 && toplevel_execute_ctrl5_up_RD_ENABLE_lane0) && (toplevel_execute_ctrl5_down_RD_PHYS_lane0 == toplevel_execute_ctrl1_down_RS2_PHYS_lane1)) && 1'b1);
    toplevel_execute_lane1_bypasser_integer_RS2_bypassEnables[7] = (((toplevel_execute_ctrl5_up_LANE_SEL_lane1 && toplevel_execute_ctrl5_up_RD_ENABLE_lane1) && (toplevel_execute_ctrl5_down_RD_PHYS_lane1 == toplevel_execute_ctrl1_down_RS2_PHYS_lane1)) && 1'b1);
    toplevel_execute_lane1_bypasser_integer_RS2_bypassEnables[8] = 1'b1;
  end

  assign _zz_toplevel_execute_lane1_bypasser_integer_RS2_bypassEnables_bools_0 = toplevel_execute_lane1_bypasser_integer_RS2_bypassEnables;
  assign toplevel_execute_lane1_bypasser_integer_RS2_bypassEnables_bools_0 = _zz_toplevel_execute_lane1_bypasser_integer_RS2_bypassEnables_bools_0[0];
  assign toplevel_execute_lane1_bypasser_integer_RS2_bypassEnables_bools_1 = _zz_toplevel_execute_lane1_bypasser_integer_RS2_bypassEnables_bools_0[1];
  assign toplevel_execute_lane1_bypasser_integer_RS2_bypassEnables_bools_2 = _zz_toplevel_execute_lane1_bypasser_integer_RS2_bypassEnables_bools_0[2];
  assign toplevel_execute_lane1_bypasser_integer_RS2_bypassEnables_bools_3 = _zz_toplevel_execute_lane1_bypasser_integer_RS2_bypassEnables_bools_0[3];
  assign toplevel_execute_lane1_bypasser_integer_RS2_bypassEnables_bools_4 = _zz_toplevel_execute_lane1_bypasser_integer_RS2_bypassEnables_bools_0[4];
  assign toplevel_execute_lane1_bypasser_integer_RS2_bypassEnables_bools_5 = _zz_toplevel_execute_lane1_bypasser_integer_RS2_bypassEnables_bools_0[5];
  assign toplevel_execute_lane1_bypasser_integer_RS2_bypassEnables_bools_6 = _zz_toplevel_execute_lane1_bypasser_integer_RS2_bypassEnables_bools_0[6];
  assign toplevel_execute_lane1_bypasser_integer_RS2_bypassEnables_bools_7 = _zz_toplevel_execute_lane1_bypasser_integer_RS2_bypassEnables_bools_0[7];
  assign toplevel_execute_lane1_bypasser_integer_RS2_bypassEnables_bools_8 = _zz_toplevel_execute_lane1_bypasser_integer_RS2_bypassEnables_bools_0[8];
  always @(*) begin
    _zz_toplevel_execute_lane1_bypasser_integer_RS2_sel[0] = (toplevel_execute_lane1_bypasser_integer_RS2_bypassEnables_bools_0 && (! 1'b0));
    _zz_toplevel_execute_lane1_bypasser_integer_RS2_sel[1] = (toplevel_execute_lane1_bypasser_integer_RS2_bypassEnables_bools_1 && (! toplevel_execute_lane1_bypasser_integer_RS2_bypassEnables_bools_0));
    _zz_toplevel_execute_lane1_bypasser_integer_RS2_sel[2] = (toplevel_execute_lane1_bypasser_integer_RS2_bypassEnables_bools_2 && (! toplevel_execute_lane1_bypasser_integer_RS2_bypassEnables_range_0_to_1));
    _zz_toplevel_execute_lane1_bypasser_integer_RS2_sel[3] = (toplevel_execute_lane1_bypasser_integer_RS2_bypassEnables_bools_3 && (! toplevel_execute_lane1_bypasser_integer_RS2_bypassEnables_range_0_to_2));
    _zz_toplevel_execute_lane1_bypasser_integer_RS2_sel[4] = (toplevel_execute_lane1_bypasser_integer_RS2_bypassEnables_bools_4 && (! toplevel_execute_lane1_bypasser_integer_RS2_bypassEnables_range_0_to_3));
    _zz_toplevel_execute_lane1_bypasser_integer_RS2_sel[5] = (toplevel_execute_lane1_bypasser_integer_RS2_bypassEnables_bools_5 && (! (toplevel_execute_lane1_bypasser_integer_RS2_bypassEnables_bools_4 || toplevel_execute_lane1_bypasser_integer_RS2_bypassEnables_range_0_to_3)));
    _zz_toplevel_execute_lane1_bypasser_integer_RS2_sel[6] = (toplevel_execute_lane1_bypasser_integer_RS2_bypassEnables_bools_6 && (! (toplevel_execute_lane1_bypasser_integer_RS2_bypassEnables_range_4_to_5 || toplevel_execute_lane1_bypasser_integer_RS2_bypassEnables_range_0_to_3)));
    _zz_toplevel_execute_lane1_bypasser_integer_RS2_sel[7] = (toplevel_execute_lane1_bypasser_integer_RS2_bypassEnables_bools_7 && (! (toplevel_execute_lane1_bypasser_integer_RS2_bypassEnables_range_4_to_6 || toplevel_execute_lane1_bypasser_integer_RS2_bypassEnables_range_0_to_3)));
    _zz_toplevel_execute_lane1_bypasser_integer_RS2_sel[8] = (toplevel_execute_lane1_bypasser_integer_RS2_bypassEnables_bools_8 && (! (toplevel_execute_lane1_bypasser_integer_RS2_bypassEnables_range_4_to_7 || toplevel_execute_lane1_bypasser_integer_RS2_bypassEnables_range_0_to_3)));
  end

  assign toplevel_execute_lane1_bypasser_integer_RS2_bypassEnables_range_0_to_1 = (|{toplevel_execute_lane1_bypasser_integer_RS2_bypassEnables_bools_1,toplevel_execute_lane1_bypasser_integer_RS2_bypassEnables_bools_0});
  assign toplevel_execute_lane1_bypasser_integer_RS2_bypassEnables_range_0_to_2 = (|{toplevel_execute_lane1_bypasser_integer_RS2_bypassEnables_bools_2,{toplevel_execute_lane1_bypasser_integer_RS2_bypassEnables_bools_1,toplevel_execute_lane1_bypasser_integer_RS2_bypassEnables_bools_0}});
  assign toplevel_execute_lane1_bypasser_integer_RS2_bypassEnables_range_0_to_3 = (|{toplevel_execute_lane1_bypasser_integer_RS2_bypassEnables_bools_3,{toplevel_execute_lane1_bypasser_integer_RS2_bypassEnables_bools_2,{toplevel_execute_lane1_bypasser_integer_RS2_bypassEnables_bools_1,toplevel_execute_lane1_bypasser_integer_RS2_bypassEnables_bools_0}}});
  assign toplevel_execute_lane1_bypasser_integer_RS2_bypassEnables_range_4_to_5 = (|{toplevel_execute_lane1_bypasser_integer_RS2_bypassEnables_bools_5,toplevel_execute_lane1_bypasser_integer_RS2_bypassEnables_bools_4});
  assign toplevel_execute_lane1_bypasser_integer_RS2_bypassEnables_range_4_to_6 = (|{toplevel_execute_lane1_bypasser_integer_RS2_bypassEnables_bools_6,{toplevel_execute_lane1_bypasser_integer_RS2_bypassEnables_bools_5,toplevel_execute_lane1_bypasser_integer_RS2_bypassEnables_bools_4}});
  assign toplevel_execute_lane1_bypasser_integer_RS2_bypassEnables_range_4_to_7 = (|{toplevel_execute_lane1_bypasser_integer_RS2_bypassEnables_bools_7,{toplevel_execute_lane1_bypasser_integer_RS2_bypassEnables_bools_6,{toplevel_execute_lane1_bypasser_integer_RS2_bypassEnables_bools_5,toplevel_execute_lane1_bypasser_integer_RS2_bypassEnables_bools_4}}});
  assign toplevel_execute_lane1_bypasser_integer_RS2_sel = _zz_toplevel_execute_lane1_bypasser_integer_RS2_sel;
  assign _zz_toplevel_execute_ctrl1_down_integer_RS2_lane1 = toplevel_execute_lane1_bypasser_integer_RS2_sel[8 : 1];
  always @(*) begin
    _zz_toplevel_execute_ctrl1_down_integer_RS2_lane1_1 = ((((_zz__zz_toplevel_execute_ctrl1_down_integer_RS2_lane1_1 ? toplevel_execute_ctrl2_down_lane1_integer_WriteBackPlugin_logic_DATA_lane1 : _zz__zz_toplevel_execute_ctrl1_down_integer_RS2_lane1_1_1) | (_zz__zz_toplevel_execute_ctrl1_down_integer_RS2_lane1_1_2 ? toplevel_execute_ctrl3_down_lane0_integer_WriteBackPlugin_logic_DATA_lane0 : _zz__zz_toplevel_execute_ctrl1_down_integer_RS2_lane1_1_3)) | ((_zz__zz_toplevel_execute_ctrl1_down_integer_RS2_lane1_1_4 ? toplevel_execute_ctrl3_down_lane1_integer_WriteBackPlugin_logic_DATA_lane1 : _zz__zz_toplevel_execute_ctrl1_down_integer_RS2_lane1_1_5) | (_zz__zz_toplevel_execute_ctrl1_down_integer_RS2_lane1_1_6 ? toplevel_execute_ctrl4_down_lane0_integer_WriteBackPlugin_logic_DATA_lane0 : _zz__zz_toplevel_execute_ctrl1_down_integer_RS2_lane1_1_7))) | (((_zz__zz_toplevel_execute_ctrl1_down_integer_RS2_lane1_1_8 ? toplevel_execute_ctrl4_down_lane1_integer_WriteBackPlugin_logic_DATA_lane1 : _zz__zz_toplevel_execute_ctrl1_down_integer_RS2_lane1_1_9) | (_zz__zz_toplevel_execute_ctrl1_down_integer_RS2_lane1_1_10 ? toplevel_execute_ctrl5_down_lane0_integer_WriteBackPlugin_logic_DATA_lane0 : _zz__zz_toplevel_execute_ctrl1_down_integer_RS2_lane1_1_11)) | ((_zz__zz_toplevel_execute_ctrl1_down_integer_RS2_lane1_1_12 ? toplevel_execute_ctrl5_down_lane1_integer_WriteBackPlugin_logic_DATA_lane1 : _zz__zz_toplevel_execute_ctrl1_down_integer_RS2_lane1_1_13) | (_zz__zz_toplevel_execute_ctrl1_down_integer_RS2_lane1_1_14 ? toplevel_execute_lane1_bypasser_integer_RS2_port_data : _zz__zz_toplevel_execute_ctrl1_down_integer_RS2_lane1_1_15))));
    if(when_ExecuteLanePlugin_l190_3) begin
      _zz_toplevel_execute_ctrl1_down_integer_RS2_lane1_1 = toplevel_execute_ctrl2_down_lane0_integer_WriteBackPlugin_logic_DATA_lane0;
    end
  end

  assign toplevel_execute_ctrl1_down_integer_RS2_lane1 = _zz_toplevel_execute_ctrl1_down_integer_RS2_lane1_1;
  assign when_ExecuteLanePlugin_l190_3 = toplevel_execute_lane1_bypasser_integer_RS2_sel[0];
  assign toplevel_execute_lane1_bypasser_integer_RS2_along_bypasses_0_checks_0_selfHit = (((toplevel_execute_ctrl3_up_LANE_SEL_lane0 && toplevel_execute_ctrl3_up_RD_ENABLE_lane0) && (toplevel_execute_ctrl3_down_RD_PHYS_lane0 == toplevel_execute_ctrl2_down_RS2_PHYS_lane1)) && 1'b1);
  assign toplevel_execute_lane1_bypasser_integer_RS2_along_bypasses_0_checks_0_hit = (toplevel_execute_lane1_bypasser_integer_RS2_along_bypasses_0_checks_0_selfHit && (! 1'b0));
  assign toplevel_execute_lane1_bypasser_integer_RS2_along_bypasses_0_checks_1_selfHit = (((toplevel_execute_ctrl4_up_LANE_SEL_lane0 && toplevel_execute_ctrl4_up_RD_ENABLE_lane0) && (toplevel_execute_ctrl4_down_RD_PHYS_lane0 == toplevel_execute_ctrl2_down_RS2_PHYS_lane1)) && 1'b1);
  assign toplevel_execute_lane1_bypasser_integer_RS2_along_bypasses_0_checks_1_youngerHits_0 = (((toplevel_execute_ctrl3_up_LANE_SEL_lane0 && toplevel_execute_ctrl3_up_RD_ENABLE_lane0) && (toplevel_execute_ctrl3_down_RD_PHYS_lane0 == toplevel_execute_ctrl2_down_RS2_PHYS_lane1)) && 1'b1);
  assign toplevel_execute_lane1_bypasser_integer_RS2_along_bypasses_0_checks_1_youngerHits_1 = (((toplevel_execute_ctrl3_up_LANE_SEL_lane1 && toplevel_execute_ctrl3_up_RD_ENABLE_lane1) && (toplevel_execute_ctrl3_down_RD_PHYS_lane1 == toplevel_execute_ctrl2_down_RS2_PHYS_lane1)) && 1'b1);
  assign toplevel_execute_lane1_bypasser_integer_RS2_along_bypasses_0_checks_1_hit = (toplevel_execute_lane1_bypasser_integer_RS2_along_bypasses_0_checks_1_selfHit && (! (|{toplevel_execute_lane1_bypasser_integer_RS2_along_bypasses_0_checks_1_youngerHits_1,toplevel_execute_lane1_bypasser_integer_RS2_along_bypasses_0_checks_1_youngerHits_0})));
  assign toplevel_execute_lane1_bypasser_integer_RS2_along_bypasses_0_checks_2_selfHit = (((toplevel_execute_ctrl3_up_LANE_SEL_lane1 && toplevel_execute_ctrl3_up_RD_ENABLE_lane1) && (toplevel_execute_ctrl3_down_RD_PHYS_lane1 == toplevel_execute_ctrl2_down_RS2_PHYS_lane1)) && 1'b1);
  assign toplevel_execute_lane1_bypasser_integer_RS2_along_bypasses_0_checks_2_hit = (toplevel_execute_lane1_bypasser_integer_RS2_along_bypasses_0_checks_2_selfHit && (! 1'b0));
  assign toplevel_execute_lane1_bypasser_integer_RS2_along_bypasses_0_checks_3_selfHit = (((toplevel_execute_ctrl4_up_LANE_SEL_lane1 && toplevel_execute_ctrl4_up_RD_ENABLE_lane1) && (toplevel_execute_ctrl4_down_RD_PHYS_lane1 == toplevel_execute_ctrl2_down_RS2_PHYS_lane1)) && 1'b1);
  assign toplevel_execute_lane1_bypasser_integer_RS2_along_bypasses_0_checks_3_youngerHits_0 = (((toplevel_execute_ctrl3_up_LANE_SEL_lane0 && toplevel_execute_ctrl3_up_RD_ENABLE_lane0) && (toplevel_execute_ctrl3_down_RD_PHYS_lane0 == toplevel_execute_ctrl2_down_RS2_PHYS_lane1)) && 1'b1);
  assign toplevel_execute_lane1_bypasser_integer_RS2_along_bypasses_0_checks_3_youngerHits_1 = (((toplevel_execute_ctrl3_up_LANE_SEL_lane1 && toplevel_execute_ctrl3_up_RD_ENABLE_lane1) && (toplevel_execute_ctrl3_down_RD_PHYS_lane1 == toplevel_execute_ctrl2_down_RS2_PHYS_lane1)) && 1'b1);
  assign toplevel_execute_lane1_bypasser_integer_RS2_along_bypasses_0_checks_3_hit = (toplevel_execute_lane1_bypasser_integer_RS2_along_bypasses_0_checks_3_selfHit && (! (|{toplevel_execute_lane1_bypasser_integer_RS2_along_bypasses_0_checks_3_youngerHits_1,toplevel_execute_lane1_bypasser_integer_RS2_along_bypasses_0_checks_3_youngerHits_0})));
  assign toplevel_execute_lane1_bypasser_integer_RS2_along_bypasses_0_hits = {toplevel_execute_lane1_bypasser_integer_RS2_along_bypasses_0_checks_3_hit,{toplevel_execute_lane1_bypasser_integer_RS2_along_bypasses_0_checks_2_hit,{toplevel_execute_lane1_bypasser_integer_RS2_along_bypasses_0_checks_1_hit,toplevel_execute_lane1_bypasser_integer_RS2_along_bypasses_0_checks_0_hit}}};
  assign _zz_toplevel_execute_ctrl2_integer_RS2_lane1_bypass = {toplevel_execute_lane1_bypasser_integer_RS2_along_bypasses_0_hits,(! (|toplevel_execute_lane1_bypasser_integer_RS2_along_bypasses_0_hits))};
  assign toplevel_execute_ctrl2_integer_RS2_lane1_bypass = ((((_zz_toplevel_execute_ctrl2_integer_RS2_lane1_bypass[0] ? toplevel_execute_ctrl2_up_integer_RS2_lane1 : 32'h0) | (_zz_toplevel_execute_ctrl2_integer_RS2_lane1_bypass[1] ? toplevel_execute_ctrl3_down_lane0_integer_WriteBackPlugin_logic_DATA_lane0 : 32'h0)) | ((_zz_toplevel_execute_ctrl2_integer_RS2_lane1_bypass[2] ? toplevel_execute_ctrl4_down_lane0_integer_WriteBackPlugin_logic_DATA_lane0 : 32'h0) | (_zz_toplevel_execute_ctrl2_integer_RS2_lane1_bypass[3] ? toplevel_execute_ctrl3_down_lane1_integer_WriteBackPlugin_logic_DATA_lane1 : 32'h0))) | (_zz_toplevel_execute_ctrl2_integer_RS2_lane1_bypass[4] ? toplevel_execute_ctrl4_down_lane1_integer_WriteBackPlugin_logic_DATA_lane1 : 32'h0));
  assign toplevel_execute_lane1_bypasser_integer_RS2_along_bypasses_1_checks_0_selfHit = (((toplevel_execute_ctrl4_up_LANE_SEL_lane0 && toplevel_execute_ctrl4_up_RD_ENABLE_lane0) && (toplevel_execute_ctrl4_down_RD_PHYS_lane0 == toplevel_execute_ctrl3_down_RS2_PHYS_lane1)) && 1'b1);
  assign toplevel_execute_lane1_bypasser_integer_RS2_along_bypasses_1_checks_0_hit = (toplevel_execute_lane1_bypasser_integer_RS2_along_bypasses_1_checks_0_selfHit && (! 1'b0));
  assign toplevel_execute_lane1_bypasser_integer_RS2_along_bypasses_1_checks_1_selfHit = (((toplevel_execute_ctrl4_up_LANE_SEL_lane1 && toplevel_execute_ctrl4_up_RD_ENABLE_lane1) && (toplevel_execute_ctrl4_down_RD_PHYS_lane1 == toplevel_execute_ctrl3_down_RS2_PHYS_lane1)) && 1'b1);
  assign toplevel_execute_lane1_bypasser_integer_RS2_along_bypasses_1_checks_1_hit = (toplevel_execute_lane1_bypasser_integer_RS2_along_bypasses_1_checks_1_selfHit && (! 1'b0));
  assign toplevel_execute_lane1_bypasser_integer_RS2_along_bypasses_1_hits = {toplevel_execute_lane1_bypasser_integer_RS2_along_bypasses_1_checks_1_hit,toplevel_execute_lane1_bypasser_integer_RS2_along_bypasses_1_checks_0_hit};
  assign _zz_toplevel_execute_ctrl3_integer_RS2_lane1_bypass = {toplevel_execute_lane1_bypasser_integer_RS2_along_bypasses_1_hits,(! (|toplevel_execute_lane1_bypasser_integer_RS2_along_bypasses_1_hits))};
  assign toplevel_execute_ctrl3_integer_RS2_lane1_bypass = (((_zz_toplevel_execute_ctrl3_integer_RS2_lane1_bypass[0] ? toplevel_execute_ctrl3_up_integer_RS2_lane1 : 32'h0) | (_zz_toplevel_execute_ctrl3_integer_RS2_lane1_bypass[1] ? toplevel_execute_ctrl4_down_lane0_integer_WriteBackPlugin_logic_DATA_lane0 : 32'h0)) | (_zz_toplevel_execute_ctrl3_integer_RS2_lane1_bypass[2] ? toplevel_execute_ctrl4_down_lane1_integer_WriteBackPlugin_logic_DATA_lane1 : 32'h0));
  assign execute_lane1_logic_completions_onCtrl_0_port_valid = (((toplevel_execute_ctrl2_down_LANE_SEL_lane1 && toplevel_execute_ctrl2_down_isReady) && (! toplevel_execute_lane1_ctrls_2_downIsCancel)) && toplevel_execute_ctrl2_down_execute_lane1_logic_completions_onCtrl_0_ENABLE_lane1);
  assign execute_lane1_logic_completions_onCtrl_0_port_payload_uopId = toplevel_execute_ctrl2_down_Decode_UOP_ID_lane1;
  assign execute_lane1_logic_completions_onCtrl_0_port_payload_trap = toplevel_execute_ctrl2_down_TRAP_lane1;
  assign execute_lane1_logic_completions_onCtrl_0_port_payload_commit = toplevel_execute_ctrl2_down_COMMIT_lane1;
  assign execute_lane1_logic_completions_onCtrl_1_port_valid = (((toplevel_execute_ctrl3_down_LANE_SEL_lane1 && toplevel_execute_ctrl3_down_isReady) && (! toplevel_execute_lane1_ctrls_3_downIsCancel)) && toplevel_execute_ctrl3_down_execute_lane1_logic_completions_onCtrl_1_ENABLE_lane1);
  assign execute_lane1_logic_completions_onCtrl_1_port_payload_uopId = toplevel_execute_ctrl3_down_Decode_UOP_ID_lane1;
  assign execute_lane1_logic_completions_onCtrl_1_port_payload_trap = toplevel_execute_ctrl3_down_TRAP_lane1;
  assign execute_lane1_logic_completions_onCtrl_1_port_payload_commit = toplevel_execute_ctrl3_down_COMMIT_lane1;
  assign execute_lane1_logic_completions_onCtrl_2_port_valid = (((toplevel_execute_ctrl4_down_LANE_SEL_lane1 && toplevel_execute_ctrl4_down_isReady) && (! toplevel_execute_lane1_ctrls_4_downIsCancel)) && toplevel_execute_ctrl4_down_execute_lane1_logic_completions_onCtrl_2_ENABLE_lane1);
  assign execute_lane1_logic_completions_onCtrl_2_port_payload_uopId = toplevel_execute_ctrl4_down_Decode_UOP_ID_lane1;
  assign execute_lane1_logic_completions_onCtrl_2_port_payload_trap = toplevel_execute_ctrl4_down_TRAP_lane1;
  assign execute_lane1_logic_completions_onCtrl_2_port_payload_commit = toplevel_execute_ctrl4_down_COMMIT_lane1;
  assign execute_lane1_logic_decoding_decodingBits = {toplevel_execute_ctrl1_down_execute_lane1_LAYER_SEL_lane1,toplevel_execute_ctrl1_down_Decode_UOP_lane1};
  assign _zz_toplevel_execute_ctrl1_down_execute_lane1_logic_completions_onCtrl_0_ENABLE_lane1 = ((execute_lane1_logic_decoding_decodingBits & 33'h100001040) == 33'h100000000);
  assign _zz_toplevel_execute_ctrl1_down_execute_lane1_logic_completions_onCtrl_0_ENABLE_lane1_1 = ((execute_lane1_logic_decoding_decodingBits & 33'h100000044) == 33'h100000004);
  assign _zz_toplevel_execute_ctrl1_down_execute_lane1_logic_completions_onCtrl_0_ENABLE_lane1_2 = ((execute_lane1_logic_decoding_decodingBits & 33'h100002040) == 33'h100002000);
  always @(*) begin
    toplevel_execute_ctrl1_down_early1_IntAluPlugin_SEL_lane1 = _zz_toplevel_execute_ctrl1_down_early1_IntAluPlugin_SEL_lane1[0];
    if(toplevel_execute_ctrl1_down_TRAP_lane1) begin
      toplevel_execute_ctrl1_down_early1_IntAluPlugin_SEL_lane1 = 1'b0;
    end
  end

  always @(*) begin
    toplevel_execute_ctrl1_down_early1_BarrelShifterPlugin_SEL_lane1 = _zz_toplevel_execute_ctrl1_down_early1_BarrelShifterPlugin_SEL_lane1[0];
    if(toplevel_execute_ctrl1_down_TRAP_lane1) begin
      toplevel_execute_ctrl1_down_early1_BarrelShifterPlugin_SEL_lane1 = 1'b0;
    end
  end

  assign _zz_toplevel_execute_ctrl1_down_execute_lane1_logic_completions_onCtrl_1_ENABLE_lane1 = ((execute_lane1_logic_decoding_decodingBits & 33'h100000010) == 33'h100000000);
  always @(*) begin
    toplevel_execute_ctrl1_down_early1_BranchPlugin_SEL_lane1 = _zz_toplevel_execute_ctrl1_down_early1_BranchPlugin_SEL_lane1[0];
    if(toplevel_execute_ctrl1_down_TRAP_lane1) begin
      toplevel_execute_ctrl1_down_early1_BranchPlugin_SEL_lane1 = 1'b0;
    end
  end

  always @(*) begin
    toplevel_execute_ctrl1_down_late1_IntAluPlugin_SEL_lane1 = _zz_toplevel_execute_ctrl1_down_late1_IntAluPlugin_SEL_lane1[0];
    if(toplevel_execute_ctrl1_down_TRAP_lane1) begin
      toplevel_execute_ctrl1_down_late1_IntAluPlugin_SEL_lane1 = 1'b0;
    end
  end

  always @(*) begin
    toplevel_execute_ctrl1_down_late1_BarrelShifterPlugin_SEL_lane1 = _zz_toplevel_execute_ctrl1_down_late1_BarrelShifterPlugin_SEL_lane1[0];
    if(toplevel_execute_ctrl1_down_TRAP_lane1) begin
      toplevel_execute_ctrl1_down_late1_BarrelShifterPlugin_SEL_lane1 = 1'b0;
    end
  end

  assign _zz_toplevel_execute_ctrl1_down_late1_BranchPlugin_SEL_lane1 = ((execute_lane1_logic_decoding_decodingBits & 33'h100000010) == 33'h0);
  always @(*) begin
    toplevel_execute_ctrl1_down_late1_BranchPlugin_SEL_lane1 = _zz_toplevel_execute_ctrl1_down_late1_BranchPlugin_SEL_lane1_1[0];
    if(toplevel_execute_ctrl1_down_TRAP_lane1) begin
      toplevel_execute_ctrl1_down_late1_BranchPlugin_SEL_lane1 = 1'b0;
    end
  end

  assign _zz_toplevel_execute_ctrl1_down_late1_SrcPlugin_logic_SRC2_CTRL_lane1 = ((execute_lane1_logic_decoding_decodingBits & 33'h000000004) == 33'h000000004);
  always @(*) begin
    toplevel_execute_ctrl1_down_lane1_integer_WriteBackPlugin_SEL_lane1 = _zz_toplevel_execute_ctrl1_down_lane1_integer_WriteBackPlugin_SEL_lane1[0];
    if(toplevel_execute_ctrl1_down_TRAP_lane1) begin
      toplevel_execute_ctrl1_down_lane1_integer_WriteBackPlugin_SEL_lane1 = 1'b0;
    end
  end

  always @(*) begin
    toplevel_execute_ctrl1_down_COMPLETION_AT_2_lane1 = _zz_toplevel_execute_ctrl1_down_COMPLETION_AT_2_lane1[0];
    if(toplevel_execute_ctrl1_down_TRAP_lane1) begin
      toplevel_execute_ctrl1_down_COMPLETION_AT_2_lane1 = 1'b0;
    end
  end

  assign _zz_toplevel_execute_ctrl1_down_execute_lane1_logic_completions_onCtrl_1_ENABLE_lane1_1 = ((execute_lane1_logic_decoding_decodingBits & 33'h100003004) == 33'h100001000);
  always @(*) begin
    toplevel_execute_ctrl1_down_COMPLETION_AT_3_lane1 = _zz_toplevel_execute_ctrl1_down_COMPLETION_AT_3_lane1[0];
    if(toplevel_execute_ctrl1_down_TRAP_lane1) begin
      toplevel_execute_ctrl1_down_COMPLETION_AT_3_lane1 = 1'b0;
    end
  end

  assign _zz_toplevel_execute_ctrl1_down_execute_lane1_logic_completions_onCtrl_2_ENABLE_lane1 = ((execute_lane1_logic_decoding_decodingBits & 33'h100000000) == 33'h0);
  always @(*) begin
    toplevel_execute_ctrl1_down_COMPLETION_AT_4_lane1 = _zz_toplevel_execute_ctrl1_down_COMPLETION_AT_4_lane1[0];
    if(toplevel_execute_ctrl1_down_TRAP_lane1) begin
      toplevel_execute_ctrl1_down_COMPLETION_AT_4_lane1 = 1'b0;
    end
  end

  always @(*) begin
    toplevel_execute_ctrl1_down_execute_lane1_logic_completions_onCtrl_0_ENABLE_lane1 = _zz_toplevel_execute_ctrl1_down_execute_lane1_logic_completions_onCtrl_0_ENABLE_lane1_3[0];
    if(toplevel_execute_ctrl1_down_TRAP_lane1) begin
      toplevel_execute_ctrl1_down_execute_lane1_logic_completions_onCtrl_0_ENABLE_lane1 = 1'b0;
    end
  end

  always @(*) begin
    toplevel_execute_ctrl1_down_execute_lane1_logic_completions_onCtrl_1_ENABLE_lane1 = _zz_toplevel_execute_ctrl1_down_execute_lane1_logic_completions_onCtrl_1_ENABLE_lane1_2[0];
    if(toplevel_execute_ctrl1_down_TRAP_lane1) begin
      toplevel_execute_ctrl1_down_execute_lane1_logic_completions_onCtrl_1_ENABLE_lane1 = 1'b0;
    end
  end

  always @(*) begin
    toplevel_execute_ctrl1_down_execute_lane1_logic_completions_onCtrl_2_ENABLE_lane1 = _zz_toplevel_execute_ctrl1_down_execute_lane1_logic_completions_onCtrl_2_ENABLE_lane1_1[0];
    if(toplevel_execute_ctrl1_down_TRAP_lane1) begin
      toplevel_execute_ctrl1_down_execute_lane1_logic_completions_onCtrl_2_ENABLE_lane1 = 1'b0;
    end
  end

  assign _zz_toplevel_execute_ctrl1_down_late1_IntAluPlugin_ALU_ADD_SUB_lane1 = ((execute_lane1_logic_decoding_decodingBits & 33'h000006000) == 33'h0);
  assign toplevel_execute_ctrl1_down_early1_IntAluPlugin_ALU_ADD_SUB_lane1 = _zz_toplevel_execute_ctrl1_down_early1_IntAluPlugin_ALU_ADD_SUB_lane1[0];
  assign _zz_toplevel_execute_ctrl1_down_late1_IntAluPlugin_ALU_SLTX_lane1 = ((execute_lane1_logic_decoding_decodingBits & 33'h000006004) == 33'h000002000);
  assign toplevel_execute_ctrl1_down_early1_IntAluPlugin_ALU_SLTX_lane1 = _zz_toplevel_execute_ctrl1_down_early1_IntAluPlugin_ALU_SLTX_lane1[0];
  assign _zz_toplevel_execute_ctrl1_down_late1_IntAluPlugin_ALU_BITWISE_CTRL_lane1 = ((execute_lane1_logic_decoding_decodingBits & 33'h000003000) == 33'h000002000);
  assign _zz_toplevel_execute_ctrl1_down_BarrelShifterPlugin_LEFT_lane1 = ((execute_lane1_logic_decoding_decodingBits & 33'h000004000) == 33'h0);
  assign _zz_toplevel_execute_ctrl1_down_late1_IntAluPlugin_ALU_BITWISE_CTRL_lane1_1 = ((execute_lane1_logic_decoding_decodingBits & 33'h000001000) == 33'h000001000);
  assign _zz_toplevel_execute_ctrl1_down_early1_IntAluPlugin_ALU_BITWISE_CTRL_lane1_1 = {(|{_zz_toplevel_execute_ctrl1_down_late1_IntAluPlugin_ALU_BITWISE_CTRL_lane1_1,{_zz_toplevel_execute_ctrl1_down_late1_SrcPlugin_logic_SRC2_CTRL_lane1,_zz_toplevel_execute_ctrl1_down_BarrelShifterPlugin_LEFT_lane1}}),(|{_zz_toplevel_execute_ctrl1_down_late1_SrcPlugin_logic_SRC2_CTRL_lane1,{_zz_toplevel_execute_ctrl1_down_BarrelShifterPlugin_LEFT_lane1,_zz_toplevel_execute_ctrl1_down_late1_IntAluPlugin_ALU_BITWISE_CTRL_lane1}})};
  assign _zz_toplevel_execute_ctrl1_down_early1_IntAluPlugin_ALU_BITWISE_CTRL_lane1 = _zz_toplevel_execute_ctrl1_down_early1_IntAluPlugin_ALU_BITWISE_CTRL_lane1_1;
  assign _zz_toplevel_execute_ctrl1_down_early1_IntAluPlugin_ALU_BITWISE_CTRL_lane1_2 = _zz_toplevel_execute_ctrl1_down_early1_IntAluPlugin_ALU_BITWISE_CTRL_lane1;
  assign toplevel_execute_ctrl1_down_early1_IntAluPlugin_ALU_BITWISE_CTRL_lane1 = _zz_toplevel_execute_ctrl1_down_early1_IntAluPlugin_ALU_BITWISE_CTRL_lane1_2;
  assign _zz_toplevel_execute_ctrl1_down_SrcStageables_REVERT_lane1 = ((execute_lane1_logic_decoding_decodingBits & 33'h000000010) == 33'h0);
  assign toplevel_execute_ctrl1_down_SrcStageables_REVERT_lane1 = _zz_toplevel_execute_ctrl1_down_SrcStageables_REVERT_lane1_1[0];
  assign toplevel_execute_ctrl1_down_SrcStageables_ZERO_lane1 = _zz_toplevel_execute_ctrl1_down_SrcStageables_ZERO_lane1[0];
  assign toplevel_execute_ctrl1_down_early1_SrcPlugin_logic_SRC1_CTRL_lane1 = (|((execute_lane1_logic_decoding_decodingBits & 33'h000000044) == 33'h000000004));
  assign _zz_toplevel_execute_ctrl1_down_late1_SrcPlugin_logic_SRC2_CTRL_lane1_1 = ((execute_lane1_logic_decoding_decodingBits & 33'h000000024) == 33'h0);
  assign toplevel_execute_ctrl1_down_early1_SrcPlugin_logic_SRC2_CTRL_lane1 = {(|_zz_toplevel_execute_ctrl1_down_late1_SrcPlugin_logic_SRC2_CTRL_lane1),(|_zz_toplevel_execute_ctrl1_down_late1_SrcPlugin_logic_SRC2_CTRL_lane1_1)};
  assign toplevel_execute_ctrl1_down_lane1_IntFormatPlugin_logic_SIGNED_lane1 = _zz_toplevel_execute_ctrl1_down_lane1_IntFormatPlugin_logic_SIGNED_lane1[0];
  assign toplevel_execute_ctrl1_down_BYPASSED_AT_2_lane1 = _zz_toplevel_execute_ctrl1_down_BYPASSED_AT_2_lane1[0];
  assign toplevel_execute_ctrl1_down_BYPASSED_AT_3_lane1 = _zz_toplevel_execute_ctrl1_down_BYPASSED_AT_3_lane1[0];
  assign toplevel_execute_ctrl1_down_MAY_FLUSH_PRECISE_3_lane1 = _zz_toplevel_execute_ctrl1_down_MAY_FLUSH_PRECISE_3_lane1[0];
  assign toplevel_execute_ctrl1_down_MAY_FLUSH_PRECISE_4_lane1 = _zz_toplevel_execute_ctrl1_down_MAY_FLUSH_PRECISE_4_lane1[0];
  assign toplevel_execute_ctrl1_down_SrcStageables_UNSIGNED_lane1 = _zz_toplevel_execute_ctrl1_down_SrcStageables_UNSIGNED_lane1[0];
  assign toplevel_execute_ctrl1_down_BarrelShifterPlugin_LEFT_lane1 = _zz_toplevel_execute_ctrl1_down_BarrelShifterPlugin_LEFT_lane1_1[0];
  assign toplevel_execute_ctrl1_down_BarrelShifterPlugin_SIGNED_lane1 = _zz_toplevel_execute_ctrl1_down_BarrelShifterPlugin_SIGNED_lane1[0];
  assign _zz_toplevel_execute_ctrl1_down_BranchPlugin_BRANCH_CTRL_lane1_1 = {(|((execute_lane1_logic_decoding_decodingBits & 33'h00000000c) == 33'h000000004)),(|((execute_lane1_logic_decoding_decodingBits & 33'h000000008) == 33'h000000008))};
  assign _zz_toplevel_execute_ctrl1_down_BranchPlugin_BRANCH_CTRL_lane1 = _zz_toplevel_execute_ctrl1_down_BranchPlugin_BRANCH_CTRL_lane1_1;
  assign _zz_toplevel_execute_ctrl1_down_BranchPlugin_BRANCH_CTRL_lane1_2 = _zz_toplevel_execute_ctrl1_down_BranchPlugin_BRANCH_CTRL_lane1;
  assign toplevel_execute_ctrl1_down_BranchPlugin_BRANCH_CTRL_lane1 = _zz_toplevel_execute_ctrl1_down_BranchPlugin_BRANCH_CTRL_lane1_2;
  assign toplevel_execute_ctrl1_down_late1_IntAluPlugin_ALU_ADD_SUB_lane1 = _zz_toplevel_execute_ctrl1_down_late1_IntAluPlugin_ALU_ADD_SUB_lane1_1[0];
  assign toplevel_execute_ctrl1_down_late1_IntAluPlugin_ALU_SLTX_lane1 = _zz_toplevel_execute_ctrl1_down_late1_IntAluPlugin_ALU_SLTX_lane1_1[0];
  assign _zz_toplevel_execute_ctrl1_down_late1_IntAluPlugin_ALU_BITWISE_CTRL_lane1_3 = {(|{_zz_toplevel_execute_ctrl1_down_late1_IntAluPlugin_ALU_BITWISE_CTRL_lane1_1,{_zz_toplevel_execute_ctrl1_down_late1_SrcPlugin_logic_SRC2_CTRL_lane1,_zz_toplevel_execute_ctrl1_down_BarrelShifterPlugin_LEFT_lane1}}),(|{_zz_toplevel_execute_ctrl1_down_late1_SrcPlugin_logic_SRC2_CTRL_lane1,{_zz_toplevel_execute_ctrl1_down_BarrelShifterPlugin_LEFT_lane1,_zz_toplevel_execute_ctrl1_down_late1_IntAluPlugin_ALU_BITWISE_CTRL_lane1}})};
  assign _zz_toplevel_execute_ctrl1_down_late1_IntAluPlugin_ALU_BITWISE_CTRL_lane1_2 = _zz_toplevel_execute_ctrl1_down_late1_IntAluPlugin_ALU_BITWISE_CTRL_lane1_3;
  assign _zz_toplevel_execute_ctrl1_down_late1_IntAluPlugin_ALU_BITWISE_CTRL_lane1_4 = _zz_toplevel_execute_ctrl1_down_late1_IntAluPlugin_ALU_BITWISE_CTRL_lane1_2;
  assign toplevel_execute_ctrl1_down_late1_IntAluPlugin_ALU_BITWISE_CTRL_lane1 = _zz_toplevel_execute_ctrl1_down_late1_IntAluPlugin_ALU_BITWISE_CTRL_lane1_4;
  assign toplevel_execute_ctrl1_down_late1_SrcPlugin_logic_SRC1_CTRL_lane1 = (|_zz_toplevel_execute_ctrl1_down_late1_SrcPlugin_logic_SRC2_CTRL_lane1);
  assign toplevel_execute_ctrl1_down_late1_SrcPlugin_logic_SRC2_CTRL_lane1 = {(|_zz_toplevel_execute_ctrl1_down_late1_SrcPlugin_logic_SRC2_CTRL_lane1),(|_zz_toplevel_execute_ctrl1_down_late1_SrcPlugin_logic_SRC2_CTRL_lane1_1)};
  assign when_ExecuteLanePlugin_l300_5 = (|{(late1_BranchPlugin_logic_flushPort_valid && 1'b1),{(early1_BranchPlugin_logic_flushPort_valid && 1'b1),{(late0_BranchPlugin_logic_flushPort_valid && 1'b1),{(early0_EnvPlugin_logic_flushPort_valid && 1'b1),{(CsrAccessPlugin_logic_flushPort_valid && 1'b1),{(early0_BranchPlugin_logic_flushPort_valid && 1'b1),(LsuPlugin_logic_flushPort_valid && 1'b1)}}}}}});
  assign toplevel_execute_lane1_ctrls_0_downIsCancel = 1'b0;
  assign toplevel_execute_lane1_ctrls_0_upIsCancel = when_ExecuteLanePlugin_l300_5;
  assign when_ExecuteLanePlugin_l300_6 = (|{(late1_BranchPlugin_logic_flushPort_valid && 1'b1),{(early1_BranchPlugin_logic_flushPort_valid && 1'b1),{(late0_BranchPlugin_logic_flushPort_valid && 1'b1),{(early0_EnvPlugin_logic_flushPort_valid && 1'b1),{(CsrAccessPlugin_logic_flushPort_valid && 1'b1),{(early0_BranchPlugin_logic_flushPort_valid && 1'b1),(LsuPlugin_logic_flushPort_valid && 1'b1)}}}}}});
  assign toplevel_execute_lane1_ctrls_1_downIsCancel = 1'b0;
  assign toplevel_execute_lane1_ctrls_1_upIsCancel = when_ExecuteLanePlugin_l300_6;
  assign when_ExecuteLanePlugin_l300_7 = (|{(late1_BranchPlugin_logic_flushPort_valid && 1'b1),{(early1_BranchPlugin_logic_flushPort_valid && 1'b1),{(late0_BranchPlugin_logic_flushPort_valid && 1'b1),{((early0_EnvPlugin_logic_flushPort_valid && 1'b1) && ((early0_EnvPlugin_logic_flushPort_payload_laneAge < toplevel_execute_ctrl2_down_LANE_AGE_lane1) || (_zz_when_ExecuteLanePlugin_l300_7 && early0_EnvPlugin_logic_flushPort_payload_self))),{((CsrAccessPlugin_logic_flushPort_valid && _zz_when_ExecuteLanePlugin_l300_7_1) && (_zz_when_ExecuteLanePlugin_l300_7_2 || _zz_when_ExecuteLanePlugin_l300_7_3)),{(early0_BranchPlugin_logic_flushPort_valid && _zz_when_ExecuteLanePlugin_l300_7_4),(LsuPlugin_logic_flushPort_valid && _zz_when_ExecuteLanePlugin_l300_7_5)}}}}}});
  assign toplevel_execute_lane1_ctrls_2_downIsCancel = 1'b0;
  assign toplevel_execute_lane1_ctrls_2_upIsCancel = when_ExecuteLanePlugin_l300_7;
  assign when_ExecuteLanePlugin_l300_8 = (|{(late1_BranchPlugin_logic_flushPort_valid && 1'b1),{((early1_BranchPlugin_logic_flushPort_valid && 1'b1) && ((early1_BranchPlugin_logic_flushPort_payload_laneAge < toplevel_execute_ctrl3_down_LANE_AGE_lane1) || ((early1_BranchPlugin_logic_flushPort_payload_laneAge == toplevel_execute_ctrl3_down_LANE_AGE_lane1) && early1_BranchPlugin_logic_flushPort_payload_self))),{(late0_BranchPlugin_logic_flushPort_valid && 1'b1),{((early0_BranchPlugin_logic_flushPort_valid && _zz_when_ExecuteLanePlugin_l300_8) && (_zz_when_ExecuteLanePlugin_l300_8_1 || _zz_when_ExecuteLanePlugin_l300_8_2)),(LsuPlugin_logic_flushPort_valid && 1'b1)}}}});
  assign toplevel_execute_lane1_ctrls_3_downIsCancel = 1'b0;
  assign toplevel_execute_lane1_ctrls_3_upIsCancel = when_ExecuteLanePlugin_l300_8;
  assign when_ExecuteLanePlugin_l300_9 = (|{((late1_BranchPlugin_logic_flushPort_valid && 1'b1) && ((late1_BranchPlugin_logic_flushPort_payload_laneAge < toplevel_execute_ctrl4_down_LANE_AGE_lane1) || ((late1_BranchPlugin_logic_flushPort_payload_laneAge == toplevel_execute_ctrl4_down_LANE_AGE_lane1) && late1_BranchPlugin_logic_flushPort_payload_self))),{((late0_BranchPlugin_logic_flushPort_valid && 1'b1) && ((late0_BranchPlugin_logic_flushPort_payload_laneAge < toplevel_execute_ctrl4_down_LANE_AGE_lane1) || (_zz_when_ExecuteLanePlugin_l300_9 && late0_BranchPlugin_logic_flushPort_payload_self))),((LsuPlugin_logic_flushPort_valid && 1'b1) && ((LsuPlugin_logic_flushPort_payload_laneAge < toplevel_execute_ctrl4_down_LANE_AGE_lane1) || (_zz_when_ExecuteLanePlugin_l300_9_1 && LsuPlugin_logic_flushPort_payload_self)))}});
  assign toplevel_execute_lane1_ctrls_4_downIsCancel = 1'b0;
  assign toplevel_execute_lane1_ctrls_4_upIsCancel = when_ExecuteLanePlugin_l300_9;
  assign toplevel_execute_lane1_ctrls_5_downIsCancel = 1'b0;
  assign toplevel_execute_lane1_ctrls_5_upIsCancel = 1'b0;
  assign execute_lane1_logic_trapPending[0] = (|{((toplevel_execute_ctrl4_up_LANE_SEL_lane1 && 1'b1) && toplevel_execute_ctrl4_down_TRAP_lane1),{((toplevel_execute_ctrl3_up_LANE_SEL_lane1 && 1'b1) && toplevel_execute_ctrl3_down_TRAP_lane1),{((toplevel_execute_ctrl2_up_LANE_SEL_lane1 && 1'b1) && toplevel_execute_ctrl2_down_TRAP_lane1),((toplevel_execute_ctrl1_up_LANE_SEL_lane1 && 1'b1) && toplevel_execute_ctrl1_down_TRAP_lane1)}}});
  assign toplevel_execute_ctrl2_up_COMMIT_lane1 = (! toplevel_execute_ctrl2_up_TRAP_lane1);
  assign integer_RegFilePlugin_logic_writeMerges_0_bus_valid = (|lane0_integer_WriteBackPlugin_logic_write_port_valid);
  assign integer_RegFilePlugin_logic_writeMerges_0_bus_address = lane0_integer_WriteBackPlugin_logic_write_port_address;
  assign integer_RegFilePlugin_logic_writeMerges_0_bus_data = lane0_integer_WriteBackPlugin_logic_write_port_data;
  assign integer_RegFilePlugin_logic_writeMerges_0_bus_uopId = lane0_integer_WriteBackPlugin_logic_write_port_uopId;
  assign integer_RegFilePlugin_logic_writeMerges_1_bus_valid = (|lane1_integer_WriteBackPlugin_logic_write_port_valid);
  assign integer_RegFilePlugin_logic_writeMerges_1_bus_address = lane1_integer_WriteBackPlugin_logic_write_port_address;
  assign integer_RegFilePlugin_logic_writeMerges_1_bus_data = lane1_integer_WriteBackPlugin_logic_write_port_data;
  assign integer_RegFilePlugin_logic_writeMerges_1_bus_uopId = lane1_integer_WriteBackPlugin_logic_write_port_uopId;
  assign toplevel_execute_lane1_bypasser_integer_RS1_port_data = integer_RegFilePlugin_logic_regfile_fpga_io_reads_0_data;
  assign toplevel_execute_lane0_bypasser_integer_RS1_port_data = integer_RegFilePlugin_logic_regfile_fpga_io_reads_1_data;
  assign toplevel_execute_lane0_bypasser_integer_RS2_port_data = integer_RegFilePlugin_logic_regfile_fpga_io_reads_2_data;
  assign toplevel_execute_lane1_bypasser_integer_RS2_port_data = integer_RegFilePlugin_logic_regfile_fpga_io_reads_3_data;
  always @(*) begin
    integer_RegFilePlugin_logic_regfile_fpga_io_writes_0_valid = integer_RegFilePlugin_logic_writeMerges_0_bus_valid;
    if(when_RegFilePlugin_l127) begin
      integer_RegFilePlugin_logic_regfile_fpga_io_writes_0_valid = 1'b1;
    end
  end

  always @(*) begin
    integer_RegFilePlugin_logic_regfile_fpga_io_writes_0_address = integer_RegFilePlugin_logic_writeMerges_0_bus_address;
    if(when_RegFilePlugin_l127) begin
      integer_RegFilePlugin_logic_regfile_fpga_io_writes_0_address = integer_RegFilePlugin_logic_initalizer_counter[4:0];
    end
  end

  always @(*) begin
    integer_RegFilePlugin_logic_regfile_fpga_io_writes_0_data = integer_RegFilePlugin_logic_writeMerges_0_bus_data;
    if(when_RegFilePlugin_l127) begin
      integer_RegFilePlugin_logic_regfile_fpga_io_writes_0_data = 32'h0;
    end
  end

  assign integer_RegFilePlugin_logic_initalizer_done = integer_RegFilePlugin_logic_initalizer_counter[5];
  assign when_RegFilePlugin_l127 = (! integer_RegFilePlugin_logic_initalizer_done);
  assign integer_write_0_valid = integer_RegFilePlugin_logic_writeMerges_0_bus_valid;
  assign integer_write_0_address = integer_RegFilePlugin_logic_writeMerges_0_bus_address;
  assign integer_write_0_data = integer_RegFilePlugin_logic_writeMerges_0_bus_data;
  assign integer_write_0_uopId = integer_RegFilePlugin_logic_writeMerges_0_bus_uopId;
  assign integer_write_1_valid = integer_RegFilePlugin_logic_writeMerges_1_bus_valid;
  assign integer_write_1_address = integer_RegFilePlugin_logic_writeMerges_1_bus_address;
  assign integer_write_1_data = integer_RegFilePlugin_logic_writeMerges_1_bus_data;
  assign integer_write_1_uopId = integer_RegFilePlugin_logic_writeMerges_1_bus_uopId;
  assign execute_freeze_valid = (|{CsrAccessPlugin_logic_fsm_inject_iLogic_freeze,{LsuPlugin_logic_onCtrl_rva_freezeIt,{LsuPlugin_logic_onCtrl_io_freezeIt,{early0_DivPlugin_logic_processing_freeze,((toplevel_execute_ctrl4_up_LANE_SEL_lane0 && toplevel_execute_ctrl4_down_MulPlugin_HIGH_lane0) && (! early0_MulPlugin_logic_writeback_buffer_valid))}}}});
  assign toplevel_execute_ctrl5_down_ready = (! execute_freeze_valid);
  assign FetchL1Plugin_pmaBuilder_addressBits = FetchL1Plugin_logic_ctrl_pmaPort_cmd_address;
  assign _zz_FetchL1Plugin_logic_ctrl_pmaPort_rsp_io = ((FetchL1Plugin_pmaBuilder_addressBits & 32'h0) == 32'h0);
  assign FetchL1Plugin_pmaBuilder_onTransfers_0_addressHit = _zz_FetchL1Plugin_pmaBuilder_onTransfers_0_addressHit[0];
  assign FetchL1Plugin_pmaBuilder_onTransfers_0_argsHit = (|1'b1);
  assign FetchL1Plugin_pmaBuilder_onTransfers_0_hit = (FetchL1Plugin_pmaBuilder_onTransfers_0_argsHit && FetchL1Plugin_pmaBuilder_onTransfers_0_addressHit);
  assign FetchL1Plugin_logic_ctrl_pmaPort_rsp_fault = (! ((|{((FetchL1Plugin_pmaBuilder_addressBits & 32'hf8000000) == 32'h80000000),((FetchL1Plugin_pmaBuilder_addressBits & 32'hffffc000) == 32'h40000000)}) && (|FetchL1Plugin_pmaBuilder_onTransfers_0_hit)));
  assign FetchL1Plugin_logic_ctrl_pmaPort_rsp_io = (! _zz_FetchL1Plugin_logic_ctrl_pmaPort_rsp_io_1[0]);
  assign LsuPlugin_pmaBuilder_l1_addressBits = LsuPlugin_logic_onPma_cached_cmd_address;
  assign LsuPlugin_pmaBuilder_l1_argsBits = LsuPlugin_logic_onPma_cached_cmd_op;
  assign _zz_LsuPlugin_logic_onPma_cached_rsp_io = ((LsuPlugin_pmaBuilder_l1_addressBits & 32'h0) == 32'h0);
  assign LsuPlugin_pmaBuilder_l1_onTransfers_0_addressHit = _zz_LsuPlugin_pmaBuilder_l1_onTransfers_0_addressHit[0];
  assign LsuPlugin_pmaBuilder_l1_onTransfers_0_argsHit = (|((LsuPlugin_pmaBuilder_l1_argsBits & 1'b0) == 1'b0));
  assign LsuPlugin_pmaBuilder_l1_onTransfers_0_hit = (LsuPlugin_pmaBuilder_l1_onTransfers_0_argsHit && LsuPlugin_pmaBuilder_l1_onTransfers_0_addressHit);
  assign LsuPlugin_logic_onPma_cached_rsp_fault = (! ((|{((LsuPlugin_pmaBuilder_l1_addressBits & 32'hf8000000) == 32'h80000000),((LsuPlugin_pmaBuilder_l1_addressBits & 32'hffffc000) == 32'h40000000)}) && (|LsuPlugin_pmaBuilder_l1_onTransfers_0_hit)));
  assign LsuPlugin_logic_onPma_cached_rsp_io = (! _zz_LsuPlugin_logic_onPma_cached_rsp_io_1[0]);
  assign LsuPlugin_pmaBuilder_io_addressBits = LsuPlugin_logic_onPma_io_cmd_address;
  assign LsuPlugin_pmaBuilder_io_argsBits = {LsuPlugin_logic_onPma_io_cmd_size,LsuPlugin_logic_onPma_io_cmd_op};
  assign LsuPlugin_pmaBuilder_io_onTransfers_0_addressHit = _zz_LsuPlugin_pmaBuilder_io_onTransfers_0_addressHit[0];
  assign LsuPlugin_pmaBuilder_io_onTransfers_0_argsHit = (|{((LsuPlugin_pmaBuilder_io_argsBits & 3'b100) == 3'b100),((LsuPlugin_pmaBuilder_io_argsBits & 3'b001) == 3'b000)});
  assign LsuPlugin_pmaBuilder_io_onTransfers_0_hit = (LsuPlugin_pmaBuilder_io_onTransfers_0_argsHit && LsuPlugin_pmaBuilder_io_onTransfers_0_addressHit);
  assign _zz_LsuPlugin_logic_onPma_io_rsp_io = ((LsuPlugin_pmaBuilder_io_addressBits & 32'h80000000) == 32'h80000000);
  assign _zz_LsuPlugin_logic_onPma_io_rsp_io_1 = ((LsuPlugin_pmaBuilder_io_addressBits & 32'h40000000) == 32'h40000000);
  assign LsuPlugin_pmaBuilder_io_onTransfers_1_addressHit = _zz_LsuPlugin_pmaBuilder_io_onTransfers_1_addressHit[0];
  assign LsuPlugin_pmaBuilder_io_onTransfers_1_argsHit = (|((LsuPlugin_pmaBuilder_io_argsBits & 3'b000) == 3'b000));
  assign LsuPlugin_pmaBuilder_io_onTransfers_1_hit = (LsuPlugin_pmaBuilder_io_onTransfers_1_argsHit && LsuPlugin_pmaBuilder_io_onTransfers_1_addressHit);
  assign LsuPlugin_logic_onPma_io_rsp_fault = (! ((|{((LsuPlugin_pmaBuilder_io_addressBits & 32'h78000000) == 32'h0),((LsuPlugin_pmaBuilder_io_addressBits & 32'hffffc000) == 32'h40000000)}) && (|{LsuPlugin_pmaBuilder_io_onTransfers_1_hit,LsuPlugin_pmaBuilder_io_onTransfers_0_hit})));
  assign LsuPlugin_logic_onPma_io_rsp_io = (! _zz_LsuPlugin_logic_onPma_io_rsp_io_2[0]);
  assign WhiteboxerPlugin_logic_completions_ports_5_valid = execute_lane1_logic_completions_onCtrl_0_port_valid;
  assign WhiteboxerPlugin_logic_completions_ports_5_payload_uopId = execute_lane1_logic_completions_onCtrl_0_port_payload_uopId;
  assign WhiteboxerPlugin_logic_completions_ports_5_payload_trap = execute_lane1_logic_completions_onCtrl_0_port_payload_trap;
  assign WhiteboxerPlugin_logic_completions_ports_5_payload_commit = execute_lane1_logic_completions_onCtrl_0_port_payload_commit;
  assign WhiteboxerPlugin_logic_completions_ports_6_valid = execute_lane1_logic_completions_onCtrl_1_port_valid;
  assign WhiteboxerPlugin_logic_completions_ports_6_payload_uopId = execute_lane1_logic_completions_onCtrl_1_port_payload_uopId;
  assign WhiteboxerPlugin_logic_completions_ports_6_payload_trap = execute_lane1_logic_completions_onCtrl_1_port_payload_trap;
  assign WhiteboxerPlugin_logic_completions_ports_6_payload_commit = execute_lane1_logic_completions_onCtrl_1_port_payload_commit;
  assign WhiteboxerPlugin_logic_completions_ports_7_valid = execute_lane1_logic_completions_onCtrl_2_port_valid;
  assign WhiteboxerPlugin_logic_completions_ports_7_payload_uopId = execute_lane1_logic_completions_onCtrl_2_port_payload_uopId;
  assign WhiteboxerPlugin_logic_completions_ports_7_payload_trap = execute_lane1_logic_completions_onCtrl_2_port_payload_trap;
  assign WhiteboxerPlugin_logic_completions_ports_7_payload_commit = execute_lane1_logic_completions_onCtrl_2_port_payload_commit;
  assign WhiteboxerPlugin_logic_commits_ports_0_oh_0 = ((((toplevel_execute_ctrl4_down_LANE_SEL_lane0 && toplevel_execute_ctrl4_down_isReady) && (! toplevel_execute_lane0_ctrls_4_downIsCancel)) && toplevel_execute_ctrl4_down_COMMIT_lane0) && (toplevel_execute_ctrl4_down_LANE_AGE_lane0 == 1'b0));
  assign WhiteboxerPlugin_logic_commits_ports_0_oh_1 = ((((toplevel_execute_ctrl4_down_LANE_SEL_lane1 && toplevel_execute_ctrl4_down_isReady) && (! toplevel_execute_lane1_ctrls_4_downIsCancel)) && toplevel_execute_ctrl4_down_COMMIT_lane1) && (toplevel_execute_ctrl4_down_LANE_AGE_lane1 == 1'b0));
  assign WhiteboxerPlugin_logic_commits_ports_0_valid = (|{WhiteboxerPlugin_logic_commits_ports_0_oh_1,WhiteboxerPlugin_logic_commits_ports_0_oh_0});
  assign WhiteboxerPlugin_logic_commits_ports_0_pc = ((WhiteboxerPlugin_logic_commits_ports_0_oh_0 ? toplevel_execute_ctrl4_down_PC_lane0 : 32'h0) | (WhiteboxerPlugin_logic_commits_ports_0_oh_1 ? toplevel_execute_ctrl4_down_PC_lane1 : 32'h0));
  assign WhiteboxerPlugin_logic_commits_ports_0_uop = ((WhiteboxerPlugin_logic_commits_ports_0_oh_0 ? toplevel_execute_ctrl4_down_Decode_UOP_lane0 : 32'h0) | (WhiteboxerPlugin_logic_commits_ports_0_oh_1 ? toplevel_execute_ctrl4_down_Decode_UOP_lane1 : 32'h0));
  assign WhiteboxerPlugin_logic_commits_ports_1_oh_0 = ((((toplevel_execute_ctrl4_down_LANE_SEL_lane0 && toplevel_execute_ctrl4_down_isReady) && (! toplevel_execute_lane0_ctrls_4_downIsCancel)) && toplevel_execute_ctrl4_down_COMMIT_lane0) && (toplevel_execute_ctrl4_down_LANE_AGE_lane0 == 1'b1));
  assign WhiteboxerPlugin_logic_commits_ports_1_oh_1 = ((((toplevel_execute_ctrl4_down_LANE_SEL_lane1 && toplevel_execute_ctrl4_down_isReady) && (! toplevel_execute_lane1_ctrls_4_downIsCancel)) && toplevel_execute_ctrl4_down_COMMIT_lane1) && (toplevel_execute_ctrl4_down_LANE_AGE_lane1 == 1'b1));
  assign WhiteboxerPlugin_logic_commits_ports_1_valid = (|{WhiteboxerPlugin_logic_commits_ports_1_oh_1,WhiteboxerPlugin_logic_commits_ports_1_oh_0});
  assign WhiteboxerPlugin_logic_commits_ports_1_pc = ((WhiteboxerPlugin_logic_commits_ports_1_oh_0 ? toplevel_execute_ctrl4_down_PC_lane0 : 32'h0) | (WhiteboxerPlugin_logic_commits_ports_1_oh_1 ? toplevel_execute_ctrl4_down_PC_lane1 : 32'h0));
  assign WhiteboxerPlugin_logic_commits_ports_1_uop = ((WhiteboxerPlugin_logic_commits_ports_1_oh_0 ? toplevel_execute_ctrl4_down_Decode_UOP_lane0 : 32'h0) | (WhiteboxerPlugin_logic_commits_ports_1_oh_1 ? toplevel_execute_ctrl4_down_Decode_UOP_lane1 : 32'h0));
  assign WhiteboxerPlugin_logic_reschedules_flushes_0_valid = BtbPlugin_logic_flushPort_valid;
  assign WhiteboxerPlugin_logic_reschedules_flushes_0_payload_self = BtbPlugin_logic_flushPort_payload_self;
  assign WhiteboxerPlugin_logic_reschedules_flushes_1_valid = LsuPlugin_logic_flushPort_valid;
  assign WhiteboxerPlugin_logic_reschedules_flushes_1_payload_uopId = LsuPlugin_logic_flushPort_payload_uopId;
  assign WhiteboxerPlugin_logic_reschedules_flushes_1_payload_laneAge = LsuPlugin_logic_flushPort_payload_laneAge;
  assign WhiteboxerPlugin_logic_reschedules_flushes_1_payload_self = LsuPlugin_logic_flushPort_payload_self;
  assign WhiteboxerPlugin_logic_reschedules_flushes_2_valid = early0_BranchPlugin_logic_flushPort_valid;
  assign WhiteboxerPlugin_logic_reschedules_flushes_2_payload_uopId = early0_BranchPlugin_logic_flushPort_payload_uopId;
  assign WhiteboxerPlugin_logic_reschedules_flushes_2_payload_laneAge = early0_BranchPlugin_logic_flushPort_payload_laneAge;
  assign WhiteboxerPlugin_logic_reschedules_flushes_2_payload_self = early0_BranchPlugin_logic_flushPort_payload_self;
  assign WhiteboxerPlugin_logic_reschedules_flushes_3_valid = CsrAccessPlugin_logic_flushPort_valid;
  assign WhiteboxerPlugin_logic_reschedules_flushes_3_payload_uopId = CsrAccessPlugin_logic_flushPort_payload_uopId;
  assign WhiteboxerPlugin_logic_reschedules_flushes_3_payload_laneAge = CsrAccessPlugin_logic_flushPort_payload_laneAge;
  assign WhiteboxerPlugin_logic_reschedules_flushes_3_payload_self = CsrAccessPlugin_logic_flushPort_payload_self;
  assign WhiteboxerPlugin_logic_reschedules_flushes_4_valid = early0_EnvPlugin_logic_flushPort_valid;
  assign WhiteboxerPlugin_logic_reschedules_flushes_4_payload_uopId = early0_EnvPlugin_logic_flushPort_payload_uopId;
  assign WhiteboxerPlugin_logic_reschedules_flushes_4_payload_laneAge = early0_EnvPlugin_logic_flushPort_payload_laneAge;
  assign WhiteboxerPlugin_logic_reschedules_flushes_4_payload_self = early0_EnvPlugin_logic_flushPort_payload_self;
  assign WhiteboxerPlugin_logic_reschedules_flushes_5_valid = late0_BranchPlugin_logic_flushPort_valid;
  assign WhiteboxerPlugin_logic_reschedules_flushes_5_payload_uopId = late0_BranchPlugin_logic_flushPort_payload_uopId;
  assign WhiteboxerPlugin_logic_reschedules_flushes_5_payload_laneAge = late0_BranchPlugin_logic_flushPort_payload_laneAge;
  assign WhiteboxerPlugin_logic_reschedules_flushes_5_payload_self = late0_BranchPlugin_logic_flushPort_payload_self;
  assign WhiteboxerPlugin_logic_reschedules_flushes_6_valid = early1_BranchPlugin_logic_flushPort_valid;
  assign WhiteboxerPlugin_logic_reschedules_flushes_6_payload_uopId = early1_BranchPlugin_logic_flushPort_payload_uopId;
  assign WhiteboxerPlugin_logic_reschedules_flushes_6_payload_laneAge = early1_BranchPlugin_logic_flushPort_payload_laneAge;
  assign WhiteboxerPlugin_logic_reschedules_flushes_6_payload_self = early1_BranchPlugin_logic_flushPort_payload_self;
  assign WhiteboxerPlugin_logic_reschedules_flushes_7_valid = late1_BranchPlugin_logic_flushPort_valid;
  assign WhiteboxerPlugin_logic_reschedules_flushes_7_payload_uopId = late1_BranchPlugin_logic_flushPort_payload_uopId;
  assign WhiteboxerPlugin_logic_reschedules_flushes_7_payload_laneAge = late1_BranchPlugin_logic_flushPort_payload_laneAge;
  assign WhiteboxerPlugin_logic_reschedules_flushes_7_payload_self = late1_BranchPlugin_logic_flushPort_payload_self;
  assign WhiteboxerPlugin_logic_reschedules_flushes_8_valid = DecoderPlugin_logic_laneLogic_0_flushPort_valid;
  assign WhiteboxerPlugin_logic_reschedules_flushes_8_payload_uopId = DecoderPlugin_logic_laneLogic_0_flushPort_payload_uopId;
  assign WhiteboxerPlugin_logic_reschedules_flushes_8_payload_laneAge = DecoderPlugin_logic_laneLogic_0_flushPort_payload_laneAge;
  assign WhiteboxerPlugin_logic_reschedules_flushes_8_payload_self = DecoderPlugin_logic_laneLogic_0_flushPort_payload_self;
  assign WhiteboxerPlugin_logic_reschedules_flushes_9_valid = DecoderPlugin_logic_laneLogic_1_flushPort_valid;
  assign WhiteboxerPlugin_logic_reschedules_flushes_9_payload_uopId = DecoderPlugin_logic_laneLogic_1_flushPort_payload_uopId;
  assign WhiteboxerPlugin_logic_reschedules_flushes_9_payload_laneAge = DecoderPlugin_logic_laneLogic_1_flushPort_payload_laneAge;
  assign WhiteboxerPlugin_logic_reschedules_flushes_9_payload_self = DecoderPlugin_logic_laneLogic_1_flushPort_payload_self;
  assign WhiteboxerPlugin_logic_prediction_learns_0_valid = late0_BranchPlugin_logic_jumpLogic_learn_valid;
  assign WhiteboxerPlugin_logic_prediction_learns_0_payload_pcOnLastSlice = late0_BranchPlugin_logic_jumpLogic_learn_payload_pcOnLastSlice;
  assign WhiteboxerPlugin_logic_prediction_learns_0_payload_pcTarget = late0_BranchPlugin_logic_jumpLogic_learn_payload_pcTarget;
  assign WhiteboxerPlugin_logic_prediction_learns_0_payload_taken = late0_BranchPlugin_logic_jumpLogic_learn_payload_taken;
  assign WhiteboxerPlugin_logic_prediction_learns_0_payload_isBranch = late0_BranchPlugin_logic_jumpLogic_learn_payload_isBranch;
  assign WhiteboxerPlugin_logic_prediction_learns_0_payload_isPush = late0_BranchPlugin_logic_jumpLogic_learn_payload_isPush;
  assign WhiteboxerPlugin_logic_prediction_learns_0_payload_isPop = late0_BranchPlugin_logic_jumpLogic_learn_payload_isPop;
  assign WhiteboxerPlugin_logic_prediction_learns_0_payload_wasWrong = late0_BranchPlugin_logic_jumpLogic_learn_payload_wasWrong;
  assign WhiteboxerPlugin_logic_prediction_learns_0_payload_badPredictedTarget = late0_BranchPlugin_logic_jumpLogic_learn_payload_badPredictedTarget;
  assign WhiteboxerPlugin_logic_prediction_learns_0_payload_history = late0_BranchPlugin_logic_jumpLogic_learn_payload_history;
  assign WhiteboxerPlugin_logic_prediction_learns_0_payload_uopId = late0_BranchPlugin_logic_jumpLogic_learn_payload_uopId;
  assign WhiteboxerPlugin_logic_prediction_learns_0_payload_ctx_GSharePlugin_GSHARE_COUNTER_0 = late0_BranchPlugin_logic_jumpLogic_learn_payload_ctx_GSharePlugin_GSHARE_COUNTER_0;
  assign WhiteboxerPlugin_logic_prediction_learns_0_payload_ctx_GSharePlugin_GSHARE_COUNTER_1 = late0_BranchPlugin_logic_jumpLogic_learn_payload_ctx_GSharePlugin_GSHARE_COUNTER_1;
  assign WhiteboxerPlugin_logic_prediction_learns_0_payload_ctx_GSharePlugin_GSHARE_COUNTER_2 = late0_BranchPlugin_logic_jumpLogic_learn_payload_ctx_GSharePlugin_GSHARE_COUNTER_2;
  assign WhiteboxerPlugin_logic_prediction_learns_0_payload_ctx_GSharePlugin_GSHARE_COUNTER_3 = late0_BranchPlugin_logic_jumpLogic_learn_payload_ctx_GSharePlugin_GSHARE_COUNTER_3;
  assign WhiteboxerPlugin_logic_prediction_learns_1_valid = late1_BranchPlugin_logic_jumpLogic_learn_valid;
  assign WhiteboxerPlugin_logic_prediction_learns_1_payload_pcOnLastSlice = late1_BranchPlugin_logic_jumpLogic_learn_payload_pcOnLastSlice;
  assign WhiteboxerPlugin_logic_prediction_learns_1_payload_pcTarget = late1_BranchPlugin_logic_jumpLogic_learn_payload_pcTarget;
  assign WhiteboxerPlugin_logic_prediction_learns_1_payload_taken = late1_BranchPlugin_logic_jumpLogic_learn_payload_taken;
  assign WhiteboxerPlugin_logic_prediction_learns_1_payload_isBranch = late1_BranchPlugin_logic_jumpLogic_learn_payload_isBranch;
  assign WhiteboxerPlugin_logic_prediction_learns_1_payload_isPush = late1_BranchPlugin_logic_jumpLogic_learn_payload_isPush;
  assign WhiteboxerPlugin_logic_prediction_learns_1_payload_isPop = late1_BranchPlugin_logic_jumpLogic_learn_payload_isPop;
  assign WhiteboxerPlugin_logic_prediction_learns_1_payload_wasWrong = late1_BranchPlugin_logic_jumpLogic_learn_payload_wasWrong;
  assign WhiteboxerPlugin_logic_prediction_learns_1_payload_badPredictedTarget = late1_BranchPlugin_logic_jumpLogic_learn_payload_badPredictedTarget;
  assign WhiteboxerPlugin_logic_prediction_learns_1_payload_history = late1_BranchPlugin_logic_jumpLogic_learn_payload_history;
  assign WhiteboxerPlugin_logic_prediction_learns_1_payload_uopId = late1_BranchPlugin_logic_jumpLogic_learn_payload_uopId;
  assign WhiteboxerPlugin_logic_prediction_learns_1_payload_ctx_GSharePlugin_GSHARE_COUNTER_0 = late1_BranchPlugin_logic_jumpLogic_learn_payload_ctx_GSharePlugin_GSHARE_COUNTER_0;
  assign WhiteboxerPlugin_logic_prediction_learns_1_payload_ctx_GSharePlugin_GSHARE_COUNTER_1 = late1_BranchPlugin_logic_jumpLogic_learn_payload_ctx_GSharePlugin_GSHARE_COUNTER_1;
  assign WhiteboxerPlugin_logic_prediction_learns_1_payload_ctx_GSharePlugin_GSHARE_COUNTER_2 = late1_BranchPlugin_logic_jumpLogic_learn_payload_ctx_GSharePlugin_GSHARE_COUNTER_2;
  assign WhiteboxerPlugin_logic_prediction_learns_1_payload_ctx_GSharePlugin_GSHARE_COUNTER_3 = late1_BranchPlugin_logic_jumpLogic_learn_payload_ctx_GSharePlugin_GSHARE_COUNTER_3;
  assign WhiteboxerPlugin_logic_loadExecute_fire = (((((((toplevel_execute_ctrl4_down_LANE_SEL_lane0 && toplevel_execute_ctrl4_down_isReady) && (! toplevel_execute_lane0_ctrls_4_downIsCancel)) && toplevel_execute_ctrl4_down_AguPlugin_SEL_lane0) && toplevel_execute_ctrl4_down_AguPlugin_LOAD_lane0) && (! toplevel_execute_ctrl4_down_LsuPlugin_logic_LSU_PREFETCH_lane0)) && (! toplevel_execute_ctrl4_down_TRAP_lane0)) && (! toplevel_execute_ctrl4_down_LsuPlugin_logic_onPma_IO_lane0));
  assign WhiteboxerPlugin_logic_loadExecute_uopId = toplevel_execute_ctrl4_down_Decode_UOP_ID_lane0;
  assign WhiteboxerPlugin_logic_loadExecute_size = toplevel_execute_ctrl4_down_AguPlugin_SIZE_lane0;
  assign WhiteboxerPlugin_logic_loadExecute_address = toplevel_execute_ctrl4_down_LsuL1_PHYSICAL_ADDRESS_lane0;
  assign WhiteboxerPlugin_logic_loadExecute_data = lane0_IntFormatPlugin_logic_stages_2_wb_payload;
  assign WhiteboxerPlugin_logic_storeCommit_fire = LsuPlugin_logic_onWb_storeFire;
  assign WhiteboxerPlugin_logic_storeCommit_uopId = toplevel_execute_ctrl4_down_Decode_UOP_ID_lane0;
  assign WhiteboxerPlugin_logic_storeCommit_size = toplevel_execute_ctrl4_down_AguPlugin_SIZE_lane0;
  assign WhiteboxerPlugin_logic_storeCommit_address = toplevel_execute_ctrl4_down_MMU_TRANSLATED_lane0;
  assign WhiteboxerPlugin_logic_storeCommit_data = toplevel_execute_ctrl4_down_LsuL1_WRITE_DATA_lane0;
  assign WhiteboxerPlugin_logic_storeCommit_storeId = toplevel_execute_ctrl4_down_Decode_STORE_ID_lane0;
  assign WhiteboxerPlugin_logic_storeCommit_amo = 1'b0;
  assign WhiteboxerPlugin_logic_storeConditional_fire = (((((toplevel_execute_ctrl4_down_LANE_SEL_lane0 && toplevel_execute_ctrl4_down_isReady) && (! toplevel_execute_lane0_ctrls_4_downIsCancel)) && toplevel_execute_ctrl4_down_AguPlugin_SEL_lane0) && (toplevel_execute_ctrl4_down_AguPlugin_ATOMIC_lane0 && (! toplevel_execute_ctrl4_down_AguPlugin_LOAD_lane0))) && (! toplevel_execute_ctrl4_down_TRAP_lane0));
  assign WhiteboxerPlugin_logic_storeConditional_uopId = toplevel_execute_ctrl4_down_Decode_UOP_ID_lane0;
  assign WhiteboxerPlugin_logic_storeConditional_miss = toplevel_execute_ctrl4_down_LsuPlugin_logic_onCtrl_SC_MISS_lane0;
  assign WhiteboxerPlugin_logic_storeBroadcast_fire = LsuPlugin_logic_onWb_storeBroadcast;
  assign WhiteboxerPlugin_logic_storeBroadcast_storeId = toplevel_execute_ctrl4_down_Decode_STORE_ID_lane0;
  assign TrapPlugin_logic_initHold = (|{(! CsrRamPlugin_logic_flush_done),{((! LsuL1Plugin_logic_initializer_done) || LsuL1Plugin_logic_initializerMem_busy),{(! integer_RegFilePlugin_logic_initalizer_done),{(FetchL1Plugin_logic_invalidate_firstEver || FetchL1Plugin_logic_initializer_busy),{GSharePlugin_logic_initializer_busy,BtbPlugin_logic_initializer_busy}}}}});
  assign WhiteboxerPlugin_logic_wfi = TrapPlugin_logic_harts_0_trap_fsm_wfi;
  assign WhiteboxerPlugin_logic_perf_executeFreezed = execute_freeze_valid;
  assign WhiteboxerPlugin_logic_perf_dispatchHazards = (|{(DispatchPlugin_logic_candidates_2_ctx_valid && (! DispatchPlugin_logic_candidates_2_fire)),{(DispatchPlugin_logic_candidates_1_ctx_valid && (! DispatchPlugin_logic_candidates_1_fire)),(DispatchPlugin_logic_candidates_0_ctx_valid && (! DispatchPlugin_logic_candidates_0_fire))}});
  assign WhiteboxerPlugin_logic_perf_candidatesCount = _zz_WhiteboxerPlugin_logic_perf_candidatesCount;
  assign WhiteboxerPlugin_logic_perf_dispatchFeedCount = _zz_WhiteboxerPlugin_logic_perf_dispatchFeedCount;
  always @(*) begin
    _zz_WhiteboxerPlugin_logic_perf_executeFreezedCounter = 1'b0;
    if(WhiteboxerPlugin_logic_perf_executeFreezed) begin
      _zz_WhiteboxerPlugin_logic_perf_executeFreezedCounter = 1'b1;
    end
  end

  always @(*) begin
    _zz_WhiteboxerPlugin_logic_perf_executeFreezedCounter_1 = (_zz_WhiteboxerPlugin_logic_perf_executeFreezedCounter_2 + _zz__zz_WhiteboxerPlugin_logic_perf_executeFreezedCounter_1);
    if(1'b0) begin
      _zz_WhiteboxerPlugin_logic_perf_executeFreezedCounter_1 = 60'h0;
    end
  end

  assign WhiteboxerPlugin_logic_perf_executeFreezedCounter = _zz_WhiteboxerPlugin_logic_perf_executeFreezedCounter_2;
  always @(*) begin
    _zz_WhiteboxerPlugin_logic_perf_dispatchHazardsCounter = 1'b0;
    if(WhiteboxerPlugin_logic_perf_dispatchHazards) begin
      _zz_WhiteboxerPlugin_logic_perf_dispatchHazardsCounter = 1'b1;
    end
  end

  always @(*) begin
    _zz_WhiteboxerPlugin_logic_perf_dispatchHazardsCounter_1 = (_zz_WhiteboxerPlugin_logic_perf_dispatchHazardsCounter_2 + _zz__zz_WhiteboxerPlugin_logic_perf_dispatchHazardsCounter_1);
    if(1'b0) begin
      _zz_WhiteboxerPlugin_logic_perf_dispatchHazardsCounter_1 = 60'h0;
    end
  end

  assign WhiteboxerPlugin_logic_perf_dispatchHazardsCounter = _zz_WhiteboxerPlugin_logic_perf_dispatchHazardsCounter_2;
  assign when_Utils_l585 = (WhiteboxerPlugin_logic_perf_candidatesCount == 2'b00);
  always @(*) begin
    _zz_WhiteboxerPlugin_logic_perf_candidatesCountCounters_0 = 1'b0;
    if(when_Utils_l585) begin
      _zz_WhiteboxerPlugin_logic_perf_candidatesCountCounters_0 = 1'b1;
    end
  end

  always @(*) begin
    _zz_WhiteboxerPlugin_logic_perf_candidatesCountCounters_0_1 = (_zz_WhiteboxerPlugin_logic_perf_candidatesCountCounters_0_2 + _zz__zz_WhiteboxerPlugin_logic_perf_candidatesCountCounters_0_1);
    if(1'b0) begin
      _zz_WhiteboxerPlugin_logic_perf_candidatesCountCounters_0_1 = 60'h0;
    end
  end

  assign WhiteboxerPlugin_logic_perf_candidatesCountCounters_0 = _zz_WhiteboxerPlugin_logic_perf_candidatesCountCounters_0_2;
  assign when_Utils_l585_1 = (WhiteboxerPlugin_logic_perf_candidatesCount == 2'b01);
  always @(*) begin
    _zz_WhiteboxerPlugin_logic_perf_candidatesCountCounters_1 = 1'b0;
    if(when_Utils_l585_1) begin
      _zz_WhiteboxerPlugin_logic_perf_candidatesCountCounters_1 = 1'b1;
    end
  end

  always @(*) begin
    _zz_WhiteboxerPlugin_logic_perf_candidatesCountCounters_1_1 = (_zz_WhiteboxerPlugin_logic_perf_candidatesCountCounters_1_2 + _zz__zz_WhiteboxerPlugin_logic_perf_candidatesCountCounters_1_1);
    if(1'b0) begin
      _zz_WhiteboxerPlugin_logic_perf_candidatesCountCounters_1_1 = 60'h0;
    end
  end

  assign WhiteboxerPlugin_logic_perf_candidatesCountCounters_1 = _zz_WhiteboxerPlugin_logic_perf_candidatesCountCounters_1_2;
  assign when_Utils_l585_2 = (WhiteboxerPlugin_logic_perf_candidatesCount == 2'b10);
  always @(*) begin
    _zz_WhiteboxerPlugin_logic_perf_candidatesCountCounters_2 = 1'b0;
    if(when_Utils_l585_2) begin
      _zz_WhiteboxerPlugin_logic_perf_candidatesCountCounters_2 = 1'b1;
    end
  end

  always @(*) begin
    _zz_WhiteboxerPlugin_logic_perf_candidatesCountCounters_2_1 = (_zz_WhiteboxerPlugin_logic_perf_candidatesCountCounters_2_2 + _zz__zz_WhiteboxerPlugin_logic_perf_candidatesCountCounters_2_1);
    if(1'b0) begin
      _zz_WhiteboxerPlugin_logic_perf_candidatesCountCounters_2_1 = 60'h0;
    end
  end

  assign WhiteboxerPlugin_logic_perf_candidatesCountCounters_2 = _zz_WhiteboxerPlugin_logic_perf_candidatesCountCounters_2_2;
  assign when_Utils_l585_3 = (WhiteboxerPlugin_logic_perf_candidatesCount == 2'b11);
  always @(*) begin
    _zz_WhiteboxerPlugin_logic_perf_candidatesCountCounters_3 = 1'b0;
    if(when_Utils_l585_3) begin
      _zz_WhiteboxerPlugin_logic_perf_candidatesCountCounters_3 = 1'b1;
    end
  end

  always @(*) begin
    _zz_WhiteboxerPlugin_logic_perf_candidatesCountCounters_3_1 = (_zz_WhiteboxerPlugin_logic_perf_candidatesCountCounters_3_2 + _zz__zz_WhiteboxerPlugin_logic_perf_candidatesCountCounters_3_1);
    if(1'b0) begin
      _zz_WhiteboxerPlugin_logic_perf_candidatesCountCounters_3_1 = 60'h0;
    end
  end

  assign WhiteboxerPlugin_logic_perf_candidatesCountCounters_3 = _zz_WhiteboxerPlugin_logic_perf_candidatesCountCounters_3_2;
  assign when_Utils_l585_4 = (WhiteboxerPlugin_logic_perf_dispatchFeedCount == 2'b00);
  always @(*) begin
    _zz_WhiteboxerPlugin_logic_perf_dispatchFeedCounters_0 = 1'b0;
    if(when_Utils_l585_4) begin
      _zz_WhiteboxerPlugin_logic_perf_dispatchFeedCounters_0 = 1'b1;
    end
  end

  always @(*) begin
    _zz_WhiteboxerPlugin_logic_perf_dispatchFeedCounters_0_1 = (_zz_WhiteboxerPlugin_logic_perf_dispatchFeedCounters_0_2 + _zz__zz_WhiteboxerPlugin_logic_perf_dispatchFeedCounters_0_1);
    if(1'b0) begin
      _zz_WhiteboxerPlugin_logic_perf_dispatchFeedCounters_0_1 = 60'h0;
    end
  end

  assign WhiteboxerPlugin_logic_perf_dispatchFeedCounters_0 = _zz_WhiteboxerPlugin_logic_perf_dispatchFeedCounters_0_2;
  assign when_Utils_l585_5 = (WhiteboxerPlugin_logic_perf_dispatchFeedCount == 2'b01);
  always @(*) begin
    _zz_WhiteboxerPlugin_logic_perf_dispatchFeedCounters_1 = 1'b0;
    if(when_Utils_l585_5) begin
      _zz_WhiteboxerPlugin_logic_perf_dispatchFeedCounters_1 = 1'b1;
    end
  end

  always @(*) begin
    _zz_WhiteboxerPlugin_logic_perf_dispatchFeedCounters_1_1 = (_zz_WhiteboxerPlugin_logic_perf_dispatchFeedCounters_1_2 + _zz__zz_WhiteboxerPlugin_logic_perf_dispatchFeedCounters_1_1);
    if(1'b0) begin
      _zz_WhiteboxerPlugin_logic_perf_dispatchFeedCounters_1_1 = 60'h0;
    end
  end

  assign WhiteboxerPlugin_logic_perf_dispatchFeedCounters_1 = _zz_WhiteboxerPlugin_logic_perf_dispatchFeedCounters_1_2;
  assign when_Utils_l585_6 = (WhiteboxerPlugin_logic_perf_dispatchFeedCount == 2'b10);
  always @(*) begin
    _zz_WhiteboxerPlugin_logic_perf_dispatchFeedCounters_2 = 1'b0;
    if(when_Utils_l585_6) begin
      _zz_WhiteboxerPlugin_logic_perf_dispatchFeedCounters_2 = 1'b1;
    end
  end

  always @(*) begin
    _zz_WhiteboxerPlugin_logic_perf_dispatchFeedCounters_2_1 = (_zz_WhiteboxerPlugin_logic_perf_dispatchFeedCounters_2_2 + _zz__zz_WhiteboxerPlugin_logic_perf_dispatchFeedCounters_2_1);
    if(1'b0) begin
      _zz_WhiteboxerPlugin_logic_perf_dispatchFeedCounters_2_1 = 60'h0;
    end
  end

  assign WhiteboxerPlugin_logic_perf_dispatchFeedCounters_2 = _zz_WhiteboxerPlugin_logic_perf_dispatchFeedCounters_2_2;
  assign WhiteboxerPlugin_logic_trap_ports_0_valid = TrapPlugin_logic_harts_0_trap_whitebox_trap;
  assign WhiteboxerPlugin_logic_trap_ports_0_interrupt = TrapPlugin_logic_harts_0_trap_whitebox_interrupt;
  assign WhiteboxerPlugin_logic_trap_ports_0_cause = TrapPlugin_logic_harts_0_trap_whitebox_code;
  assign fetch_logic_ctrls_2_up_forgetOne = (|fetch_logic_ctrls_2_forgetsSingleRequest_FetchPipelinePlugin_l46);
  assign fetch_logic_ctrls_2_up_cancel = (|fetch_logic_flushes_1_doIt);
  assign fetch_logic_ctrls_1_up_forgetOne = (|fetch_logic_ctrls_1_throwWhen_FetchPipelinePlugin_l44);
  assign fetch_logic_ctrls_1_up_cancel = (|fetch_logic_ctrls_1_throwWhen_FetchPipelinePlugin_l44);
  assign fetch_logic_ctrls_0_down_ready = fetch_logic_ctrls_1_up_ready;
  assign fetch_logic_ctrls_1_down_ready = fetch_logic_ctrls_2_up_ready;
  always @(*) begin
    fetch_logic_ctrls_0_down_valid = fetch_logic_ctrls_0_up_valid;
    if(when_CtrlLink_l150) begin
      fetch_logic_ctrls_0_down_valid = 1'b0;
    end
  end

  always @(*) begin
    fetch_logic_ctrls_0_up_ready = fetch_logic_ctrls_0_down_isReady;
    if(when_CtrlLink_l150) begin
      fetch_logic_ctrls_0_up_ready = 1'b0;
    end
  end

  assign when_CtrlLink_l150 = (|{fetch_logic_ctrls_0_haltRequest_PcPlugin_l136,{fetch_logic_ctrls_0_haltRequest_BtbPlugin_l171,{fetch_logic_ctrls_0_haltRequest_FetchL1Plugin_l317,fetch_logic_ctrls_0_haltRequest_FetchL1Plugin_l233}}});
  assign fetch_logic_ctrls_0_down_Fetch_WORD_PC = fetch_logic_ctrls_0_up_Fetch_WORD_PC;
  assign fetch_logic_ctrls_0_down_Fetch_PC_FAULT = fetch_logic_ctrls_0_up_Fetch_PC_FAULT;
  assign fetch_logic_ctrls_0_down_Fetch_ID = fetch_logic_ctrls_0_up_Fetch_ID;
  always @(*) begin
    fetch_logic_ctrls_1_down_valid = fetch_logic_ctrls_1_up_valid;
    if(when_CtrlLink_l157) begin
      fetch_logic_ctrls_1_down_valid = 1'b0;
    end
  end

  assign fetch_logic_ctrls_1_up_ready = fetch_logic_ctrls_1_down_isReady;
  assign when_CtrlLink_l157 = (|fetch_logic_ctrls_1_throwWhen_FetchPipelinePlugin_l44);
  assign fetch_logic_ctrls_1_down_Fetch_WORD_PC = fetch_logic_ctrls_1_up_Fetch_WORD_PC;
  assign fetch_logic_ctrls_1_down_Fetch_PC_FAULT = fetch_logic_ctrls_1_up_Fetch_PC_FAULT;
  assign fetch_logic_ctrls_1_down_Fetch_ID = fetch_logic_ctrls_1_up_Fetch_ID;
  assign fetch_logic_ctrls_1_down_FetchL1Plugin_logic_cmd_PLRU_BYPASS_VALID = fetch_logic_ctrls_1_up_FetchL1Plugin_logic_cmd_PLRU_BYPASS_VALID;
  assign fetch_logic_ctrls_1_down_FetchL1Plugin_logic_cmd_PLRU_BYPASS_DATA_0 = fetch_logic_ctrls_1_up_FetchL1Plugin_logic_cmd_PLRU_BYPASS_DATA_0;
  assign fetch_logic_ctrls_1_down_FetchL1Plugin_logic_cmd_TAGS_UPDATE = fetch_logic_ctrls_1_up_FetchL1Plugin_logic_cmd_TAGS_UPDATE;
  assign fetch_logic_ctrls_1_down_FetchL1Plugin_logic_cmd_TAGS_UPDATE_ADDRESS = fetch_logic_ctrls_1_up_FetchL1Plugin_logic_cmd_TAGS_UPDATE_ADDRESS;
  assign fetch_logic_ctrls_1_down_GSharePlugin_logic_HASH = fetch_logic_ctrls_1_up_GSharePlugin_logic_HASH;
  assign fetch_logic_ctrls_1_down_Prediction_BRANCH_HISTORY = fetch_logic_ctrls_1_up_Prediction_BRANCH_HISTORY;
  assign fetch_logic_ctrls_1_down_GSharePlugin_logic_BYPASS_valid = fetch_logic_ctrls_1_up_GSharePlugin_logic_BYPASS_valid;
  assign fetch_logic_ctrls_1_down_GSharePlugin_logic_BYPASS_payload_address = fetch_logic_ctrls_1_up_GSharePlugin_logic_BYPASS_payload_address;
  assign fetch_logic_ctrls_1_down_GSharePlugin_logic_BYPASS_payload_data_0 = fetch_logic_ctrls_1_up_GSharePlugin_logic_BYPASS_payload_data_0;
  assign fetch_logic_ctrls_1_down_GSharePlugin_logic_BYPASS_payload_data_1 = fetch_logic_ctrls_1_up_GSharePlugin_logic_BYPASS_payload_data_1;
  assign fetch_logic_ctrls_1_down_GSharePlugin_logic_BYPASS_payload_data_2 = fetch_logic_ctrls_1_up_GSharePlugin_logic_BYPASS_payload_data_2;
  assign fetch_logic_ctrls_1_down_GSharePlugin_logic_BYPASS_payload_data_3 = fetch_logic_ctrls_1_up_GSharePlugin_logic_BYPASS_payload_data_3;
  assign fetch_logic_ctrls_1_down_BtbPlugin_logic_readCmd_HAZARDS = fetch_logic_ctrls_1_up_BtbPlugin_logic_readCmd_HAZARDS;
  assign fetch_logic_ctrls_2_down_valid = fetch_logic_ctrls_2_up_valid;
  assign fetch_logic_ctrls_2_up_ready = fetch_logic_ctrls_2_down_isReady;
  assign fetch_logic_ctrls_2_down_Fetch_WORD_PC = fetch_logic_ctrls_2_up_Fetch_WORD_PC;
  assign fetch_logic_ctrls_2_down_Fetch_PC_FAULT = fetch_logic_ctrls_2_up_Fetch_PC_FAULT;
  assign fetch_logic_ctrls_2_down_Fetch_ID = fetch_logic_ctrls_2_up_Fetch_ID;
  assign fetch_logic_ctrls_2_down_Prediction_BRANCH_HISTORY = fetch_logic_ctrls_2_up_Prediction_BRANCH_HISTORY;
  assign fetch_logic_ctrls_2_down_FetchL1Plugin_logic_WAYS_TAGS_0_loaded = fetch_logic_ctrls_2_up_FetchL1Plugin_logic_WAYS_TAGS_0_loaded;
  assign fetch_logic_ctrls_2_down_FetchL1Plugin_logic_WAYS_TAGS_0_error = fetch_logic_ctrls_2_up_FetchL1Plugin_logic_WAYS_TAGS_0_error;
  assign fetch_logic_ctrls_2_down_FetchL1Plugin_logic_WAYS_TAGS_0_address = fetch_logic_ctrls_2_up_FetchL1Plugin_logic_WAYS_TAGS_0_address;
  assign fetch_logic_ctrls_2_down_FetchL1Plugin_logic_WAYS_TAGS_1_loaded = fetch_logic_ctrls_2_up_FetchL1Plugin_logic_WAYS_TAGS_1_loaded;
  assign fetch_logic_ctrls_2_down_FetchL1Plugin_logic_WAYS_TAGS_1_error = fetch_logic_ctrls_2_up_FetchL1Plugin_logic_WAYS_TAGS_1_error;
  assign fetch_logic_ctrls_2_down_FetchL1Plugin_logic_WAYS_TAGS_1_address = fetch_logic_ctrls_2_up_FetchL1Plugin_logic_WAYS_TAGS_1_address;
  assign fetch_logic_ctrls_2_down_FetchL1Plugin_logic_PLRU_BYPASSED_0 = fetch_logic_ctrls_2_up_FetchL1Plugin_logic_PLRU_BYPASSED_0;
  assign fetch_logic_ctrls_2_down_FetchL1Plugin_logic_BANKS_MUXES_0 = fetch_logic_ctrls_2_up_FetchL1Plugin_logic_BANKS_MUXES_0;
  assign fetch_logic_ctrls_2_down_FetchL1Plugin_logic_BANKS_MUXES_1 = fetch_logic_ctrls_2_up_FetchL1Plugin_logic_BANKS_MUXES_1;
  assign fetch_logic_ctrls_2_down_FetchL1Plugin_logic_HAZARD = fetch_logic_ctrls_2_up_FetchL1Plugin_logic_HAZARD;
  assign fetch_logic_ctrls_2_down_FetchL1Plugin_logic_WAYS_HITS_0 = fetch_logic_ctrls_2_up_FetchL1Plugin_logic_WAYS_HITS_0;
  assign fetch_logic_ctrls_2_down_FetchL1Plugin_logic_WAYS_HITS_1 = fetch_logic_ctrls_2_up_FetchL1Plugin_logic_WAYS_HITS_1;
  assign fetch_logic_ctrls_2_down_MMU_BYPASS_TRANSLATION = fetch_logic_ctrls_2_up_MMU_BYPASS_TRANSLATION;
  assign fetch_logic_ctrls_2_down_FetchL1Plugin_logic_WAYS_HIT = fetch_logic_ctrls_2_up_FetchL1Plugin_logic_WAYS_HIT;
  assign fetch_logic_ctrls_2_down_GSharePlugin_GSHARE_COUNTER_0 = fetch_logic_ctrls_2_up_GSharePlugin_GSHARE_COUNTER_0;
  assign fetch_logic_ctrls_2_down_GSharePlugin_GSHARE_COUNTER_1 = fetch_logic_ctrls_2_up_GSharePlugin_GSHARE_COUNTER_1;
  assign fetch_logic_ctrls_2_down_GSharePlugin_GSHARE_COUNTER_2 = fetch_logic_ctrls_2_up_GSharePlugin_GSHARE_COUNTER_2;
  assign fetch_logic_ctrls_2_down_GSharePlugin_GSHARE_COUNTER_3 = fetch_logic_ctrls_2_up_GSharePlugin_GSHARE_COUNTER_3;
  assign fetch_logic_ctrls_2_down_BtbPlugin_logic_chunksLogic_0_readRsp_ENTRY_hash = fetch_logic_ctrls_2_up_BtbPlugin_logic_chunksLogic_0_readRsp_ENTRY_hash;
  assign fetch_logic_ctrls_2_down_BtbPlugin_logic_chunksLogic_0_readRsp_ENTRY_sliceLow = fetch_logic_ctrls_2_up_BtbPlugin_logic_chunksLogic_0_readRsp_ENTRY_sliceLow;
  assign fetch_logic_ctrls_2_down_BtbPlugin_logic_chunksLogic_0_readRsp_ENTRY_pcTarget = fetch_logic_ctrls_2_up_BtbPlugin_logic_chunksLogic_0_readRsp_ENTRY_pcTarget;
  assign fetch_logic_ctrls_2_down_BtbPlugin_logic_chunksLogic_0_readRsp_ENTRY_isBranch = fetch_logic_ctrls_2_up_BtbPlugin_logic_chunksLogic_0_readRsp_ENTRY_isBranch;
  assign fetch_logic_ctrls_2_down_BtbPlugin_logic_chunksLogic_0_readRsp_ENTRY_isPush = fetch_logic_ctrls_2_up_BtbPlugin_logic_chunksLogic_0_readRsp_ENTRY_isPush;
  assign fetch_logic_ctrls_2_down_BtbPlugin_logic_chunksLogic_0_readRsp_ENTRY_isPop = fetch_logic_ctrls_2_up_BtbPlugin_logic_chunksLogic_0_readRsp_ENTRY_isPop;
  assign fetch_logic_ctrls_2_down_BtbPlugin_logic_chunksLogic_0_hitCalc_HIT = fetch_logic_ctrls_2_up_BtbPlugin_logic_chunksLogic_0_hitCalc_HIT;
  assign fetch_logic_ctrls_2_down_BtbPlugin_logic_chunksLogic_1_readRsp_ENTRY_hash = fetch_logic_ctrls_2_up_BtbPlugin_logic_chunksLogic_1_readRsp_ENTRY_hash;
  assign fetch_logic_ctrls_2_down_BtbPlugin_logic_chunksLogic_1_readRsp_ENTRY_sliceLow = fetch_logic_ctrls_2_up_BtbPlugin_logic_chunksLogic_1_readRsp_ENTRY_sliceLow;
  assign fetch_logic_ctrls_2_down_BtbPlugin_logic_chunksLogic_1_readRsp_ENTRY_pcTarget = fetch_logic_ctrls_2_up_BtbPlugin_logic_chunksLogic_1_readRsp_ENTRY_pcTarget;
  assign fetch_logic_ctrls_2_down_BtbPlugin_logic_chunksLogic_1_readRsp_ENTRY_isBranch = fetch_logic_ctrls_2_up_BtbPlugin_logic_chunksLogic_1_readRsp_ENTRY_isBranch;
  assign fetch_logic_ctrls_2_down_BtbPlugin_logic_chunksLogic_1_readRsp_ENTRY_isPush = fetch_logic_ctrls_2_up_BtbPlugin_logic_chunksLogic_1_readRsp_ENTRY_isPush;
  assign fetch_logic_ctrls_2_down_BtbPlugin_logic_chunksLogic_1_readRsp_ENTRY_isPop = fetch_logic_ctrls_2_up_BtbPlugin_logic_chunksLogic_1_readRsp_ENTRY_isPop;
  assign fetch_logic_ctrls_2_down_BtbPlugin_logic_chunksLogic_1_hitCalc_HIT = fetch_logic_ctrls_2_up_BtbPlugin_logic_chunksLogic_1_hitCalc_HIT;
  assign fetch_logic_ctrls_2_down_MMU_HAZARD = fetch_logic_ctrls_2_up_MMU_HAZARD;
  assign fetch_logic_ctrls_2_down_MMU_REFILL = fetch_logic_ctrls_2_up_MMU_REFILL;
  assign fetch_logic_ctrls_2_down_MMU_TRANSLATED = fetch_logic_ctrls_2_up_MMU_TRANSLATED;
  assign fetch_logic_ctrls_2_down_MMU_ALLOW_EXECUTE = fetch_logic_ctrls_2_up_MMU_ALLOW_EXECUTE;
  assign fetch_logic_ctrls_2_down_MMU_PAGE_FAULT = fetch_logic_ctrls_2_up_MMU_PAGE_FAULT;
  assign fetch_logic_ctrls_2_down_MMU_ACCESS_FAULT = fetch_logic_ctrls_2_up_MMU_ACCESS_FAULT;
  always @(*) begin
    toplevel_decode_ctrls_0_down_ready = toplevel_decode_ctrls_1_up_ready;
    if(when_StageLink_l67) begin
      toplevel_decode_ctrls_0_down_ready = 1'b1;
    end
  end

  assign when_StageLink_l67 = (! toplevel_decode_ctrls_1_up_isValid);
  assign when_DecodePipelinePlugin_l68 = ((! toplevel_decode_ctrls_1_up_isReady) && toplevel_decode_ctrls_1_lane0_upIsCancel);
  assign when_DecodePipelinePlugin_l68_1 = ((! toplevel_decode_ctrls_1_up_isReady) && toplevel_decode_ctrls_1_lane1_upIsCancel);
  assign toplevel_decode_ctrls_0_down_valid = toplevel_decode_ctrls_0_up_valid;
  assign toplevel_decode_ctrls_0_up_ready = toplevel_decode_ctrls_0_down_isReady;
  assign toplevel_decode_ctrls_0_down_Decode_INSTRUCTION_0 = toplevel_decode_ctrls_0_up_Decode_INSTRUCTION_0;
  assign toplevel_decode_ctrls_0_down_Decode_DECOMPRESSION_FAULT_0 = toplevel_decode_ctrls_0_up_Decode_DECOMPRESSION_FAULT_0;
  assign toplevel_decode_ctrls_0_down_Decode_INSTRUCTION_RAW_0 = toplevel_decode_ctrls_0_up_Decode_INSTRUCTION_RAW_0;
  assign toplevel_decode_ctrls_0_down_Decode_INSTRUCTION_SLICE_COUNT_0 = toplevel_decode_ctrls_0_up_Decode_INSTRUCTION_SLICE_COUNT_0;
  assign toplevel_decode_ctrls_0_down_PC_0 = toplevel_decode_ctrls_0_up_PC_0;
  assign toplevel_decode_ctrls_0_down_Decode_DOP_ID_0 = toplevel_decode_ctrls_0_up_Decode_DOP_ID_0;
  assign toplevel_decode_ctrls_0_down_Fetch_ID_0 = toplevel_decode_ctrls_0_up_Fetch_ID_0;
  assign toplevel_decode_ctrls_0_down_GSharePlugin_GSHARE_COUNTER_0_0 = toplevel_decode_ctrls_0_up_GSharePlugin_GSHARE_COUNTER_0_0;
  assign toplevel_decode_ctrls_0_down_GSharePlugin_GSHARE_COUNTER_0_1 = toplevel_decode_ctrls_0_up_GSharePlugin_GSHARE_COUNTER_0_1;
  assign toplevel_decode_ctrls_0_down_GSharePlugin_GSHARE_COUNTER_0_2 = toplevel_decode_ctrls_0_up_GSharePlugin_GSHARE_COUNTER_0_2;
  assign toplevel_decode_ctrls_0_down_GSharePlugin_GSHARE_COUNTER_0_3 = toplevel_decode_ctrls_0_up_GSharePlugin_GSHARE_COUNTER_0_3;
  assign toplevel_decode_ctrls_0_down_Prediction_BRANCH_HISTORY_0 = toplevel_decode_ctrls_0_up_Prediction_BRANCH_HISTORY_0;
  assign toplevel_decode_ctrls_0_down_TRAP_0 = toplevel_decode_ctrls_0_up_TRAP_0;
  assign toplevel_decode_ctrls_0_down_Prediction_ALIGNED_JUMPED_0 = toplevel_decode_ctrls_0_up_Prediction_ALIGNED_JUMPED_0;
  assign toplevel_decode_ctrls_0_down_Prediction_ALIGNED_JUMPED_PC_0 = toplevel_decode_ctrls_0_up_Prediction_ALIGNED_JUMPED_PC_0;
  assign toplevel_decode_ctrls_0_down_Prediction_ALIGNED_SLICES_BRANCH_0 = toplevel_decode_ctrls_0_up_Prediction_ALIGNED_SLICES_BRANCH_0;
  assign toplevel_decode_ctrls_0_down_Prediction_ALIGNED_SLICES_TAKEN_0 = toplevel_decode_ctrls_0_up_Prediction_ALIGNED_SLICES_TAKEN_0;
  assign toplevel_decode_ctrls_0_down_Prediction_ALIGN_REDO_0 = toplevel_decode_ctrls_0_up_Prediction_ALIGN_REDO_0;
  assign toplevel_decode_ctrls_0_down_Decode_INSTRUCTION_1 = toplevel_decode_ctrls_0_up_Decode_INSTRUCTION_1;
  assign toplevel_decode_ctrls_0_down_Decode_DECOMPRESSION_FAULT_1 = toplevel_decode_ctrls_0_up_Decode_DECOMPRESSION_FAULT_1;
  assign toplevel_decode_ctrls_0_down_Decode_INSTRUCTION_RAW_1 = toplevel_decode_ctrls_0_up_Decode_INSTRUCTION_RAW_1;
  assign toplevel_decode_ctrls_0_down_Decode_INSTRUCTION_SLICE_COUNT_1 = toplevel_decode_ctrls_0_up_Decode_INSTRUCTION_SLICE_COUNT_1;
  assign toplevel_decode_ctrls_0_down_PC_1 = toplevel_decode_ctrls_0_up_PC_1;
  assign toplevel_decode_ctrls_0_down_Decode_DOP_ID_1 = toplevel_decode_ctrls_0_up_Decode_DOP_ID_1;
  assign toplevel_decode_ctrls_0_down_Fetch_ID_1 = toplevel_decode_ctrls_0_up_Fetch_ID_1;
  assign toplevel_decode_ctrls_0_down_GSharePlugin_GSHARE_COUNTER_1_0 = toplevel_decode_ctrls_0_up_GSharePlugin_GSHARE_COUNTER_1_0;
  assign toplevel_decode_ctrls_0_down_GSharePlugin_GSHARE_COUNTER_1_1 = toplevel_decode_ctrls_0_up_GSharePlugin_GSHARE_COUNTER_1_1;
  assign toplevel_decode_ctrls_0_down_GSharePlugin_GSHARE_COUNTER_1_2 = toplevel_decode_ctrls_0_up_GSharePlugin_GSHARE_COUNTER_1_2;
  assign toplevel_decode_ctrls_0_down_GSharePlugin_GSHARE_COUNTER_1_3 = toplevel_decode_ctrls_0_up_GSharePlugin_GSHARE_COUNTER_1_3;
  assign toplevel_decode_ctrls_0_down_Prediction_BRANCH_HISTORY_1 = toplevel_decode_ctrls_0_up_Prediction_BRANCH_HISTORY_1;
  assign toplevel_decode_ctrls_0_down_TRAP_1 = toplevel_decode_ctrls_0_up_TRAP_1;
  assign toplevel_decode_ctrls_0_down_Prediction_ALIGNED_JUMPED_1 = toplevel_decode_ctrls_0_up_Prediction_ALIGNED_JUMPED_1;
  assign toplevel_decode_ctrls_0_down_Prediction_ALIGNED_JUMPED_PC_1 = toplevel_decode_ctrls_0_up_Prediction_ALIGNED_JUMPED_PC_1;
  assign toplevel_decode_ctrls_0_down_Prediction_ALIGNED_SLICES_BRANCH_1 = toplevel_decode_ctrls_0_up_Prediction_ALIGNED_SLICES_BRANCH_1;
  assign toplevel_decode_ctrls_0_down_Prediction_ALIGNED_SLICES_TAKEN_1 = toplevel_decode_ctrls_0_up_Prediction_ALIGNED_SLICES_TAKEN_1;
  assign toplevel_decode_ctrls_0_down_Prediction_ALIGN_REDO_1 = toplevel_decode_ctrls_0_up_Prediction_ALIGN_REDO_1;
  assign toplevel_decode_ctrls_1_down_valid = toplevel_decode_ctrls_1_up_valid;
  assign toplevel_decode_ctrls_1_up_ready = toplevel_decode_ctrls_1_down_isReady;
  assign toplevel_decode_ctrls_1_down_Decode_INSTRUCTION_0 = toplevel_decode_ctrls_1_up_Decode_INSTRUCTION_0;
  assign toplevel_decode_ctrls_1_down_Decode_DECOMPRESSION_FAULT_0 = toplevel_decode_ctrls_1_up_Decode_DECOMPRESSION_FAULT_0;
  assign toplevel_decode_ctrls_1_down_Decode_INSTRUCTION_RAW_0 = toplevel_decode_ctrls_1_up_Decode_INSTRUCTION_RAW_0;
  assign toplevel_decode_ctrls_1_down_Decode_INSTRUCTION_SLICE_COUNT_0 = toplevel_decode_ctrls_1_up_Decode_INSTRUCTION_SLICE_COUNT_0;
  assign toplevel_decode_ctrls_1_down_PC_0 = toplevel_decode_ctrls_1_up_PC_0;
  assign toplevel_decode_ctrls_1_down_Decode_DOP_ID_0 = toplevel_decode_ctrls_1_up_Decode_DOP_ID_0;
  assign toplevel_decode_ctrls_1_down_GSharePlugin_GSHARE_COUNTER_0_0 = toplevel_decode_ctrls_1_up_GSharePlugin_GSHARE_COUNTER_0_0;
  assign toplevel_decode_ctrls_1_down_GSharePlugin_GSHARE_COUNTER_0_1 = toplevel_decode_ctrls_1_up_GSharePlugin_GSHARE_COUNTER_0_1;
  assign toplevel_decode_ctrls_1_down_GSharePlugin_GSHARE_COUNTER_0_2 = toplevel_decode_ctrls_1_up_GSharePlugin_GSHARE_COUNTER_0_2;
  assign toplevel_decode_ctrls_1_down_GSharePlugin_GSHARE_COUNTER_0_3 = toplevel_decode_ctrls_1_up_GSharePlugin_GSHARE_COUNTER_0_3;
  assign toplevel_decode_ctrls_1_down_Prediction_BRANCH_HISTORY_0 = toplevel_decode_ctrls_1_up_Prediction_BRANCH_HISTORY_0;
  assign toplevel_decode_ctrls_1_down_Prediction_ALIGNED_JUMPED_0 = toplevel_decode_ctrls_1_up_Prediction_ALIGNED_JUMPED_0;
  assign toplevel_decode_ctrls_1_down_Prediction_ALIGNED_JUMPED_PC_0 = toplevel_decode_ctrls_1_up_Prediction_ALIGNED_JUMPED_PC_0;
  assign toplevel_decode_ctrls_1_down_Prediction_ALIGNED_SLICES_BRANCH_0 = toplevel_decode_ctrls_1_up_Prediction_ALIGNED_SLICES_BRANCH_0;
  assign toplevel_decode_ctrls_1_down_Prediction_ALIGNED_SLICES_TAKEN_0 = toplevel_decode_ctrls_1_up_Prediction_ALIGNED_SLICES_TAKEN_0;
  assign toplevel_decode_ctrls_1_down_Prediction_ALIGN_REDO_0 = toplevel_decode_ctrls_1_up_Prediction_ALIGN_REDO_0;
  assign toplevel_decode_ctrls_1_down_Decode_INSTRUCTION_1 = toplevel_decode_ctrls_1_up_Decode_INSTRUCTION_1;
  assign toplevel_decode_ctrls_1_down_Decode_DECOMPRESSION_FAULT_1 = toplevel_decode_ctrls_1_up_Decode_DECOMPRESSION_FAULT_1;
  assign toplevel_decode_ctrls_1_down_Decode_INSTRUCTION_RAW_1 = toplevel_decode_ctrls_1_up_Decode_INSTRUCTION_RAW_1;
  assign toplevel_decode_ctrls_1_down_Decode_INSTRUCTION_SLICE_COUNT_1 = toplevel_decode_ctrls_1_up_Decode_INSTRUCTION_SLICE_COUNT_1;
  assign toplevel_decode_ctrls_1_down_PC_1 = toplevel_decode_ctrls_1_up_PC_1;
  assign toplevel_decode_ctrls_1_down_Decode_DOP_ID_1 = toplevel_decode_ctrls_1_up_Decode_DOP_ID_1;
  assign toplevel_decode_ctrls_1_down_GSharePlugin_GSHARE_COUNTER_1_0 = toplevel_decode_ctrls_1_up_GSharePlugin_GSHARE_COUNTER_1_0;
  assign toplevel_decode_ctrls_1_down_GSharePlugin_GSHARE_COUNTER_1_1 = toplevel_decode_ctrls_1_up_GSharePlugin_GSHARE_COUNTER_1_1;
  assign toplevel_decode_ctrls_1_down_GSharePlugin_GSHARE_COUNTER_1_2 = toplevel_decode_ctrls_1_up_GSharePlugin_GSHARE_COUNTER_1_2;
  assign toplevel_decode_ctrls_1_down_GSharePlugin_GSHARE_COUNTER_1_3 = toplevel_decode_ctrls_1_up_GSharePlugin_GSHARE_COUNTER_1_3;
  assign toplevel_decode_ctrls_1_down_Prediction_BRANCH_HISTORY_1 = toplevel_decode_ctrls_1_up_Prediction_BRANCH_HISTORY_1;
  assign toplevel_decode_ctrls_1_down_Prediction_ALIGNED_JUMPED_1 = toplevel_decode_ctrls_1_up_Prediction_ALIGNED_JUMPED_1;
  assign toplevel_decode_ctrls_1_down_Prediction_ALIGNED_JUMPED_PC_1 = toplevel_decode_ctrls_1_up_Prediction_ALIGNED_JUMPED_PC_1;
  assign toplevel_decode_ctrls_1_down_Prediction_ALIGNED_SLICES_BRANCH_1 = toplevel_decode_ctrls_1_up_Prediction_ALIGNED_SLICES_BRANCH_1;
  assign toplevel_decode_ctrls_1_down_Prediction_ALIGNED_SLICES_TAKEN_1 = toplevel_decode_ctrls_1_up_Prediction_ALIGNED_SLICES_TAKEN_1;
  assign toplevel_decode_ctrls_1_down_Prediction_ALIGN_REDO_1 = toplevel_decode_ctrls_1_up_Prediction_ALIGN_REDO_1;
  assign toplevel_execute_ctrl0_down_ready = toplevel_execute_ctrl1_up_ready;
  assign toplevel_execute_ctrl1_down_ready = toplevel_execute_ctrl2_up_ready;
  assign toplevel_execute_ctrl2_down_ready = toplevel_execute_ctrl3_up_ready;
  assign toplevel_execute_ctrl3_down_ready = toplevel_execute_ctrl4_up_ready;
  assign toplevel_execute_ctrl4_down_ready = toplevel_execute_ctrl5_up_ready;
  assign toplevel_execute_ctrl0_up_ready = toplevel_execute_ctrl0_down_isReady;
  assign toplevel_execute_ctrl0_down_Decode_UOP_lane0 = toplevel_execute_ctrl0_up_Decode_UOP_lane0;
  assign toplevel_execute_ctrl0_down_Prediction_ALIGNED_JUMPED_lane0 = toplevel_execute_ctrl0_up_Prediction_ALIGNED_JUMPED_lane0;
  assign toplevel_execute_ctrl0_down_Prediction_ALIGNED_JUMPED_PC_lane0 = toplevel_execute_ctrl0_up_Prediction_ALIGNED_JUMPED_PC_lane0;
  assign toplevel_execute_ctrl0_down_Prediction_ALIGNED_SLICES_TAKEN_lane0 = toplevel_execute_ctrl0_up_Prediction_ALIGNED_SLICES_TAKEN_lane0;
  assign toplevel_execute_ctrl0_down_Prediction_ALIGNED_SLICES_BRANCH_lane0 = toplevel_execute_ctrl0_up_Prediction_ALIGNED_SLICES_BRANCH_lane0;
  assign toplevel_execute_ctrl0_down_GSharePlugin_GSHARE_COUNTER_lane0_0 = toplevel_execute_ctrl0_up_GSharePlugin_GSHARE_COUNTER_lane0_0;
  assign toplevel_execute_ctrl0_down_GSharePlugin_GSHARE_COUNTER_lane0_1 = toplevel_execute_ctrl0_up_GSharePlugin_GSHARE_COUNTER_lane0_1;
  assign toplevel_execute_ctrl0_down_GSharePlugin_GSHARE_COUNTER_lane0_2 = toplevel_execute_ctrl0_up_GSharePlugin_GSHARE_COUNTER_lane0_2;
  assign toplevel_execute_ctrl0_down_GSharePlugin_GSHARE_COUNTER_lane0_3 = toplevel_execute_ctrl0_up_GSharePlugin_GSHARE_COUNTER_lane0_3;
  assign toplevel_execute_ctrl0_down_Prediction_BRANCH_HISTORY_lane0 = toplevel_execute_ctrl0_up_Prediction_BRANCH_HISTORY_lane0;
  assign toplevel_execute_ctrl0_down_Decode_INSTRUCTION_SLICE_COUNT_lane0 = toplevel_execute_ctrl0_up_Decode_INSTRUCTION_SLICE_COUNT_lane0;
  assign toplevel_execute_ctrl0_down_PC_lane0 = toplevel_execute_ctrl0_up_PC_lane0;
  assign toplevel_execute_ctrl0_down_TRAP_lane0 = toplevel_execute_ctrl0_up_TRAP_lane0;
  assign toplevel_execute_ctrl0_down_Decode_UOP_ID_lane0 = toplevel_execute_ctrl0_up_Decode_UOP_ID_lane0;
  assign toplevel_execute_ctrl0_down_RS1_PHYS_lane0 = toplevel_execute_ctrl0_up_RS1_PHYS_lane0;
  assign toplevel_execute_ctrl0_down_RS2_PHYS_lane0 = toplevel_execute_ctrl0_up_RS2_PHYS_lane0;
  assign toplevel_execute_ctrl0_down_RD_PHYS_lane0 = toplevel_execute_ctrl0_up_RD_PHYS_lane0;
  assign toplevel_execute_ctrl0_down_LANE_AGE_lane0 = toplevel_execute_ctrl0_up_LANE_AGE_lane0;
  assign toplevel_execute_ctrl0_down_COMPLETED_lane0 = toplevel_execute_ctrl0_up_COMPLETED_lane0;
  assign toplevel_execute_ctrl0_down_execute_lane0_LAYER_SEL_lane0 = toplevel_execute_ctrl0_up_execute_lane0_LAYER_SEL_lane0;
  assign toplevel_execute_ctrl0_down_Decode_UOP_lane1 = toplevel_execute_ctrl0_up_Decode_UOP_lane1;
  assign toplevel_execute_ctrl0_down_Prediction_ALIGNED_JUMPED_lane1 = toplevel_execute_ctrl0_up_Prediction_ALIGNED_JUMPED_lane1;
  assign toplevel_execute_ctrl0_down_Prediction_ALIGNED_JUMPED_PC_lane1 = toplevel_execute_ctrl0_up_Prediction_ALIGNED_JUMPED_PC_lane1;
  assign toplevel_execute_ctrl0_down_Prediction_ALIGNED_SLICES_TAKEN_lane1 = toplevel_execute_ctrl0_up_Prediction_ALIGNED_SLICES_TAKEN_lane1;
  assign toplevel_execute_ctrl0_down_Prediction_ALIGNED_SLICES_BRANCH_lane1 = toplevel_execute_ctrl0_up_Prediction_ALIGNED_SLICES_BRANCH_lane1;
  assign toplevel_execute_ctrl0_down_GSharePlugin_GSHARE_COUNTER_lane1_0 = toplevel_execute_ctrl0_up_GSharePlugin_GSHARE_COUNTER_lane1_0;
  assign toplevel_execute_ctrl0_down_GSharePlugin_GSHARE_COUNTER_lane1_1 = toplevel_execute_ctrl0_up_GSharePlugin_GSHARE_COUNTER_lane1_1;
  assign toplevel_execute_ctrl0_down_GSharePlugin_GSHARE_COUNTER_lane1_2 = toplevel_execute_ctrl0_up_GSharePlugin_GSHARE_COUNTER_lane1_2;
  assign toplevel_execute_ctrl0_down_GSharePlugin_GSHARE_COUNTER_lane1_3 = toplevel_execute_ctrl0_up_GSharePlugin_GSHARE_COUNTER_lane1_3;
  assign toplevel_execute_ctrl0_down_Prediction_BRANCH_HISTORY_lane1 = toplevel_execute_ctrl0_up_Prediction_BRANCH_HISTORY_lane1;
  assign toplevel_execute_ctrl0_down_Decode_INSTRUCTION_SLICE_COUNT_lane1 = toplevel_execute_ctrl0_up_Decode_INSTRUCTION_SLICE_COUNT_lane1;
  assign toplevel_execute_ctrl0_down_PC_lane1 = toplevel_execute_ctrl0_up_PC_lane1;
  assign toplevel_execute_ctrl0_down_TRAP_lane1 = toplevel_execute_ctrl0_up_TRAP_lane1;
  assign toplevel_execute_ctrl0_down_Decode_UOP_ID_lane1 = toplevel_execute_ctrl0_up_Decode_UOP_ID_lane1;
  assign toplevel_execute_ctrl0_down_RS1_PHYS_lane1 = toplevel_execute_ctrl0_up_RS1_PHYS_lane1;
  assign toplevel_execute_ctrl0_down_RS2_PHYS_lane1 = toplevel_execute_ctrl0_up_RS2_PHYS_lane1;
  assign toplevel_execute_ctrl0_down_RD_PHYS_lane1 = toplevel_execute_ctrl0_up_RD_PHYS_lane1;
  assign toplevel_execute_ctrl0_down_LANE_AGE_lane1 = toplevel_execute_ctrl0_up_LANE_AGE_lane1;
  assign toplevel_execute_ctrl0_down_COMPLETED_lane1 = toplevel_execute_ctrl0_up_COMPLETED_lane1;
  assign toplevel_execute_ctrl0_down_execute_lane1_LAYER_SEL_lane1 = toplevel_execute_ctrl0_up_execute_lane1_LAYER_SEL_lane1;
  assign toplevel_execute_ctrl1_up_ready = toplevel_execute_ctrl1_down_isReady;
  assign toplevel_execute_ctrl1_down_Decode_UOP_lane0 = toplevel_execute_ctrl1_up_Decode_UOP_lane0;
  assign toplevel_execute_ctrl1_down_Prediction_ALIGNED_JUMPED_lane0 = toplevel_execute_ctrl1_up_Prediction_ALIGNED_JUMPED_lane0;
  assign toplevel_execute_ctrl1_down_Prediction_ALIGNED_JUMPED_PC_lane0 = toplevel_execute_ctrl1_up_Prediction_ALIGNED_JUMPED_PC_lane0;
  assign toplevel_execute_ctrl1_down_Prediction_ALIGNED_SLICES_TAKEN_lane0 = toplevel_execute_ctrl1_up_Prediction_ALIGNED_SLICES_TAKEN_lane0;
  assign toplevel_execute_ctrl1_down_Prediction_ALIGNED_SLICES_BRANCH_lane0 = toplevel_execute_ctrl1_up_Prediction_ALIGNED_SLICES_BRANCH_lane0;
  assign toplevel_execute_ctrl1_down_GSharePlugin_GSHARE_COUNTER_lane0_0 = toplevel_execute_ctrl1_up_GSharePlugin_GSHARE_COUNTER_lane0_0;
  assign toplevel_execute_ctrl1_down_GSharePlugin_GSHARE_COUNTER_lane0_1 = toplevel_execute_ctrl1_up_GSharePlugin_GSHARE_COUNTER_lane0_1;
  assign toplevel_execute_ctrl1_down_GSharePlugin_GSHARE_COUNTER_lane0_2 = toplevel_execute_ctrl1_up_GSharePlugin_GSHARE_COUNTER_lane0_2;
  assign toplevel_execute_ctrl1_down_GSharePlugin_GSHARE_COUNTER_lane0_3 = toplevel_execute_ctrl1_up_GSharePlugin_GSHARE_COUNTER_lane0_3;
  assign toplevel_execute_ctrl1_down_Prediction_BRANCH_HISTORY_lane0 = toplevel_execute_ctrl1_up_Prediction_BRANCH_HISTORY_lane0;
  assign toplevel_execute_ctrl1_down_Decode_INSTRUCTION_SLICE_COUNT_lane0 = toplevel_execute_ctrl1_up_Decode_INSTRUCTION_SLICE_COUNT_lane0;
  assign toplevel_execute_ctrl1_down_PC_lane0 = toplevel_execute_ctrl1_up_PC_lane0;
  assign toplevel_execute_ctrl1_down_TRAP_lane0 = toplevel_execute_ctrl1_up_TRAP_lane0;
  assign toplevel_execute_ctrl1_down_Decode_UOP_ID_lane0 = toplevel_execute_ctrl1_up_Decode_UOP_ID_lane0;
  assign toplevel_execute_ctrl1_down_RS1_PHYS_lane0 = toplevel_execute_ctrl1_up_RS1_PHYS_lane0;
  assign toplevel_execute_ctrl1_down_RS2_PHYS_lane0 = toplevel_execute_ctrl1_up_RS2_PHYS_lane0;
  assign toplevel_execute_ctrl1_down_RD_PHYS_lane0 = toplevel_execute_ctrl1_up_RD_PHYS_lane0;
  assign toplevel_execute_ctrl1_down_LANE_AGE_lane0 = toplevel_execute_ctrl1_up_LANE_AGE_lane0;
  assign toplevel_execute_ctrl1_down_COMPLETED_lane0 = toplevel_execute_ctrl1_up_COMPLETED_lane0;
  assign toplevel_execute_ctrl1_down_execute_lane0_LAYER_SEL_lane0 = toplevel_execute_ctrl1_up_execute_lane0_LAYER_SEL_lane0;
  assign toplevel_execute_ctrl1_down_Decode_UOP_lane1 = toplevel_execute_ctrl1_up_Decode_UOP_lane1;
  assign toplevel_execute_ctrl1_down_Prediction_ALIGNED_JUMPED_lane1 = toplevel_execute_ctrl1_up_Prediction_ALIGNED_JUMPED_lane1;
  assign toplevel_execute_ctrl1_down_Prediction_ALIGNED_JUMPED_PC_lane1 = toplevel_execute_ctrl1_up_Prediction_ALIGNED_JUMPED_PC_lane1;
  assign toplevel_execute_ctrl1_down_Prediction_ALIGNED_SLICES_TAKEN_lane1 = toplevel_execute_ctrl1_up_Prediction_ALIGNED_SLICES_TAKEN_lane1;
  assign toplevel_execute_ctrl1_down_Prediction_ALIGNED_SLICES_BRANCH_lane1 = toplevel_execute_ctrl1_up_Prediction_ALIGNED_SLICES_BRANCH_lane1;
  assign toplevel_execute_ctrl1_down_GSharePlugin_GSHARE_COUNTER_lane1_0 = toplevel_execute_ctrl1_up_GSharePlugin_GSHARE_COUNTER_lane1_0;
  assign toplevel_execute_ctrl1_down_GSharePlugin_GSHARE_COUNTER_lane1_1 = toplevel_execute_ctrl1_up_GSharePlugin_GSHARE_COUNTER_lane1_1;
  assign toplevel_execute_ctrl1_down_GSharePlugin_GSHARE_COUNTER_lane1_2 = toplevel_execute_ctrl1_up_GSharePlugin_GSHARE_COUNTER_lane1_2;
  assign toplevel_execute_ctrl1_down_GSharePlugin_GSHARE_COUNTER_lane1_3 = toplevel_execute_ctrl1_up_GSharePlugin_GSHARE_COUNTER_lane1_3;
  assign toplevel_execute_ctrl1_down_Prediction_BRANCH_HISTORY_lane1 = toplevel_execute_ctrl1_up_Prediction_BRANCH_HISTORY_lane1;
  assign toplevel_execute_ctrl1_down_Decode_INSTRUCTION_SLICE_COUNT_lane1 = toplevel_execute_ctrl1_up_Decode_INSTRUCTION_SLICE_COUNT_lane1;
  assign toplevel_execute_ctrl1_down_PC_lane1 = toplevel_execute_ctrl1_up_PC_lane1;
  assign toplevel_execute_ctrl1_down_TRAP_lane1 = toplevel_execute_ctrl1_up_TRAP_lane1;
  assign toplevel_execute_ctrl1_down_Decode_UOP_ID_lane1 = toplevel_execute_ctrl1_up_Decode_UOP_ID_lane1;
  assign toplevel_execute_ctrl1_down_RS1_PHYS_lane1 = toplevel_execute_ctrl1_up_RS1_PHYS_lane1;
  assign toplevel_execute_ctrl1_down_RS2_PHYS_lane1 = toplevel_execute_ctrl1_up_RS2_PHYS_lane1;
  assign toplevel_execute_ctrl1_down_RD_PHYS_lane1 = toplevel_execute_ctrl1_up_RD_PHYS_lane1;
  assign toplevel_execute_ctrl1_down_LANE_AGE_lane1 = toplevel_execute_ctrl1_up_LANE_AGE_lane1;
  assign toplevel_execute_ctrl1_down_COMPLETED_lane1 = toplevel_execute_ctrl1_up_COMPLETED_lane1;
  assign toplevel_execute_ctrl1_down_execute_lane1_LAYER_SEL_lane1 = toplevel_execute_ctrl1_up_execute_lane1_LAYER_SEL_lane1;
  assign toplevel_execute_ctrl1_down_AguPlugin_SIZE_lane0 = toplevel_execute_ctrl1_up_AguPlugin_SIZE_lane0;
  assign toplevel_execute_ctrl2_up_ready = toplevel_execute_ctrl2_down_isReady;
  assign toplevel_execute_ctrl2_down_Decode_UOP_lane0 = toplevel_execute_ctrl2_up_Decode_UOP_lane0;
  assign toplevel_execute_ctrl2_down_Prediction_ALIGNED_JUMPED_lane0 = toplevel_execute_ctrl2_up_Prediction_ALIGNED_JUMPED_lane0;
  assign toplevel_execute_ctrl2_down_Prediction_ALIGNED_JUMPED_PC_lane0 = toplevel_execute_ctrl2_up_Prediction_ALIGNED_JUMPED_PC_lane0;
  assign toplevel_execute_ctrl2_down_Prediction_ALIGNED_SLICES_TAKEN_lane0 = toplevel_execute_ctrl2_up_Prediction_ALIGNED_SLICES_TAKEN_lane0;
  assign toplevel_execute_ctrl2_down_Prediction_ALIGNED_SLICES_BRANCH_lane0 = toplevel_execute_ctrl2_up_Prediction_ALIGNED_SLICES_BRANCH_lane0;
  assign toplevel_execute_ctrl2_down_GSharePlugin_GSHARE_COUNTER_lane0_0 = toplevel_execute_ctrl2_up_GSharePlugin_GSHARE_COUNTER_lane0_0;
  assign toplevel_execute_ctrl2_down_GSharePlugin_GSHARE_COUNTER_lane0_1 = toplevel_execute_ctrl2_up_GSharePlugin_GSHARE_COUNTER_lane0_1;
  assign toplevel_execute_ctrl2_down_GSharePlugin_GSHARE_COUNTER_lane0_2 = toplevel_execute_ctrl2_up_GSharePlugin_GSHARE_COUNTER_lane0_2;
  assign toplevel_execute_ctrl2_down_GSharePlugin_GSHARE_COUNTER_lane0_3 = toplevel_execute_ctrl2_up_GSharePlugin_GSHARE_COUNTER_lane0_3;
  assign toplevel_execute_ctrl2_down_Prediction_BRANCH_HISTORY_lane0 = toplevel_execute_ctrl2_up_Prediction_BRANCH_HISTORY_lane0;
  assign toplevel_execute_ctrl2_down_Decode_INSTRUCTION_SLICE_COUNT_lane0 = toplevel_execute_ctrl2_up_Decode_INSTRUCTION_SLICE_COUNT_lane0;
  assign toplevel_execute_ctrl2_down_PC_lane0 = toplevel_execute_ctrl2_up_PC_lane0;
  assign toplevel_execute_ctrl2_down_Decode_UOP_ID_lane0 = toplevel_execute_ctrl2_up_Decode_UOP_ID_lane0;
  assign toplevel_execute_ctrl2_down_RS1_PHYS_lane0 = toplevel_execute_ctrl2_up_RS1_PHYS_lane0;
  assign toplevel_execute_ctrl2_down_RS2_PHYS_lane0 = toplevel_execute_ctrl2_up_RS2_PHYS_lane0;
  assign toplevel_execute_ctrl2_down_RD_PHYS_lane0 = toplevel_execute_ctrl2_up_RD_PHYS_lane0;
  assign toplevel_execute_ctrl2_down_LANE_AGE_lane0 = toplevel_execute_ctrl2_up_LANE_AGE_lane0;
  assign toplevel_execute_ctrl2_down_Decode_UOP_lane1 = toplevel_execute_ctrl2_up_Decode_UOP_lane1;
  assign toplevel_execute_ctrl2_down_Prediction_ALIGNED_JUMPED_lane1 = toplevel_execute_ctrl2_up_Prediction_ALIGNED_JUMPED_lane1;
  assign toplevel_execute_ctrl2_down_Prediction_ALIGNED_JUMPED_PC_lane1 = toplevel_execute_ctrl2_up_Prediction_ALIGNED_JUMPED_PC_lane1;
  assign toplevel_execute_ctrl2_down_Prediction_ALIGNED_SLICES_TAKEN_lane1 = toplevel_execute_ctrl2_up_Prediction_ALIGNED_SLICES_TAKEN_lane1;
  assign toplevel_execute_ctrl2_down_Prediction_ALIGNED_SLICES_BRANCH_lane1 = toplevel_execute_ctrl2_up_Prediction_ALIGNED_SLICES_BRANCH_lane1;
  assign toplevel_execute_ctrl2_down_GSharePlugin_GSHARE_COUNTER_lane1_0 = toplevel_execute_ctrl2_up_GSharePlugin_GSHARE_COUNTER_lane1_0;
  assign toplevel_execute_ctrl2_down_GSharePlugin_GSHARE_COUNTER_lane1_1 = toplevel_execute_ctrl2_up_GSharePlugin_GSHARE_COUNTER_lane1_1;
  assign toplevel_execute_ctrl2_down_GSharePlugin_GSHARE_COUNTER_lane1_2 = toplevel_execute_ctrl2_up_GSharePlugin_GSHARE_COUNTER_lane1_2;
  assign toplevel_execute_ctrl2_down_GSharePlugin_GSHARE_COUNTER_lane1_3 = toplevel_execute_ctrl2_up_GSharePlugin_GSHARE_COUNTER_lane1_3;
  assign toplevel_execute_ctrl2_down_Prediction_BRANCH_HISTORY_lane1 = toplevel_execute_ctrl2_up_Prediction_BRANCH_HISTORY_lane1;
  assign toplevel_execute_ctrl2_down_Decode_INSTRUCTION_SLICE_COUNT_lane1 = toplevel_execute_ctrl2_up_Decode_INSTRUCTION_SLICE_COUNT_lane1;
  assign toplevel_execute_ctrl2_down_PC_lane1 = toplevel_execute_ctrl2_up_PC_lane1;
  assign toplevel_execute_ctrl2_down_TRAP_lane1 = toplevel_execute_ctrl2_up_TRAP_lane1;
  assign toplevel_execute_ctrl2_down_Decode_UOP_ID_lane1 = toplevel_execute_ctrl2_up_Decode_UOP_ID_lane1;
  assign toplevel_execute_ctrl2_down_RS1_PHYS_lane1 = toplevel_execute_ctrl2_up_RS1_PHYS_lane1;
  assign toplevel_execute_ctrl2_down_RS2_PHYS_lane1 = toplevel_execute_ctrl2_up_RS2_PHYS_lane1;
  assign toplevel_execute_ctrl2_down_RD_PHYS_lane1 = toplevel_execute_ctrl2_up_RD_PHYS_lane1;
  assign toplevel_execute_ctrl2_down_LANE_AGE_lane1 = toplevel_execute_ctrl2_up_LANE_AGE_lane1;
  assign toplevel_execute_ctrl2_down_AguPlugin_SIZE_lane0 = toplevel_execute_ctrl2_up_AguPlugin_SIZE_lane0;
  assign toplevel_execute_ctrl2_down_early0_SrcPlugin_SRC1_lane0 = toplevel_execute_ctrl2_up_early0_SrcPlugin_SRC1_lane0;
  assign toplevel_execute_ctrl2_down_early0_SrcPlugin_SRC2_lane0 = toplevel_execute_ctrl2_up_early0_SrcPlugin_SRC2_lane0;
  assign toplevel_execute_ctrl2_down_early1_SrcPlugin_SRC1_lane1 = toplevel_execute_ctrl2_up_early1_SrcPlugin_SRC1_lane1;
  assign toplevel_execute_ctrl2_down_early1_SrcPlugin_SRC2_lane1 = toplevel_execute_ctrl2_up_early1_SrcPlugin_SRC2_lane1;
  assign toplevel_execute_ctrl2_down_MAY_FLUSH_PRECISE_3_lane0 = toplevel_execute_ctrl2_up_MAY_FLUSH_PRECISE_3_lane0;
  assign toplevel_execute_ctrl2_down_MAY_FLUSH_PRECISE_3_lane1 = toplevel_execute_ctrl2_up_MAY_FLUSH_PRECISE_3_lane1;
  assign toplevel_execute_ctrl2_down_early0_IntAluPlugin_SEL_lane0 = toplevel_execute_ctrl2_up_early0_IntAluPlugin_SEL_lane0;
  assign toplevel_execute_ctrl2_down_early0_BarrelShifterPlugin_SEL_lane0 = toplevel_execute_ctrl2_up_early0_BarrelShifterPlugin_SEL_lane0;
  assign toplevel_execute_ctrl2_down_early0_BranchPlugin_SEL_lane0 = toplevel_execute_ctrl2_up_early0_BranchPlugin_SEL_lane0;
  assign toplevel_execute_ctrl2_down_early0_MulPlugin_SEL_lane0 = toplevel_execute_ctrl2_up_early0_MulPlugin_SEL_lane0;
  assign toplevel_execute_ctrl2_down_early0_DivPlugin_SEL_lane0 = toplevel_execute_ctrl2_up_early0_DivPlugin_SEL_lane0;
  assign toplevel_execute_ctrl2_down_early0_EnvPlugin_SEL_lane0 = toplevel_execute_ctrl2_up_early0_EnvPlugin_SEL_lane0;
  assign toplevel_execute_ctrl2_down_late0_IntAluPlugin_SEL_lane0 = toplevel_execute_ctrl2_up_late0_IntAluPlugin_SEL_lane0;
  assign toplevel_execute_ctrl2_down_late0_BarrelShifterPlugin_SEL_lane0 = toplevel_execute_ctrl2_up_late0_BarrelShifterPlugin_SEL_lane0;
  assign toplevel_execute_ctrl2_down_late0_BranchPlugin_SEL_lane0 = toplevel_execute_ctrl2_up_late0_BranchPlugin_SEL_lane0;
  assign toplevel_execute_ctrl2_down_MulPlugin_HIGH_lane0 = toplevel_execute_ctrl2_up_MulPlugin_HIGH_lane0;
  assign toplevel_execute_ctrl2_down_CsrAccessPlugin_SEL_lane0 = toplevel_execute_ctrl2_up_CsrAccessPlugin_SEL_lane0;
  assign toplevel_execute_ctrl2_down_AguPlugin_SEL_lane0 = toplevel_execute_ctrl2_up_AguPlugin_SEL_lane0;
  assign toplevel_execute_ctrl2_down_LsuPlugin_logic_FENCE_lane0 = toplevel_execute_ctrl2_up_LsuPlugin_logic_FENCE_lane0;
  assign toplevel_execute_ctrl2_down_lane0_integer_WriteBackPlugin_SEL_lane0 = toplevel_execute_ctrl2_up_lane0_integer_WriteBackPlugin_SEL_lane0;
  assign toplevel_execute_ctrl2_down_COMPLETION_AT_2_lane0 = toplevel_execute_ctrl2_up_COMPLETION_AT_2_lane0;
  assign toplevel_execute_ctrl2_down_COMPLETION_AT_3_lane0 = toplevel_execute_ctrl2_up_COMPLETION_AT_3_lane0;
  assign toplevel_execute_ctrl2_down_COMPLETION_AT_4_lane0 = toplevel_execute_ctrl2_up_COMPLETION_AT_4_lane0;
  assign toplevel_execute_ctrl2_down_execute_lane0_logic_completions_onCtrl_0_ENABLE_lane0 = toplevel_execute_ctrl2_up_execute_lane0_logic_completions_onCtrl_0_ENABLE_lane0;
  assign toplevel_execute_ctrl2_down_execute_lane0_logic_completions_onCtrl_1_ENABLE_lane0 = toplevel_execute_ctrl2_up_execute_lane0_logic_completions_onCtrl_1_ENABLE_lane0;
  assign toplevel_execute_ctrl2_down_execute_lane0_logic_completions_onCtrl_2_ENABLE_lane0 = toplevel_execute_ctrl2_up_execute_lane0_logic_completions_onCtrl_2_ENABLE_lane0;
  assign toplevel_execute_ctrl2_down_early0_IntAluPlugin_ALU_ADD_SUB_lane0 = toplevel_execute_ctrl2_up_early0_IntAluPlugin_ALU_ADD_SUB_lane0;
  assign toplevel_execute_ctrl2_down_early0_IntAluPlugin_ALU_SLTX_lane0 = toplevel_execute_ctrl2_up_early0_IntAluPlugin_ALU_SLTX_lane0;
  assign toplevel_execute_ctrl2_down_early0_IntAluPlugin_ALU_BITWISE_CTRL_lane0 = toplevel_execute_ctrl2_up_early0_IntAluPlugin_ALU_BITWISE_CTRL_lane0;
  assign toplevel_execute_ctrl2_down_SrcStageables_REVERT_lane0 = toplevel_execute_ctrl2_up_SrcStageables_REVERT_lane0;
  assign toplevel_execute_ctrl2_down_SrcStageables_ZERO_lane0 = toplevel_execute_ctrl2_up_SrcStageables_ZERO_lane0;
  assign toplevel_execute_ctrl2_down_lane0_IntFormatPlugin_logic_SIGNED_lane0 = toplevel_execute_ctrl2_up_lane0_IntFormatPlugin_logic_SIGNED_lane0;
  assign toplevel_execute_ctrl2_down_lane0_IntFormatPlugin_logic_WIDTH_ID_lane0 = toplevel_execute_ctrl2_up_lane0_IntFormatPlugin_logic_WIDTH_ID_lane0;
  assign toplevel_execute_ctrl2_down_BYPASSED_AT_3_lane0 = toplevel_execute_ctrl2_up_BYPASSED_AT_3_lane0;
  assign toplevel_execute_ctrl2_down_SrcStageables_UNSIGNED_lane0 = toplevel_execute_ctrl2_up_SrcStageables_UNSIGNED_lane0;
  assign toplevel_execute_ctrl2_down_BarrelShifterPlugin_LEFT_lane0 = toplevel_execute_ctrl2_up_BarrelShifterPlugin_LEFT_lane0;
  assign toplevel_execute_ctrl2_down_BarrelShifterPlugin_SIGNED_lane0 = toplevel_execute_ctrl2_up_BarrelShifterPlugin_SIGNED_lane0;
  assign toplevel_execute_ctrl2_down_BranchPlugin_BRANCH_CTRL_lane0 = toplevel_execute_ctrl2_up_BranchPlugin_BRANCH_CTRL_lane0;
  assign toplevel_execute_ctrl2_down_RsUnsignedPlugin_RS1_SIGNED_lane0 = toplevel_execute_ctrl2_up_RsUnsignedPlugin_RS1_SIGNED_lane0;
  assign toplevel_execute_ctrl2_down_RsUnsignedPlugin_RS2_SIGNED_lane0 = toplevel_execute_ctrl2_up_RsUnsignedPlugin_RS2_SIGNED_lane0;
  assign toplevel_execute_ctrl2_down_DivPlugin_REM_lane0 = toplevel_execute_ctrl2_up_DivPlugin_REM_lane0;
  assign toplevel_execute_ctrl2_down_CsrAccessPlugin_CSR_IMM_lane0 = toplevel_execute_ctrl2_up_CsrAccessPlugin_CSR_IMM_lane0;
  assign toplevel_execute_ctrl2_down_CsrAccessPlugin_CSR_MASK_lane0 = toplevel_execute_ctrl2_up_CsrAccessPlugin_CSR_MASK_lane0;
  assign toplevel_execute_ctrl2_down_CsrAccessPlugin_CSR_CLEAR_lane0 = toplevel_execute_ctrl2_up_CsrAccessPlugin_CSR_CLEAR_lane0;
  assign toplevel_execute_ctrl2_down_AguPlugin_LOAD_lane0 = toplevel_execute_ctrl2_up_AguPlugin_LOAD_lane0;
  assign toplevel_execute_ctrl2_down_AguPlugin_STORE_lane0 = toplevel_execute_ctrl2_up_AguPlugin_STORE_lane0;
  assign toplevel_execute_ctrl2_down_AguPlugin_ATOMIC_lane0 = toplevel_execute_ctrl2_up_AguPlugin_ATOMIC_lane0;
  assign toplevel_execute_ctrl2_down_AguPlugin_FLOAT_lane0 = toplevel_execute_ctrl2_up_AguPlugin_FLOAT_lane0;
  assign toplevel_execute_ctrl2_down_LsuPlugin_logic_LSU_PREFETCH_lane0 = toplevel_execute_ctrl2_up_LsuPlugin_logic_LSU_PREFETCH_lane0;
  assign toplevel_execute_ctrl2_down_early0_EnvPlugin_OP_lane0 = toplevel_execute_ctrl2_up_early0_EnvPlugin_OP_lane0;
  assign toplevel_execute_ctrl2_down_late0_IntAluPlugin_ALU_ADD_SUB_lane0 = toplevel_execute_ctrl2_up_late0_IntAluPlugin_ALU_ADD_SUB_lane0;
  assign toplevel_execute_ctrl2_down_late0_IntAluPlugin_ALU_SLTX_lane0 = toplevel_execute_ctrl2_up_late0_IntAluPlugin_ALU_SLTX_lane0;
  assign toplevel_execute_ctrl2_down_late0_IntAluPlugin_ALU_BITWISE_CTRL_lane0 = toplevel_execute_ctrl2_up_late0_IntAluPlugin_ALU_BITWISE_CTRL_lane0;
  assign toplevel_execute_ctrl2_down_late0_SrcPlugin_logic_SRC1_CTRL_lane0 = toplevel_execute_ctrl2_up_late0_SrcPlugin_logic_SRC1_CTRL_lane0;
  assign toplevel_execute_ctrl2_down_late0_SrcPlugin_logic_SRC2_CTRL_lane0 = toplevel_execute_ctrl2_up_late0_SrcPlugin_logic_SRC2_CTRL_lane0;
  assign toplevel_execute_ctrl2_down_early1_IntAluPlugin_SEL_lane1 = toplevel_execute_ctrl2_up_early1_IntAluPlugin_SEL_lane1;
  assign toplevel_execute_ctrl2_down_early1_BarrelShifterPlugin_SEL_lane1 = toplevel_execute_ctrl2_up_early1_BarrelShifterPlugin_SEL_lane1;
  assign toplevel_execute_ctrl2_down_early1_BranchPlugin_SEL_lane1 = toplevel_execute_ctrl2_up_early1_BranchPlugin_SEL_lane1;
  assign toplevel_execute_ctrl2_down_late1_IntAluPlugin_SEL_lane1 = toplevel_execute_ctrl2_up_late1_IntAluPlugin_SEL_lane1;
  assign toplevel_execute_ctrl2_down_late1_BarrelShifterPlugin_SEL_lane1 = toplevel_execute_ctrl2_up_late1_BarrelShifterPlugin_SEL_lane1;
  assign toplevel_execute_ctrl2_down_late1_BranchPlugin_SEL_lane1 = toplevel_execute_ctrl2_up_late1_BranchPlugin_SEL_lane1;
  assign toplevel_execute_ctrl2_down_lane1_integer_WriteBackPlugin_SEL_lane1 = toplevel_execute_ctrl2_up_lane1_integer_WriteBackPlugin_SEL_lane1;
  assign toplevel_execute_ctrl2_down_COMPLETION_AT_2_lane1 = toplevel_execute_ctrl2_up_COMPLETION_AT_2_lane1;
  assign toplevel_execute_ctrl2_down_COMPLETION_AT_3_lane1 = toplevel_execute_ctrl2_up_COMPLETION_AT_3_lane1;
  assign toplevel_execute_ctrl2_down_COMPLETION_AT_4_lane1 = toplevel_execute_ctrl2_up_COMPLETION_AT_4_lane1;
  assign toplevel_execute_ctrl2_down_execute_lane1_logic_completions_onCtrl_0_ENABLE_lane1 = toplevel_execute_ctrl2_up_execute_lane1_logic_completions_onCtrl_0_ENABLE_lane1;
  assign toplevel_execute_ctrl2_down_execute_lane1_logic_completions_onCtrl_1_ENABLE_lane1 = toplevel_execute_ctrl2_up_execute_lane1_logic_completions_onCtrl_1_ENABLE_lane1;
  assign toplevel_execute_ctrl2_down_execute_lane1_logic_completions_onCtrl_2_ENABLE_lane1 = toplevel_execute_ctrl2_up_execute_lane1_logic_completions_onCtrl_2_ENABLE_lane1;
  assign toplevel_execute_ctrl2_down_early1_IntAluPlugin_ALU_ADD_SUB_lane1 = toplevel_execute_ctrl2_up_early1_IntAluPlugin_ALU_ADD_SUB_lane1;
  assign toplevel_execute_ctrl2_down_early1_IntAluPlugin_ALU_SLTX_lane1 = toplevel_execute_ctrl2_up_early1_IntAluPlugin_ALU_SLTX_lane1;
  assign toplevel_execute_ctrl2_down_early1_IntAluPlugin_ALU_BITWISE_CTRL_lane1 = toplevel_execute_ctrl2_up_early1_IntAluPlugin_ALU_BITWISE_CTRL_lane1;
  assign toplevel_execute_ctrl2_down_SrcStageables_REVERT_lane1 = toplevel_execute_ctrl2_up_SrcStageables_REVERT_lane1;
  assign toplevel_execute_ctrl2_down_SrcStageables_ZERO_lane1 = toplevel_execute_ctrl2_up_SrcStageables_ZERO_lane1;
  assign toplevel_execute_ctrl2_down_BYPASSED_AT_3_lane1 = toplevel_execute_ctrl2_up_BYPASSED_AT_3_lane1;
  assign toplevel_execute_ctrl2_down_SrcStageables_UNSIGNED_lane1 = toplevel_execute_ctrl2_up_SrcStageables_UNSIGNED_lane1;
  assign toplevel_execute_ctrl2_down_BarrelShifterPlugin_LEFT_lane1 = toplevel_execute_ctrl2_up_BarrelShifterPlugin_LEFT_lane1;
  assign toplevel_execute_ctrl2_down_BarrelShifterPlugin_SIGNED_lane1 = toplevel_execute_ctrl2_up_BarrelShifterPlugin_SIGNED_lane1;
  assign toplevel_execute_ctrl2_down_BranchPlugin_BRANCH_CTRL_lane1 = toplevel_execute_ctrl2_up_BranchPlugin_BRANCH_CTRL_lane1;
  assign toplevel_execute_ctrl2_down_late1_IntAluPlugin_ALU_ADD_SUB_lane1 = toplevel_execute_ctrl2_up_late1_IntAluPlugin_ALU_ADD_SUB_lane1;
  assign toplevel_execute_ctrl2_down_late1_IntAluPlugin_ALU_SLTX_lane1 = toplevel_execute_ctrl2_up_late1_IntAluPlugin_ALU_SLTX_lane1;
  assign toplevel_execute_ctrl2_down_late1_IntAluPlugin_ALU_BITWISE_CTRL_lane1 = toplevel_execute_ctrl2_up_late1_IntAluPlugin_ALU_BITWISE_CTRL_lane1;
  assign toplevel_execute_ctrl2_down_late1_SrcPlugin_logic_SRC1_CTRL_lane1 = toplevel_execute_ctrl2_up_late1_SrcPlugin_logic_SRC1_CTRL_lane1;
  assign toplevel_execute_ctrl2_down_late1_SrcPlugin_logic_SRC2_CTRL_lane1 = toplevel_execute_ctrl2_up_late1_SrcPlugin_logic_SRC2_CTRL_lane1;
  assign toplevel_execute_ctrl2_down_COMMIT_lane1 = toplevel_execute_ctrl2_up_COMMIT_lane1;
  assign toplevel_execute_ctrl3_up_ready = toplevel_execute_ctrl3_down_isReady;
  assign toplevel_execute_ctrl3_down_Decode_UOP_lane0 = toplevel_execute_ctrl3_up_Decode_UOP_lane0;
  assign toplevel_execute_ctrl3_down_Prediction_ALIGNED_JUMPED_lane0 = toplevel_execute_ctrl3_up_Prediction_ALIGNED_JUMPED_lane0;
  assign toplevel_execute_ctrl3_down_Prediction_ALIGNED_JUMPED_PC_lane0 = toplevel_execute_ctrl3_up_Prediction_ALIGNED_JUMPED_PC_lane0;
  assign toplevel_execute_ctrl3_down_Prediction_ALIGNED_SLICES_TAKEN_lane0 = toplevel_execute_ctrl3_up_Prediction_ALIGNED_SLICES_TAKEN_lane0;
  assign toplevel_execute_ctrl3_down_Prediction_ALIGNED_SLICES_BRANCH_lane0 = toplevel_execute_ctrl3_up_Prediction_ALIGNED_SLICES_BRANCH_lane0;
  assign toplevel_execute_ctrl3_down_GSharePlugin_GSHARE_COUNTER_lane0_0 = toplevel_execute_ctrl3_up_GSharePlugin_GSHARE_COUNTER_lane0_0;
  assign toplevel_execute_ctrl3_down_GSharePlugin_GSHARE_COUNTER_lane0_1 = toplevel_execute_ctrl3_up_GSharePlugin_GSHARE_COUNTER_lane0_1;
  assign toplevel_execute_ctrl3_down_GSharePlugin_GSHARE_COUNTER_lane0_2 = toplevel_execute_ctrl3_up_GSharePlugin_GSHARE_COUNTER_lane0_2;
  assign toplevel_execute_ctrl3_down_GSharePlugin_GSHARE_COUNTER_lane0_3 = toplevel_execute_ctrl3_up_GSharePlugin_GSHARE_COUNTER_lane0_3;
  assign toplevel_execute_ctrl3_down_Prediction_BRANCH_HISTORY_lane0 = toplevel_execute_ctrl3_up_Prediction_BRANCH_HISTORY_lane0;
  assign toplevel_execute_ctrl3_down_Decode_INSTRUCTION_SLICE_COUNT_lane0 = toplevel_execute_ctrl3_up_Decode_INSTRUCTION_SLICE_COUNT_lane0;
  assign toplevel_execute_ctrl3_down_PC_lane0 = toplevel_execute_ctrl3_up_PC_lane0;
  assign toplevel_execute_ctrl3_down_TRAP_lane0 = toplevel_execute_ctrl3_up_TRAP_lane0;
  assign toplevel_execute_ctrl3_down_Decode_UOP_ID_lane0 = toplevel_execute_ctrl3_up_Decode_UOP_ID_lane0;
  assign toplevel_execute_ctrl3_down_RS1_PHYS_lane0 = toplevel_execute_ctrl3_up_RS1_PHYS_lane0;
  assign toplevel_execute_ctrl3_down_RS2_PHYS_lane0 = toplevel_execute_ctrl3_up_RS2_PHYS_lane0;
  assign toplevel_execute_ctrl3_down_RD_PHYS_lane0 = toplevel_execute_ctrl3_up_RD_PHYS_lane0;
  assign toplevel_execute_ctrl3_down_LANE_AGE_lane0 = toplevel_execute_ctrl3_up_LANE_AGE_lane0;
  assign toplevel_execute_ctrl3_down_Decode_UOP_lane1 = toplevel_execute_ctrl3_up_Decode_UOP_lane1;
  assign toplevel_execute_ctrl3_down_Prediction_ALIGNED_JUMPED_lane1 = toplevel_execute_ctrl3_up_Prediction_ALIGNED_JUMPED_lane1;
  assign toplevel_execute_ctrl3_down_Prediction_ALIGNED_JUMPED_PC_lane1 = toplevel_execute_ctrl3_up_Prediction_ALIGNED_JUMPED_PC_lane1;
  assign toplevel_execute_ctrl3_down_Prediction_ALIGNED_SLICES_TAKEN_lane1 = toplevel_execute_ctrl3_up_Prediction_ALIGNED_SLICES_TAKEN_lane1;
  assign toplevel_execute_ctrl3_down_Prediction_ALIGNED_SLICES_BRANCH_lane1 = toplevel_execute_ctrl3_up_Prediction_ALIGNED_SLICES_BRANCH_lane1;
  assign toplevel_execute_ctrl3_down_GSharePlugin_GSHARE_COUNTER_lane1_0 = toplevel_execute_ctrl3_up_GSharePlugin_GSHARE_COUNTER_lane1_0;
  assign toplevel_execute_ctrl3_down_GSharePlugin_GSHARE_COUNTER_lane1_1 = toplevel_execute_ctrl3_up_GSharePlugin_GSHARE_COUNTER_lane1_1;
  assign toplevel_execute_ctrl3_down_GSharePlugin_GSHARE_COUNTER_lane1_2 = toplevel_execute_ctrl3_up_GSharePlugin_GSHARE_COUNTER_lane1_2;
  assign toplevel_execute_ctrl3_down_GSharePlugin_GSHARE_COUNTER_lane1_3 = toplevel_execute_ctrl3_up_GSharePlugin_GSHARE_COUNTER_lane1_3;
  assign toplevel_execute_ctrl3_down_Prediction_BRANCH_HISTORY_lane1 = toplevel_execute_ctrl3_up_Prediction_BRANCH_HISTORY_lane1;
  assign toplevel_execute_ctrl3_down_Decode_INSTRUCTION_SLICE_COUNT_lane1 = toplevel_execute_ctrl3_up_Decode_INSTRUCTION_SLICE_COUNT_lane1;
  assign toplevel_execute_ctrl3_down_PC_lane1 = toplevel_execute_ctrl3_up_PC_lane1;
  assign toplevel_execute_ctrl3_down_TRAP_lane1 = toplevel_execute_ctrl3_up_TRAP_lane1;
  assign toplevel_execute_ctrl3_down_Decode_UOP_ID_lane1 = toplevel_execute_ctrl3_up_Decode_UOP_ID_lane1;
  assign toplevel_execute_ctrl3_down_RS1_PHYS_lane1 = toplevel_execute_ctrl3_up_RS1_PHYS_lane1;
  assign toplevel_execute_ctrl3_down_RS2_PHYS_lane1 = toplevel_execute_ctrl3_up_RS2_PHYS_lane1;
  assign toplevel_execute_ctrl3_down_RD_PHYS_lane1 = toplevel_execute_ctrl3_up_RD_PHYS_lane1;
  assign toplevel_execute_ctrl3_down_LANE_AGE_lane1 = toplevel_execute_ctrl3_up_LANE_AGE_lane1;
  assign toplevel_execute_ctrl3_down_AguPlugin_SIZE_lane0 = toplevel_execute_ctrl3_up_AguPlugin_SIZE_lane0;
  assign toplevel_execute_ctrl3_down_early0_BarrelShifterPlugin_SEL_lane0 = toplevel_execute_ctrl3_up_early0_BarrelShifterPlugin_SEL_lane0;
  assign toplevel_execute_ctrl3_down_early0_BranchPlugin_SEL_lane0 = toplevel_execute_ctrl3_up_early0_BranchPlugin_SEL_lane0;
  assign toplevel_execute_ctrl3_down_early0_MulPlugin_SEL_lane0 = toplevel_execute_ctrl3_up_early0_MulPlugin_SEL_lane0;
  assign toplevel_execute_ctrl3_down_early0_DivPlugin_SEL_lane0 = toplevel_execute_ctrl3_up_early0_DivPlugin_SEL_lane0;
  assign toplevel_execute_ctrl3_down_late0_IntAluPlugin_SEL_lane0 = toplevel_execute_ctrl3_up_late0_IntAluPlugin_SEL_lane0;
  assign toplevel_execute_ctrl3_down_late0_BarrelShifterPlugin_SEL_lane0 = toplevel_execute_ctrl3_up_late0_BarrelShifterPlugin_SEL_lane0;
  assign toplevel_execute_ctrl3_down_late0_BranchPlugin_SEL_lane0 = toplevel_execute_ctrl3_up_late0_BranchPlugin_SEL_lane0;
  assign toplevel_execute_ctrl3_down_MulPlugin_HIGH_lane0 = toplevel_execute_ctrl3_up_MulPlugin_HIGH_lane0;
  assign toplevel_execute_ctrl3_down_CsrAccessPlugin_SEL_lane0 = toplevel_execute_ctrl3_up_CsrAccessPlugin_SEL_lane0;
  assign toplevel_execute_ctrl3_down_AguPlugin_SEL_lane0 = toplevel_execute_ctrl3_up_AguPlugin_SEL_lane0;
  assign toplevel_execute_ctrl3_down_LsuPlugin_logic_FENCE_lane0 = toplevel_execute_ctrl3_up_LsuPlugin_logic_FENCE_lane0;
  assign toplevel_execute_ctrl3_down_lane0_integer_WriteBackPlugin_SEL_lane0 = toplevel_execute_ctrl3_up_lane0_integer_WriteBackPlugin_SEL_lane0;
  assign toplevel_execute_ctrl3_down_COMPLETION_AT_3_lane0 = toplevel_execute_ctrl3_up_COMPLETION_AT_3_lane0;
  assign toplevel_execute_ctrl3_down_COMPLETION_AT_4_lane0 = toplevel_execute_ctrl3_up_COMPLETION_AT_4_lane0;
  assign toplevel_execute_ctrl3_down_execute_lane0_logic_completions_onCtrl_1_ENABLE_lane0 = toplevel_execute_ctrl3_up_execute_lane0_logic_completions_onCtrl_1_ENABLE_lane0;
  assign toplevel_execute_ctrl3_down_execute_lane0_logic_completions_onCtrl_2_ENABLE_lane0 = toplevel_execute_ctrl3_up_execute_lane0_logic_completions_onCtrl_2_ENABLE_lane0;
  assign toplevel_execute_ctrl3_down_SrcStageables_REVERT_lane0 = toplevel_execute_ctrl3_up_SrcStageables_REVERT_lane0;
  assign toplevel_execute_ctrl3_down_SrcStageables_ZERO_lane0 = toplevel_execute_ctrl3_up_SrcStageables_ZERO_lane0;
  assign toplevel_execute_ctrl3_down_lane0_IntFormatPlugin_logic_SIGNED_lane0 = toplevel_execute_ctrl3_up_lane0_IntFormatPlugin_logic_SIGNED_lane0;
  assign toplevel_execute_ctrl3_down_lane0_IntFormatPlugin_logic_WIDTH_ID_lane0 = toplevel_execute_ctrl3_up_lane0_IntFormatPlugin_logic_WIDTH_ID_lane0;
  assign toplevel_execute_ctrl3_down_SrcStageables_UNSIGNED_lane0 = toplevel_execute_ctrl3_up_SrcStageables_UNSIGNED_lane0;
  assign toplevel_execute_ctrl3_down_BarrelShifterPlugin_LEFT_lane0 = toplevel_execute_ctrl3_up_BarrelShifterPlugin_LEFT_lane0;
  assign toplevel_execute_ctrl3_down_BarrelShifterPlugin_SIGNED_lane0 = toplevel_execute_ctrl3_up_BarrelShifterPlugin_SIGNED_lane0;
  assign toplevel_execute_ctrl3_down_BranchPlugin_BRANCH_CTRL_lane0 = toplevel_execute_ctrl3_up_BranchPlugin_BRANCH_CTRL_lane0;
  assign toplevel_execute_ctrl3_down_AguPlugin_LOAD_lane0 = toplevel_execute_ctrl3_up_AguPlugin_LOAD_lane0;
  assign toplevel_execute_ctrl3_down_AguPlugin_STORE_lane0 = toplevel_execute_ctrl3_up_AguPlugin_STORE_lane0;
  assign toplevel_execute_ctrl3_down_AguPlugin_ATOMIC_lane0 = toplevel_execute_ctrl3_up_AguPlugin_ATOMIC_lane0;
  assign toplevel_execute_ctrl3_down_AguPlugin_FLOAT_lane0 = toplevel_execute_ctrl3_up_AguPlugin_FLOAT_lane0;
  assign toplevel_execute_ctrl3_down_LsuPlugin_logic_LSU_PREFETCH_lane0 = toplevel_execute_ctrl3_up_LsuPlugin_logic_LSU_PREFETCH_lane0;
  assign toplevel_execute_ctrl3_down_late0_IntAluPlugin_ALU_ADD_SUB_lane0 = toplevel_execute_ctrl3_up_late0_IntAluPlugin_ALU_ADD_SUB_lane0;
  assign toplevel_execute_ctrl3_down_late0_IntAluPlugin_ALU_SLTX_lane0 = toplevel_execute_ctrl3_up_late0_IntAluPlugin_ALU_SLTX_lane0;
  assign toplevel_execute_ctrl3_down_late0_IntAluPlugin_ALU_BITWISE_CTRL_lane0 = toplevel_execute_ctrl3_up_late0_IntAluPlugin_ALU_BITWISE_CTRL_lane0;
  assign toplevel_execute_ctrl3_down_late0_SrcPlugin_logic_SRC1_CTRL_lane0 = toplevel_execute_ctrl3_up_late0_SrcPlugin_logic_SRC1_CTRL_lane0;
  assign toplevel_execute_ctrl3_down_late0_SrcPlugin_logic_SRC2_CTRL_lane0 = toplevel_execute_ctrl3_up_late0_SrcPlugin_logic_SRC2_CTRL_lane0;
  assign toplevel_execute_ctrl3_down_early1_BarrelShifterPlugin_SEL_lane1 = toplevel_execute_ctrl3_up_early1_BarrelShifterPlugin_SEL_lane1;
  assign toplevel_execute_ctrl3_down_early1_BranchPlugin_SEL_lane1 = toplevel_execute_ctrl3_up_early1_BranchPlugin_SEL_lane1;
  assign toplevel_execute_ctrl3_down_late1_IntAluPlugin_SEL_lane1 = toplevel_execute_ctrl3_up_late1_IntAluPlugin_SEL_lane1;
  assign toplevel_execute_ctrl3_down_late1_BarrelShifterPlugin_SEL_lane1 = toplevel_execute_ctrl3_up_late1_BarrelShifterPlugin_SEL_lane1;
  assign toplevel_execute_ctrl3_down_late1_BranchPlugin_SEL_lane1 = toplevel_execute_ctrl3_up_late1_BranchPlugin_SEL_lane1;
  assign toplevel_execute_ctrl3_down_lane1_integer_WriteBackPlugin_SEL_lane1 = toplevel_execute_ctrl3_up_lane1_integer_WriteBackPlugin_SEL_lane1;
  assign toplevel_execute_ctrl3_down_COMPLETION_AT_3_lane1 = toplevel_execute_ctrl3_up_COMPLETION_AT_3_lane1;
  assign toplevel_execute_ctrl3_down_COMPLETION_AT_4_lane1 = toplevel_execute_ctrl3_up_COMPLETION_AT_4_lane1;
  assign toplevel_execute_ctrl3_down_execute_lane1_logic_completions_onCtrl_1_ENABLE_lane1 = toplevel_execute_ctrl3_up_execute_lane1_logic_completions_onCtrl_1_ENABLE_lane1;
  assign toplevel_execute_ctrl3_down_execute_lane1_logic_completions_onCtrl_2_ENABLE_lane1 = toplevel_execute_ctrl3_up_execute_lane1_logic_completions_onCtrl_2_ENABLE_lane1;
  assign toplevel_execute_ctrl3_down_SrcStageables_REVERT_lane1 = toplevel_execute_ctrl3_up_SrcStageables_REVERT_lane1;
  assign toplevel_execute_ctrl3_down_SrcStageables_ZERO_lane1 = toplevel_execute_ctrl3_up_SrcStageables_ZERO_lane1;
  assign toplevel_execute_ctrl3_down_SrcStageables_UNSIGNED_lane1 = toplevel_execute_ctrl3_up_SrcStageables_UNSIGNED_lane1;
  assign toplevel_execute_ctrl3_down_BarrelShifterPlugin_LEFT_lane1 = toplevel_execute_ctrl3_up_BarrelShifterPlugin_LEFT_lane1;
  assign toplevel_execute_ctrl3_down_BarrelShifterPlugin_SIGNED_lane1 = toplevel_execute_ctrl3_up_BarrelShifterPlugin_SIGNED_lane1;
  assign toplevel_execute_ctrl3_down_BranchPlugin_BRANCH_CTRL_lane1 = toplevel_execute_ctrl3_up_BranchPlugin_BRANCH_CTRL_lane1;
  assign toplevel_execute_ctrl3_down_late1_IntAluPlugin_ALU_ADD_SUB_lane1 = toplevel_execute_ctrl3_up_late1_IntAluPlugin_ALU_ADD_SUB_lane1;
  assign toplevel_execute_ctrl3_down_late1_IntAluPlugin_ALU_SLTX_lane1 = toplevel_execute_ctrl3_up_late1_IntAluPlugin_ALU_SLTX_lane1;
  assign toplevel_execute_ctrl3_down_late1_IntAluPlugin_ALU_BITWISE_CTRL_lane1 = toplevel_execute_ctrl3_up_late1_IntAluPlugin_ALU_BITWISE_CTRL_lane1;
  assign toplevel_execute_ctrl3_down_late1_SrcPlugin_logic_SRC1_CTRL_lane1 = toplevel_execute_ctrl3_up_late1_SrcPlugin_logic_SRC1_CTRL_lane1;
  assign toplevel_execute_ctrl3_down_late1_SrcPlugin_logic_SRC2_CTRL_lane1 = toplevel_execute_ctrl3_up_late1_SrcPlugin_logic_SRC2_CTRL_lane1;
  assign toplevel_execute_ctrl3_down_COMMIT_lane0 = toplevel_execute_ctrl3_up_COMMIT_lane0;
  assign toplevel_execute_ctrl3_down_COMMIT_lane1 = toplevel_execute_ctrl3_up_COMMIT_lane1;
  assign toplevel_execute_ctrl3_down_early0_SrcPlugin_ADD_SUB_lane0 = toplevel_execute_ctrl3_up_early0_SrcPlugin_ADD_SUB_lane0;
  assign toplevel_execute_ctrl3_down_early0_SrcPlugin_LESS_lane0 = toplevel_execute_ctrl3_up_early0_SrcPlugin_LESS_lane0;
  assign toplevel_execute_ctrl3_down_early0_BarrelShifterPlugin_SHIFT_RESULT_lane0 = toplevel_execute_ctrl3_up_early0_BarrelShifterPlugin_SHIFT_RESULT_lane0;
  assign toplevel_execute_ctrl3_down_MUL_SRC1_lane0 = toplevel_execute_ctrl3_up_MUL_SRC1_lane0;
  assign toplevel_execute_ctrl3_down_MUL_SRC2_lane0 = toplevel_execute_ctrl3_up_MUL_SRC2_lane0;
  assign toplevel_execute_ctrl3_down_DivPlugin_DIV_RESULT_lane0 = toplevel_execute_ctrl3_up_DivPlugin_DIV_RESULT_lane0;
  assign toplevel_execute_ctrl3_down_early1_SrcPlugin_LESS_lane1 = toplevel_execute_ctrl3_up_early1_SrcPlugin_LESS_lane1;
  assign toplevel_execute_ctrl3_down_early1_BarrelShifterPlugin_SHIFT_RESULT_lane1 = toplevel_execute_ctrl3_up_early1_BarrelShifterPlugin_SHIFT_RESULT_lane1;
  assign toplevel_execute_ctrl3_down_early0_BranchPlugin_pcCalc_PC_TRUE_lane0 = toplevel_execute_ctrl3_up_early0_BranchPlugin_pcCalc_PC_TRUE_lane0;
  assign toplevel_execute_ctrl3_down_early0_BranchPlugin_pcCalc_PC_FALSE_lane0 = toplevel_execute_ctrl3_up_early0_BranchPlugin_pcCalc_PC_FALSE_lane0;
  assign toplevel_execute_ctrl3_down_early0_BranchPlugin_pcCalc_PC_LAST_SLICE_lane0 = toplevel_execute_ctrl3_up_early0_BranchPlugin_pcCalc_PC_LAST_SLICE_lane0;
  assign toplevel_execute_ctrl3_down_early1_BranchPlugin_pcCalc_PC_TRUE_lane1 = toplevel_execute_ctrl3_up_early1_BranchPlugin_pcCalc_PC_TRUE_lane1;
  assign toplevel_execute_ctrl3_down_early1_BranchPlugin_pcCalc_PC_FALSE_lane1 = toplevel_execute_ctrl3_up_early1_BranchPlugin_pcCalc_PC_FALSE_lane1;
  assign toplevel_execute_ctrl3_down_early1_BranchPlugin_pcCalc_PC_LAST_SLICE_lane1 = toplevel_execute_ctrl3_up_early1_BranchPlugin_pcCalc_PC_LAST_SLICE_lane1;
  assign toplevel_execute_ctrl3_down_early0_BranchPlugin_logic_alu_EQ_lane0 = toplevel_execute_ctrl3_up_early0_BranchPlugin_logic_alu_EQ_lane0;
  assign toplevel_execute_ctrl3_down_early0_BranchPlugin_logic_alu_btb_BAD_TARGET_lane0 = toplevel_execute_ctrl3_up_early0_BranchPlugin_logic_alu_btb_BAD_TARGET_lane0;
  assign toplevel_execute_ctrl3_down_early0_BranchPlugin_logic_alu_MSB_FAILED_lane0 = toplevel_execute_ctrl3_up_early0_BranchPlugin_logic_alu_MSB_FAILED_lane0;
  assign toplevel_execute_ctrl3_down_early1_BranchPlugin_logic_alu_EQ_lane1 = toplevel_execute_ctrl3_up_early1_BranchPlugin_logic_alu_EQ_lane1;
  assign toplevel_execute_ctrl3_down_early1_BranchPlugin_logic_alu_btb_BAD_TARGET_lane1 = toplevel_execute_ctrl3_up_early1_BranchPlugin_logic_alu_btb_BAD_TARGET_lane1;
  assign toplevel_execute_ctrl3_down_early1_BranchPlugin_logic_alu_MSB_FAILED_lane1 = toplevel_execute_ctrl3_up_early1_BranchPlugin_logic_alu_MSB_FAILED_lane1;
  assign toplevel_execute_ctrl3_down_LsuL1_MIXED_ADDRESS_lane0 = toplevel_execute_ctrl3_up_LsuL1_MIXED_ADDRESS_lane0;
  assign toplevel_execute_ctrl3_down_LsuL1Plugin_logic_BANK_BUSY_lane0 = toplevel_execute_ctrl3_up_LsuL1Plugin_logic_BANK_BUSY_lane0;
  assign toplevel_execute_ctrl3_down_LsuL1Plugin_logic_EVENT_WRITE_VALID_lane0 = toplevel_execute_ctrl3_up_LsuL1Plugin_logic_EVENT_WRITE_VALID_lane0;
  assign toplevel_execute_ctrl3_down_LsuL1Plugin_logic_EVENT_WRITE_ADDRESS_lane0 = toplevel_execute_ctrl3_up_LsuL1Plugin_logic_EVENT_WRITE_ADDRESS_lane0;
  assign toplevel_execute_ctrl3_down_LsuL1Plugin_logic_ls_rt0_SHARED_BYPASS_VALID_lane0 = toplevel_execute_ctrl3_up_LsuL1Plugin_logic_ls_rt0_SHARED_BYPASS_VALID_lane0;
  assign toplevel_execute_ctrl3_down_LsuL1Plugin_logic_ls_rt0_SHARED_BYPASS_VALUE_lane0_plru_0 = toplevel_execute_ctrl3_up_LsuL1Plugin_logic_ls_rt0_SHARED_BYPASS_VALUE_lane0_plru_0;
  assign toplevel_execute_ctrl3_down_LsuL1Plugin_logic_ls_rt0_SHARED_BYPASS_VALUE_lane0_dirty = toplevel_execute_ctrl3_up_LsuL1Plugin_logic_ls_rt0_SHARED_BYPASS_VALUE_lane0_dirty;
  assign toplevel_execute_ctrl3_down_LsuL1Plugin_logic_EVENT_WRITE_DATA_lane0 = toplevel_execute_ctrl3_up_LsuL1Plugin_logic_EVENT_WRITE_DATA_lane0;
  assign toplevel_execute_ctrl3_down_LsuL1Plugin_logic_EVENT_WRITE_MASK_lane0 = toplevel_execute_ctrl3_up_LsuL1Plugin_logic_EVENT_WRITE_MASK_lane0;
  assign toplevel_execute_ctrl3_down_LsuPlugin_logic_FORCE_PHYSICAL_lane0 = toplevel_execute_ctrl3_up_LsuPlugin_logic_FORCE_PHYSICAL_lane0;
  assign toplevel_execute_ctrl3_down_LsuPlugin_logic_FROM_ACCESS_lane0 = toplevel_execute_ctrl3_up_LsuPlugin_logic_FROM_ACCESS_lane0;
  assign toplevel_execute_ctrl3_down_LsuL1_MASK_lane0 = toplevel_execute_ctrl3_up_LsuL1_MASK_lane0;
  assign toplevel_execute_ctrl3_down_LsuL1_SIZE_lane0 = toplevel_execute_ctrl3_up_LsuL1_SIZE_lane0;
  assign toplevel_execute_ctrl3_down_LsuL1_LOAD_lane0 = toplevel_execute_ctrl3_up_LsuL1_LOAD_lane0;
  assign toplevel_execute_ctrl3_down_LsuL1_ATOMIC_lane0 = toplevel_execute_ctrl3_up_LsuL1_ATOMIC_lane0;
  assign toplevel_execute_ctrl3_down_LsuL1_STORE_lane0 = toplevel_execute_ctrl3_up_LsuL1_STORE_lane0;
  assign toplevel_execute_ctrl3_down_LsuL1_PREFETCH_lane0 = toplevel_execute_ctrl3_up_LsuL1_PREFETCH_lane0;
  assign toplevel_execute_ctrl3_down_LsuL1_FLUSH_lane0 = toplevel_execute_ctrl3_up_LsuL1_FLUSH_lane0;
  assign toplevel_execute_ctrl3_down_Decode_STORE_ID_lane0 = toplevel_execute_ctrl3_up_Decode_STORE_ID_lane0;
  assign toplevel_execute_ctrl3_down_LsuPlugin_logic_FROM_LSU_lane0 = toplevel_execute_ctrl3_up_LsuPlugin_logic_FROM_LSU_lane0;
  assign toplevel_execute_ctrl3_down_LsuPlugin_logic_FROM_PREFETCH_lane0 = toplevel_execute_ctrl3_up_LsuPlugin_logic_FROM_PREFETCH_lane0;
  assign toplevel_execute_ctrl4_up_ready = toplevel_execute_ctrl4_down_isReady;
  assign toplevel_execute_ctrl4_down_Decode_UOP_lane0 = toplevel_execute_ctrl4_up_Decode_UOP_lane0;
  assign toplevel_execute_ctrl4_down_Prediction_ALIGNED_JUMPED_lane0 = toplevel_execute_ctrl4_up_Prediction_ALIGNED_JUMPED_lane0;
  assign toplevel_execute_ctrl4_down_Prediction_ALIGNED_JUMPED_PC_lane0 = toplevel_execute_ctrl4_up_Prediction_ALIGNED_JUMPED_PC_lane0;
  assign toplevel_execute_ctrl4_down_Prediction_ALIGNED_SLICES_TAKEN_lane0 = toplevel_execute_ctrl4_up_Prediction_ALIGNED_SLICES_TAKEN_lane0;
  assign toplevel_execute_ctrl4_down_Prediction_ALIGNED_SLICES_BRANCH_lane0 = toplevel_execute_ctrl4_up_Prediction_ALIGNED_SLICES_BRANCH_lane0;
  assign toplevel_execute_ctrl4_down_GSharePlugin_GSHARE_COUNTER_lane0_0 = toplevel_execute_ctrl4_up_GSharePlugin_GSHARE_COUNTER_lane0_0;
  assign toplevel_execute_ctrl4_down_GSharePlugin_GSHARE_COUNTER_lane0_1 = toplevel_execute_ctrl4_up_GSharePlugin_GSHARE_COUNTER_lane0_1;
  assign toplevel_execute_ctrl4_down_GSharePlugin_GSHARE_COUNTER_lane0_2 = toplevel_execute_ctrl4_up_GSharePlugin_GSHARE_COUNTER_lane0_2;
  assign toplevel_execute_ctrl4_down_GSharePlugin_GSHARE_COUNTER_lane0_3 = toplevel_execute_ctrl4_up_GSharePlugin_GSHARE_COUNTER_lane0_3;
  assign toplevel_execute_ctrl4_down_Prediction_BRANCH_HISTORY_lane0 = toplevel_execute_ctrl4_up_Prediction_BRANCH_HISTORY_lane0;
  assign toplevel_execute_ctrl4_down_Decode_INSTRUCTION_SLICE_COUNT_lane0 = toplevel_execute_ctrl4_up_Decode_INSTRUCTION_SLICE_COUNT_lane0;
  assign toplevel_execute_ctrl4_down_PC_lane0 = toplevel_execute_ctrl4_up_PC_lane0;
  assign toplevel_execute_ctrl4_down_Decode_UOP_ID_lane0 = toplevel_execute_ctrl4_up_Decode_UOP_ID_lane0;
  assign toplevel_execute_ctrl4_down_RD_PHYS_lane0 = toplevel_execute_ctrl4_up_RD_PHYS_lane0;
  assign toplevel_execute_ctrl4_down_LANE_AGE_lane0 = toplevel_execute_ctrl4_up_LANE_AGE_lane0;
  assign toplevel_execute_ctrl4_down_Decode_UOP_lane1 = toplevel_execute_ctrl4_up_Decode_UOP_lane1;
  assign toplevel_execute_ctrl4_down_Prediction_ALIGNED_JUMPED_lane1 = toplevel_execute_ctrl4_up_Prediction_ALIGNED_JUMPED_lane1;
  assign toplevel_execute_ctrl4_down_Prediction_ALIGNED_JUMPED_PC_lane1 = toplevel_execute_ctrl4_up_Prediction_ALIGNED_JUMPED_PC_lane1;
  assign toplevel_execute_ctrl4_down_Prediction_ALIGNED_SLICES_TAKEN_lane1 = toplevel_execute_ctrl4_up_Prediction_ALIGNED_SLICES_TAKEN_lane1;
  assign toplevel_execute_ctrl4_down_Prediction_ALIGNED_SLICES_BRANCH_lane1 = toplevel_execute_ctrl4_up_Prediction_ALIGNED_SLICES_BRANCH_lane1;
  assign toplevel_execute_ctrl4_down_GSharePlugin_GSHARE_COUNTER_lane1_0 = toplevel_execute_ctrl4_up_GSharePlugin_GSHARE_COUNTER_lane1_0;
  assign toplevel_execute_ctrl4_down_GSharePlugin_GSHARE_COUNTER_lane1_1 = toplevel_execute_ctrl4_up_GSharePlugin_GSHARE_COUNTER_lane1_1;
  assign toplevel_execute_ctrl4_down_GSharePlugin_GSHARE_COUNTER_lane1_2 = toplevel_execute_ctrl4_up_GSharePlugin_GSHARE_COUNTER_lane1_2;
  assign toplevel_execute_ctrl4_down_GSharePlugin_GSHARE_COUNTER_lane1_3 = toplevel_execute_ctrl4_up_GSharePlugin_GSHARE_COUNTER_lane1_3;
  assign toplevel_execute_ctrl4_down_Prediction_BRANCH_HISTORY_lane1 = toplevel_execute_ctrl4_up_Prediction_BRANCH_HISTORY_lane1;
  assign toplevel_execute_ctrl4_down_Decode_INSTRUCTION_SLICE_COUNT_lane1 = toplevel_execute_ctrl4_up_Decode_INSTRUCTION_SLICE_COUNT_lane1;
  assign toplevel_execute_ctrl4_down_PC_lane1 = toplevel_execute_ctrl4_up_PC_lane1;
  assign toplevel_execute_ctrl4_down_TRAP_lane1 = toplevel_execute_ctrl4_up_TRAP_lane1;
  assign toplevel_execute_ctrl4_down_Decode_UOP_ID_lane1 = toplevel_execute_ctrl4_up_Decode_UOP_ID_lane1;
  assign toplevel_execute_ctrl4_down_RD_PHYS_lane1 = toplevel_execute_ctrl4_up_RD_PHYS_lane1;
  assign toplevel_execute_ctrl4_down_LANE_AGE_lane1 = toplevel_execute_ctrl4_up_LANE_AGE_lane1;
  assign toplevel_execute_ctrl4_down_AguPlugin_SIZE_lane0 = toplevel_execute_ctrl4_up_AguPlugin_SIZE_lane0;
  assign toplevel_execute_ctrl4_down_integer_RS2_lane0 = toplevel_execute_ctrl4_up_integer_RS2_lane0;
  assign toplevel_execute_ctrl4_down_early0_BranchPlugin_SEL_lane0 = toplevel_execute_ctrl4_up_early0_BranchPlugin_SEL_lane0;
  assign toplevel_execute_ctrl4_down_early0_MulPlugin_SEL_lane0 = toplevel_execute_ctrl4_up_early0_MulPlugin_SEL_lane0;
  assign toplevel_execute_ctrl4_down_late0_IntAluPlugin_SEL_lane0 = toplevel_execute_ctrl4_up_late0_IntAluPlugin_SEL_lane0;
  assign toplevel_execute_ctrl4_down_late0_BarrelShifterPlugin_SEL_lane0 = toplevel_execute_ctrl4_up_late0_BarrelShifterPlugin_SEL_lane0;
  assign toplevel_execute_ctrl4_down_late0_BranchPlugin_SEL_lane0 = toplevel_execute_ctrl4_up_late0_BranchPlugin_SEL_lane0;
  assign toplevel_execute_ctrl4_down_MulPlugin_HIGH_lane0 = toplevel_execute_ctrl4_up_MulPlugin_HIGH_lane0;
  assign toplevel_execute_ctrl4_down_AguPlugin_SEL_lane0 = toplevel_execute_ctrl4_up_AguPlugin_SEL_lane0;
  assign toplevel_execute_ctrl4_down_LsuPlugin_logic_FENCE_lane0 = toplevel_execute_ctrl4_up_LsuPlugin_logic_FENCE_lane0;
  assign toplevel_execute_ctrl4_down_lane0_integer_WriteBackPlugin_SEL_lane0 = toplevel_execute_ctrl4_up_lane0_integer_WriteBackPlugin_SEL_lane0;
  assign toplevel_execute_ctrl4_down_COMPLETION_AT_4_lane0 = toplevel_execute_ctrl4_up_COMPLETION_AT_4_lane0;
  assign toplevel_execute_ctrl4_down_execute_lane0_logic_completions_onCtrl_2_ENABLE_lane0 = toplevel_execute_ctrl4_up_execute_lane0_logic_completions_onCtrl_2_ENABLE_lane0;
  assign toplevel_execute_ctrl4_down_SrcStageables_REVERT_lane0 = toplevel_execute_ctrl4_up_SrcStageables_REVERT_lane0;
  assign toplevel_execute_ctrl4_down_SrcStageables_ZERO_lane0 = toplevel_execute_ctrl4_up_SrcStageables_ZERO_lane0;
  assign toplevel_execute_ctrl4_down_lane0_IntFormatPlugin_logic_SIGNED_lane0 = toplevel_execute_ctrl4_up_lane0_IntFormatPlugin_logic_SIGNED_lane0;
  assign toplevel_execute_ctrl4_down_lane0_IntFormatPlugin_logic_WIDTH_ID_lane0 = toplevel_execute_ctrl4_up_lane0_IntFormatPlugin_logic_WIDTH_ID_lane0;
  assign toplevel_execute_ctrl4_down_SrcStageables_UNSIGNED_lane0 = toplevel_execute_ctrl4_up_SrcStageables_UNSIGNED_lane0;
  assign toplevel_execute_ctrl4_down_BarrelShifterPlugin_LEFT_lane0 = toplevel_execute_ctrl4_up_BarrelShifterPlugin_LEFT_lane0;
  assign toplevel_execute_ctrl4_down_BarrelShifterPlugin_SIGNED_lane0 = toplevel_execute_ctrl4_up_BarrelShifterPlugin_SIGNED_lane0;
  assign toplevel_execute_ctrl4_down_BranchPlugin_BRANCH_CTRL_lane0 = toplevel_execute_ctrl4_up_BranchPlugin_BRANCH_CTRL_lane0;
  assign toplevel_execute_ctrl4_down_AguPlugin_LOAD_lane0 = toplevel_execute_ctrl4_up_AguPlugin_LOAD_lane0;
  assign toplevel_execute_ctrl4_down_AguPlugin_STORE_lane0 = toplevel_execute_ctrl4_up_AguPlugin_STORE_lane0;
  assign toplevel_execute_ctrl4_down_AguPlugin_ATOMIC_lane0 = toplevel_execute_ctrl4_up_AguPlugin_ATOMIC_lane0;
  assign toplevel_execute_ctrl4_down_AguPlugin_FLOAT_lane0 = toplevel_execute_ctrl4_up_AguPlugin_FLOAT_lane0;
  assign toplevel_execute_ctrl4_down_LsuPlugin_logic_LSU_PREFETCH_lane0 = toplevel_execute_ctrl4_up_LsuPlugin_logic_LSU_PREFETCH_lane0;
  assign toplevel_execute_ctrl4_down_late0_IntAluPlugin_ALU_ADD_SUB_lane0 = toplevel_execute_ctrl4_up_late0_IntAluPlugin_ALU_ADD_SUB_lane0;
  assign toplevel_execute_ctrl4_down_late0_IntAluPlugin_ALU_SLTX_lane0 = toplevel_execute_ctrl4_up_late0_IntAluPlugin_ALU_SLTX_lane0;
  assign toplevel_execute_ctrl4_down_late0_IntAluPlugin_ALU_BITWISE_CTRL_lane0 = toplevel_execute_ctrl4_up_late0_IntAluPlugin_ALU_BITWISE_CTRL_lane0;
  assign toplevel_execute_ctrl4_down_early1_BranchPlugin_SEL_lane1 = toplevel_execute_ctrl4_up_early1_BranchPlugin_SEL_lane1;
  assign toplevel_execute_ctrl4_down_late1_IntAluPlugin_SEL_lane1 = toplevel_execute_ctrl4_up_late1_IntAluPlugin_SEL_lane1;
  assign toplevel_execute_ctrl4_down_late1_BarrelShifterPlugin_SEL_lane1 = toplevel_execute_ctrl4_up_late1_BarrelShifterPlugin_SEL_lane1;
  assign toplevel_execute_ctrl4_down_late1_BranchPlugin_SEL_lane1 = toplevel_execute_ctrl4_up_late1_BranchPlugin_SEL_lane1;
  assign toplevel_execute_ctrl4_down_lane1_integer_WriteBackPlugin_SEL_lane1 = toplevel_execute_ctrl4_up_lane1_integer_WriteBackPlugin_SEL_lane1;
  assign toplevel_execute_ctrl4_down_COMPLETION_AT_4_lane1 = toplevel_execute_ctrl4_up_COMPLETION_AT_4_lane1;
  assign toplevel_execute_ctrl4_down_execute_lane1_logic_completions_onCtrl_2_ENABLE_lane1 = toplevel_execute_ctrl4_up_execute_lane1_logic_completions_onCtrl_2_ENABLE_lane1;
  assign toplevel_execute_ctrl4_down_SrcStageables_REVERT_lane1 = toplevel_execute_ctrl4_up_SrcStageables_REVERT_lane1;
  assign toplevel_execute_ctrl4_down_SrcStageables_ZERO_lane1 = toplevel_execute_ctrl4_up_SrcStageables_ZERO_lane1;
  assign toplevel_execute_ctrl4_down_SrcStageables_UNSIGNED_lane1 = toplevel_execute_ctrl4_up_SrcStageables_UNSIGNED_lane1;
  assign toplevel_execute_ctrl4_down_BarrelShifterPlugin_LEFT_lane1 = toplevel_execute_ctrl4_up_BarrelShifterPlugin_LEFT_lane1;
  assign toplevel_execute_ctrl4_down_BarrelShifterPlugin_SIGNED_lane1 = toplevel_execute_ctrl4_up_BarrelShifterPlugin_SIGNED_lane1;
  assign toplevel_execute_ctrl4_down_BranchPlugin_BRANCH_CTRL_lane1 = toplevel_execute_ctrl4_up_BranchPlugin_BRANCH_CTRL_lane1;
  assign toplevel_execute_ctrl4_down_late1_IntAluPlugin_ALU_ADD_SUB_lane1 = toplevel_execute_ctrl4_up_late1_IntAluPlugin_ALU_ADD_SUB_lane1;
  assign toplevel_execute_ctrl4_down_late1_IntAluPlugin_ALU_SLTX_lane1 = toplevel_execute_ctrl4_up_late1_IntAluPlugin_ALU_SLTX_lane1;
  assign toplevel_execute_ctrl4_down_late1_IntAluPlugin_ALU_BITWISE_CTRL_lane1 = toplevel_execute_ctrl4_up_late1_IntAluPlugin_ALU_BITWISE_CTRL_lane1;
  assign toplevel_execute_ctrl4_down_COMMIT_lane1 = toplevel_execute_ctrl4_up_COMMIT_lane1;
  assign toplevel_execute_ctrl4_down_early0_BranchPlugin_pcCalc_PC_TRUE_lane0 = toplevel_execute_ctrl4_up_early0_BranchPlugin_pcCalc_PC_TRUE_lane0;
  assign toplevel_execute_ctrl4_down_early0_BranchPlugin_pcCalc_PC_FALSE_lane0 = toplevel_execute_ctrl4_up_early0_BranchPlugin_pcCalc_PC_FALSE_lane0;
  assign toplevel_execute_ctrl4_down_early0_BranchPlugin_pcCalc_PC_LAST_SLICE_lane0 = toplevel_execute_ctrl4_up_early0_BranchPlugin_pcCalc_PC_LAST_SLICE_lane0;
  assign toplevel_execute_ctrl4_down_early1_BranchPlugin_pcCalc_PC_TRUE_lane1 = toplevel_execute_ctrl4_up_early1_BranchPlugin_pcCalc_PC_TRUE_lane1;
  assign toplevel_execute_ctrl4_down_early1_BranchPlugin_pcCalc_PC_FALSE_lane1 = toplevel_execute_ctrl4_up_early1_BranchPlugin_pcCalc_PC_FALSE_lane1;
  assign toplevel_execute_ctrl4_down_early1_BranchPlugin_pcCalc_PC_LAST_SLICE_lane1 = toplevel_execute_ctrl4_up_early1_BranchPlugin_pcCalc_PC_LAST_SLICE_lane1;
  assign toplevel_execute_ctrl4_down_LsuL1_MIXED_ADDRESS_lane0 = toplevel_execute_ctrl4_up_LsuL1_MIXED_ADDRESS_lane0;
  assign toplevel_execute_ctrl4_down_LsuL1Plugin_logic_EVENT_WRITE_DATA_lane0 = toplevel_execute_ctrl4_up_LsuL1Plugin_logic_EVENT_WRITE_DATA_lane0;
  assign toplevel_execute_ctrl4_down_LsuL1Plugin_logic_EVENT_WRITE_MASK_lane0 = toplevel_execute_ctrl4_up_LsuL1Plugin_logic_EVENT_WRITE_MASK_lane0;
  assign toplevel_execute_ctrl4_down_LsuPlugin_logic_FROM_ACCESS_lane0 = toplevel_execute_ctrl4_up_LsuPlugin_logic_FROM_ACCESS_lane0;
  assign toplevel_execute_ctrl4_down_LsuL1_MASK_lane0 = toplevel_execute_ctrl4_up_LsuL1_MASK_lane0;
  assign toplevel_execute_ctrl4_down_LsuL1_SIZE_lane0 = toplevel_execute_ctrl4_up_LsuL1_SIZE_lane0;
  assign toplevel_execute_ctrl4_down_LsuL1_LOAD_lane0 = toplevel_execute_ctrl4_up_LsuL1_LOAD_lane0;
  assign toplevel_execute_ctrl4_down_LsuL1_ATOMIC_lane0 = toplevel_execute_ctrl4_up_LsuL1_ATOMIC_lane0;
  assign toplevel_execute_ctrl4_down_LsuL1_STORE_lane0 = toplevel_execute_ctrl4_up_LsuL1_STORE_lane0;
  assign toplevel_execute_ctrl4_down_LsuL1_PREFETCH_lane0 = toplevel_execute_ctrl4_up_LsuL1_PREFETCH_lane0;
  assign toplevel_execute_ctrl4_down_LsuL1_FLUSH_lane0 = toplevel_execute_ctrl4_up_LsuL1_FLUSH_lane0;
  assign toplevel_execute_ctrl4_down_Decode_STORE_ID_lane0 = toplevel_execute_ctrl4_up_Decode_STORE_ID_lane0;
  assign toplevel_execute_ctrl4_down_LsuPlugin_logic_FROM_LSU_lane0 = toplevel_execute_ctrl4_up_LsuPlugin_logic_FROM_LSU_lane0;
  assign toplevel_execute_ctrl4_down_LsuPlugin_logic_FROM_PREFETCH_lane0 = toplevel_execute_ctrl4_up_LsuPlugin_logic_FROM_PREFETCH_lane0;
  assign toplevel_execute_ctrl4_down_LsuL1Plugin_logic_SHARED_lane0_plru_0 = toplevel_execute_ctrl4_up_LsuL1Plugin_logic_SHARED_lane0_plru_0;
  assign toplevel_execute_ctrl4_down_LsuL1Plugin_logic_SHARED_lane0_dirty = toplevel_execute_ctrl4_up_LsuL1Plugin_logic_SHARED_lane0_dirty;
  assign toplevel_execute_ctrl4_down_early0_MulPlugin_logic_steps_0_adders_0_lane0 = toplevel_execute_ctrl4_up_early0_MulPlugin_logic_steps_0_adders_0_lane0;
  assign toplevel_execute_ctrl4_down_early0_MulPlugin_logic_steps_0_adders_1_lane0 = toplevel_execute_ctrl4_up_early0_MulPlugin_logic_steps_0_adders_1_lane0;
  assign toplevel_execute_ctrl4_down_late0_SrcPlugin_SRC1_lane0 = toplevel_execute_ctrl4_up_late0_SrcPlugin_SRC1_lane0;
  assign toplevel_execute_ctrl4_down_late0_SrcPlugin_SRC2_lane0 = toplevel_execute_ctrl4_up_late0_SrcPlugin_SRC2_lane0;
  assign toplevel_execute_ctrl4_down_late1_SrcPlugin_SRC1_lane1 = toplevel_execute_ctrl4_up_late1_SrcPlugin_SRC1_lane1;
  assign toplevel_execute_ctrl4_down_late1_SrcPlugin_SRC2_lane1 = toplevel_execute_ctrl4_up_late1_SrcPlugin_SRC2_lane1;
  assign toplevel_execute_ctrl4_down_LsuL1Plugin_logic_BANK_BUSY_REMAPPED_lane0 = toplevel_execute_ctrl4_up_LsuL1Plugin_logic_BANK_BUSY_REMAPPED_lane0;
  assign toplevel_execute_ctrl4_down_LsuL1Plugin_logic_BANKS_MUXES_lane0_0 = toplevel_execute_ctrl4_up_LsuL1Plugin_logic_BANKS_MUXES_lane0_0;
  assign toplevel_execute_ctrl4_down_LsuL1Plugin_logic_BANKS_MUXES_lane0_1 = toplevel_execute_ctrl4_up_LsuL1Plugin_logic_BANKS_MUXES_lane0_1;
  assign toplevel_execute_ctrl4_down_LsuL1Plugin_logic_WRITE_TO_READ_HAZARDS_lane0 = toplevel_execute_ctrl4_up_LsuL1Plugin_logic_WRITE_TO_READ_HAZARDS_lane0;
  assign toplevel_execute_ctrl4_down_LsuL1_PHYSICAL_ADDRESS_lane0 = toplevel_execute_ctrl4_up_LsuL1_PHYSICAL_ADDRESS_lane0;
  assign toplevel_execute_ctrl4_down_LsuL1Plugin_logic_WAYS_TAGS_lane0_0_loaded = toplevel_execute_ctrl4_up_LsuL1Plugin_logic_WAYS_TAGS_lane0_0_loaded;
  assign toplevel_execute_ctrl4_down_LsuL1Plugin_logic_WAYS_TAGS_lane0_0_address = toplevel_execute_ctrl4_up_LsuL1Plugin_logic_WAYS_TAGS_lane0_0_address;
  assign toplevel_execute_ctrl4_down_LsuL1Plugin_logic_WAYS_TAGS_lane0_0_fault = toplevel_execute_ctrl4_up_LsuL1Plugin_logic_WAYS_TAGS_lane0_0_fault;
  assign toplevel_execute_ctrl4_down_LsuL1Plugin_logic_WAYS_TAGS_lane0_1_loaded = toplevel_execute_ctrl4_up_LsuL1Plugin_logic_WAYS_TAGS_lane0_1_loaded;
  assign toplevel_execute_ctrl4_down_LsuL1Plugin_logic_WAYS_TAGS_lane0_1_address = toplevel_execute_ctrl4_up_LsuL1Plugin_logic_WAYS_TAGS_lane0_1_address;
  assign toplevel_execute_ctrl4_down_LsuL1Plugin_logic_WAYS_TAGS_lane0_1_fault = toplevel_execute_ctrl4_up_LsuL1Plugin_logic_WAYS_TAGS_lane0_1_fault;
  assign toplevel_execute_ctrl4_down_LsuL1Plugin_logic_WAYS_HITS_lane0 = toplevel_execute_ctrl4_up_LsuL1Plugin_logic_WAYS_HITS_lane0;
  assign toplevel_execute_ctrl4_down_LsuPlugin_logic_onTrigger_HIT_lane0 = toplevel_execute_ctrl4_up_LsuPlugin_logic_onTrigger_HIT_lane0;
  assign toplevel_execute_ctrl4_down_MMU_TRANSLATED_lane0 = toplevel_execute_ctrl4_up_MMU_TRANSLATED_lane0;
  assign toplevel_execute_ctrl4_down_LsuPlugin_logic_preCtrl_MISS_ALIGNED_lane0 = toplevel_execute_ctrl4_up_LsuPlugin_logic_preCtrl_MISS_ALIGNED_lane0;
  assign toplevel_execute_ctrl4_down_LsuPlugin_logic_preCtrl_IS_AMO_lane0 = toplevel_execute_ctrl4_up_LsuPlugin_logic_preCtrl_IS_AMO_lane0;
  assign toplevel_execute_ctrl4_down_LsuPlugin_logic_onPma_CACHED_RSP_lane0_fault = toplevel_execute_ctrl4_up_LsuPlugin_logic_onPma_CACHED_RSP_lane0_fault;
  assign toplevel_execute_ctrl4_down_LsuPlugin_logic_onPma_CACHED_RSP_lane0_io = toplevel_execute_ctrl4_up_LsuPlugin_logic_onPma_CACHED_RSP_lane0_io;
  assign toplevel_execute_ctrl4_down_LsuPlugin_logic_onPma_IO_RSP_lane0_fault = toplevel_execute_ctrl4_up_LsuPlugin_logic_onPma_IO_RSP_lane0_fault;
  assign toplevel_execute_ctrl4_down_LsuPlugin_logic_onPma_IO_RSP_lane0_io = toplevel_execute_ctrl4_up_LsuPlugin_logic_onPma_IO_RSP_lane0_io;
  assign toplevel_execute_ctrl4_down_LsuPlugin_logic_onPma_IO_lane0 = toplevel_execute_ctrl4_up_LsuPlugin_logic_onPma_IO_lane0;
  assign toplevel_execute_ctrl4_down_LsuPlugin_logic_onPma_FROM_LSU_MSB_FAILED_lane0 = toplevel_execute_ctrl4_up_LsuPlugin_logic_onPma_FROM_LSU_MSB_FAILED_lane0;
  assign toplevel_execute_ctrl4_down_LsuPlugin_logic_MMU_PAGE_FAULT_lane0 = toplevel_execute_ctrl4_up_LsuPlugin_logic_MMU_PAGE_FAULT_lane0;
  assign toplevel_execute_ctrl4_down_LsuPlugin_logic_MMU_FAILURE_lane0 = toplevel_execute_ctrl4_up_LsuPlugin_logic_MMU_FAILURE_lane0;
  assign toplevel_execute_ctrl4_down_MMU_ACCESS_FAULT_lane0 = toplevel_execute_ctrl4_up_MMU_ACCESS_FAULT_lane0;
  assign toplevel_execute_ctrl4_down_MMU_REFILL_lane0 = toplevel_execute_ctrl4_up_MMU_REFILL_lane0;
  assign toplevel_execute_ctrl4_down_MMU_HAZARD_lane0 = toplevel_execute_ctrl4_up_MMU_HAZARD_lane0;
  assign toplevel_execute_ctrl4_down_MMU_BYPASS_TRANSLATION_lane0 = toplevel_execute_ctrl4_up_MMU_BYPASS_TRANSLATION_lane0;
  assign toplevel_execute_ctrl5_up_ready = toplevel_execute_ctrl5_down_isReady;
  assign toplevel_execute_ctrl5_down_LANE_SEL_lane0 = toplevel_execute_ctrl5_up_LANE_SEL_lane0;
  assign toplevel_execute_ctrl5_down_RD_PHYS_lane0 = toplevel_execute_ctrl5_up_RD_PHYS_lane0;
  assign toplevel_execute_ctrl5_down_LANE_AGE_lane0 = toplevel_execute_ctrl5_up_LANE_AGE_lane0;
  assign toplevel_execute_ctrl5_down_LANE_SEL_lane1 = toplevel_execute_ctrl5_up_LANE_SEL_lane1;
  assign toplevel_execute_ctrl5_down_RD_PHYS_lane1 = toplevel_execute_ctrl5_up_RD_PHYS_lane1;
  assign toplevel_execute_ctrl5_down_LANE_AGE_lane1 = toplevel_execute_ctrl5_up_LANE_AGE_lane1;
  assign toplevel_execute_ctrl5_down_COMMIT_lane0 = toplevel_execute_ctrl5_up_COMMIT_lane0;
  assign toplevel_execute_ctrl5_down_COMMIT_lane1 = toplevel_execute_ctrl5_up_COMMIT_lane1;
  assign toplevel_execute_ctrl5_down_lane0_integer_WriteBackPlugin_logic_DATA_lane0 = toplevel_execute_ctrl5_up_lane0_integer_WriteBackPlugin_logic_DATA_lane0;
  assign toplevel_execute_ctrl5_down_lane1_integer_WriteBackPlugin_logic_DATA_lane1 = toplevel_execute_ctrl5_up_lane1_integer_WriteBackPlugin_logic_DATA_lane1;
  assign fetch_logic_ctrls_0_down_isFiring = (fetch_logic_ctrls_0_down_isValid && fetch_logic_ctrls_0_down_isReady);
  assign fetch_logic_ctrls_0_down_isValid = fetch_logic_ctrls_0_down_valid;
  assign fetch_logic_ctrls_0_down_isReady = fetch_logic_ctrls_0_down_ready;
  assign fetch_logic_ctrls_1_up_isValid = fetch_logic_ctrls_1_up_valid;
  assign fetch_logic_ctrls_1_down_isValid = fetch_logic_ctrls_1_down_valid;
  assign fetch_logic_ctrls_1_down_isReady = fetch_logic_ctrls_1_down_ready;
  assign fetch_logic_ctrls_2_up_isValid = fetch_logic_ctrls_2_up_valid;
  assign fetch_logic_ctrls_2_up_isReady = fetch_logic_ctrls_2_up_ready;
  assign fetch_logic_ctrls_2_up_isCancel = fetch_logic_ctrls_2_up_cancel;
  assign fetch_logic_ctrls_2_up_isCanceling = (fetch_logic_ctrls_2_up_isValid && fetch_logic_ctrls_2_up_isCancel);
  assign fetch_logic_ctrls_0_up_isFiring = (fetch_logic_ctrls_0_up_isValid && fetch_logic_ctrls_0_up_isReady);
  assign fetch_logic_ctrls_0_up_isValid = fetch_logic_ctrls_0_up_valid;
  assign fetch_logic_ctrls_0_up_isReady = fetch_logic_ctrls_0_up_ready;
  assign fetch_logic_ctrls_2_down_isValid = fetch_logic_ctrls_2_down_valid;
  assign fetch_logic_ctrls_2_down_isReady = fetch_logic_ctrls_2_down_ready;
  assign fetch_logic_ctrls_2_down_isCancel = 1'b0;
  assign toplevel_decode_ctrls_0_down_isValid = toplevel_decode_ctrls_0_down_valid;
  assign toplevel_decode_ctrls_0_down_isReady = toplevel_decode_ctrls_0_down_ready;
  assign toplevel_decode_ctrls_1_up_isMoving = (toplevel_decode_ctrls_1_up_isValid && toplevel_decode_ctrls_1_up_isReady);
  assign toplevel_decode_ctrls_1_up_isValid = toplevel_decode_ctrls_1_up_valid;
  assign toplevel_decode_ctrls_1_up_isReady = toplevel_decode_ctrls_1_up_ready;
  assign toplevel_decode_ctrls_1_up_isCanceling = 1'b0;
  assign toplevel_decode_ctrls_0_up_isFiring = (toplevel_decode_ctrls_0_up_isValid && toplevel_decode_ctrls_0_up_isReady);
  assign toplevel_decode_ctrls_0_up_isMoving = (toplevel_decode_ctrls_0_up_isValid && toplevel_decode_ctrls_0_up_isReady);
  assign toplevel_decode_ctrls_0_up_isValid = toplevel_decode_ctrls_0_up_valid;
  assign toplevel_decode_ctrls_0_up_isReady = toplevel_decode_ctrls_0_up_ready;
  assign toplevel_decode_ctrls_0_up_isCancel = 1'b0;
  assign toplevel_decode_ctrls_1_down_isReady = toplevel_decode_ctrls_1_down_ready;
  assign toplevel_execute_ctrl0_down_isReady = toplevel_execute_ctrl0_down_ready;
  assign toplevel_execute_ctrl1_down_isReady = toplevel_execute_ctrl1_down_ready;
  assign toplevel_execute_ctrl2_down_isReady = toplevel_execute_ctrl2_down_ready;
  assign toplevel_execute_ctrl3_down_isReady = toplevel_execute_ctrl3_down_ready;
  assign toplevel_execute_ctrl4_down_isReady = toplevel_execute_ctrl4_down_ready;
  assign toplevel_execute_ctrl5_down_isReady = toplevel_execute_ctrl5_down_ready;
  always @(*) begin
    LsuPlugin_logic_flusher_stateNext = LsuPlugin_logic_flusher_stateReg;
    case(LsuPlugin_logic_flusher_stateReg)
      LsuPlugin_logic_flusher_enumDef_CMD : begin
        if(when_LsuPlugin_l297) begin
          LsuPlugin_logic_flusher_stateNext = LsuPlugin_logic_flusher_enumDef_COMPLETION;
        end
      end
      LsuPlugin_logic_flusher_enumDef_COMPLETION : begin
        if(when_LsuPlugin_l305) begin
          LsuPlugin_logic_flusher_stateNext = LsuPlugin_logic_flusher_enumDef_IDLE;
        end
      end
      default : begin
        if(LsuPlugin_logic_flusher_arbiter_io_output_valid) begin
          LsuPlugin_logic_flusher_stateNext = LsuPlugin_logic_flusher_enumDef_CMD;
        end
      end
    endcase
    if(LsuPlugin_logic_flusher_wantKill) begin
      LsuPlugin_logic_flusher_stateNext = LsuPlugin_logic_flusher_enumDef_IDLE;
    end
  end

  assign when_LsuPlugin_l297 = (LsuPlugin_logic_flusher_cmdCounter[6] && (! LsuPlugin_logic_flusher_inflight));
  assign when_LsuPlugin_l305 = (! (|LsuPlugin_logic_flusher_waiter));
  always @(*) begin
    TrapPlugin_logic_harts_0_trap_fsm_stateNext = TrapPlugin_logic_harts_0_trap_fsm_stateReg;
    case(TrapPlugin_logic_harts_0_trap_fsm_stateReg)
      TrapPlugin_logic_harts_0_trap_fsm_enumDef_RUNNING : begin
        if(TrapPlugin_logic_harts_0_trap_trigger_valid) begin
          TrapPlugin_logic_harts_0_trap_fsm_stateNext = TrapPlugin_logic_harts_0_trap_fsm_enumDef_PROCESS_1;
        end
      end
      TrapPlugin_logic_harts_0_trap_fsm_enumDef_PROCESS_1 : begin
        if(when_TrapPlugin_l393) begin
          TrapPlugin_logic_harts_0_trap_fsm_stateNext = TrapPlugin_logic_harts_0_trap_fsm_enumDef_TRAP_TVAL;
        end else begin
          case(TrapPlugin_logic_harts_0_trap_pending_state_code)
            4'b0000 : begin
              TrapPlugin_logic_harts_0_trap_fsm_stateNext = TrapPlugin_logic_harts_0_trap_fsm_enumDef_RUNNING;
            end
            4'b0001 : begin
              TrapPlugin_logic_harts_0_trap_fsm_stateNext = TrapPlugin_logic_harts_0_trap_fsm_enumDef_XRET_EPC;
            end
            4'b0010 : begin
              TrapPlugin_logic_harts_0_trap_fsm_stateNext = TrapPlugin_logic_harts_0_trap_fsm_enumDef_LSU_FLUSH;
            end
            4'b0100 : begin
              TrapPlugin_logic_harts_0_trap_fsm_stateNext = TrapPlugin_logic_harts_0_trap_fsm_enumDef_JUMP;
            end
            4'b0101 : begin
              TrapPlugin_logic_harts_0_trap_fsm_stateNext = TrapPlugin_logic_harts_0_trap_fsm_enumDef_JUMP;
            end
            4'b1000 : begin
              if(TrapPlugin_api_harts_0_askWake) begin
                TrapPlugin_logic_harts_0_trap_fsm_stateNext = TrapPlugin_logic_harts_0_trap_fsm_enumDef_JUMP;
              end
            end
            4'b0110 : begin
              if(TrapPlugin_logic_harts_0_trap_fsm_atsPorts_invalidate_cmd_ready) begin
                TrapPlugin_logic_harts_0_trap_fsm_stateNext = TrapPlugin_logic_harts_0_trap_fsm_enumDef_JUMP;
              end
            end
            4'b0111 : begin
              if(TrapPlugin_logic_harts_0_trap_fsm_atsPorts_refill_cmd_ready) begin
                TrapPlugin_logic_harts_0_trap_fsm_stateNext = TrapPlugin_logic_harts_0_trap_fsm_enumDef_ATS_RSP;
              end
            end
            default : begin
            end
          endcase
        end
      end
      TrapPlugin_logic_harts_0_trap_fsm_enumDef_TRAP_EPC : begin
        if(TrapPlugin_logic_harts_0_crsPorts_write_ready) begin
          TrapPlugin_logic_harts_0_trap_fsm_stateNext = TrapPlugin_logic_harts_0_trap_fsm_enumDef_TRAP_TVEC;
        end
      end
      TrapPlugin_logic_harts_0_trap_fsm_enumDef_TRAP_TVAL : begin
        if(TrapPlugin_logic_harts_0_crsPorts_write_ready) begin
          TrapPlugin_logic_harts_0_trap_fsm_stateNext = TrapPlugin_logic_harts_0_trap_fsm_enumDef_TRAP_EPC;
        end
      end
      TrapPlugin_logic_harts_0_trap_fsm_enumDef_TRAP_TVEC : begin
        if(TrapPlugin_logic_harts_0_crsPorts_read_ready) begin
          TrapPlugin_logic_harts_0_trap_fsm_stateNext = TrapPlugin_logic_harts_0_trap_fsm_enumDef_TRAP_APPLY;
        end
      end
      TrapPlugin_logic_harts_0_trap_fsm_enumDef_TRAP_APPLY : begin
        TrapPlugin_logic_harts_0_trap_fsm_stateNext = TrapPlugin_logic_harts_0_trap_fsm_enumDef_RUNNING;
      end
      TrapPlugin_logic_harts_0_trap_fsm_enumDef_XRET_EPC : begin
        if(TrapPlugin_logic_harts_0_crsPorts_read_ready) begin
          TrapPlugin_logic_harts_0_trap_fsm_stateNext = TrapPlugin_logic_harts_0_trap_fsm_enumDef_XRET_APPLY;
        end
      end
      TrapPlugin_logic_harts_0_trap_fsm_enumDef_XRET_APPLY : begin
        TrapPlugin_logic_harts_0_trap_fsm_stateNext = TrapPlugin_logic_harts_0_trap_fsm_enumDef_RUNNING;
      end
      TrapPlugin_logic_harts_0_trap_fsm_enumDef_ATS_RSP : begin
        if(TrapPlugin_logic_harts_0_trap_fsm_atsPorts_refill_rsp_valid) begin
          TrapPlugin_logic_harts_0_trap_fsm_stateNext = TrapPlugin_logic_harts_0_trap_fsm_enumDef_JUMP;
          if(when_TrapPlugin_l492) begin
            TrapPlugin_logic_harts_0_trap_fsm_stateNext = TrapPlugin_logic_harts_0_trap_fsm_enumDef_TRAP_TVAL;
          end
        end
      end
      TrapPlugin_logic_harts_0_trap_fsm_enumDef_JUMP : begin
        TrapPlugin_logic_harts_0_trap_fsm_stateNext = TrapPlugin_logic_harts_0_trap_fsm_enumDef_RUNNING;
      end
      TrapPlugin_logic_harts_0_trap_fsm_enumDef_LSU_FLUSH : begin
        if(TrapPlugin_logic_lsuL1Invalidate_0_cmd_ready) begin
          TrapPlugin_logic_harts_0_trap_fsm_stateNext = TrapPlugin_logic_harts_0_trap_fsm_enumDef_FETCH_FLUSH;
        end
      end
      TrapPlugin_logic_harts_0_trap_fsm_enumDef_FETCH_FLUSH : begin
        if(TrapPlugin_logic_fetchL1Invalidate_0_cmd_ready) begin
          TrapPlugin_logic_harts_0_trap_fsm_stateNext = TrapPlugin_logic_harts_0_trap_fsm_enumDef_JUMP;
        end
      end
      default : begin
        if(when_TrapPlugin_l348) begin
          TrapPlugin_logic_harts_0_trap_fsm_stateNext = TrapPlugin_logic_harts_0_trap_fsm_enumDef_RUNNING;
        end
      end
    endcase
    if(TrapPlugin_logic_harts_0_trap_fsm_wantKill) begin
      TrapPlugin_logic_harts_0_trap_fsm_stateNext = TrapPlugin_logic_harts_0_trap_fsm_enumDef_RESET;
    end
  end

  assign when_TrapPlugin_l393 = ((TrapPlugin_logic_harts_0_trap_pending_state_exception || TrapPlugin_logic_harts_0_trap_fsm_triggerEbreak) || TrapPlugin_logic_harts_0_trap_fsm_buffer_trap_interrupt);
  always @(*) begin
    _zz_TrapPlugin_logic_harts_0_crsPorts_write_address = 3'b101;
    case(TrapPlugin_logic_harts_0_trap_fsm_buffer_trap_targetPrivilege)
      2'b01 : begin
        _zz_TrapPlugin_logic_harts_0_crsPorts_write_address = 3'b001;
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    _zz_TrapPlugin_logic_harts_0_crsPorts_write_address_1 = 3'b110;
    case(TrapPlugin_logic_harts_0_trap_fsm_buffer_trap_targetPrivilege)
      2'b01 : begin
        _zz_TrapPlugin_logic_harts_0_crsPorts_write_address_1 = 3'b010;
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    _zz_TrapPlugin_logic_harts_0_crsPorts_read_address = 3'b111;
    case(TrapPlugin_logic_harts_0_trap_fsm_buffer_trap_targetPrivilege)
      2'b01 : begin
        _zz_TrapPlugin_logic_harts_0_crsPorts_read_address = 3'b011;
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    _zz_TrapPlugin_logic_harts_0_crsPorts_read_address_1 = 3'b101;
    case(TrapPlugin_logic_harts_0_trap_fsm_xretPrivilege)
      2'b01 : begin
        _zz_TrapPlugin_logic_harts_0_crsPorts_read_address_1 = 3'b001;
      end
      default : begin
      end
    endcase
  end

  assign when_TrapPlugin_l637 = (TrapPlugin_logic_harts_0_trap_pending_xret_targetPrivilege != 2'b11);
  assign switch_TrapPlugin_l638 = TrapPlugin_logic_harts_0_trap_pending_state_arg[1 : 0];
  assign when_TrapPlugin_l492 = (TrapPlugin_logic_harts_0_trap_fsm_atsPorts_refill_rsp_payload_pageFault || TrapPlugin_logic_harts_0_trap_fsm_atsPorts_refill_rsp_payload_accessFault);
  assign switch_TrapPlugin_l494 = {TrapPlugin_logic_harts_0_trap_fsm_atsPorts_refill_rsp_payload_pageFault,TrapPlugin_logic_harts_0_trap_pending_state_arg[1 : 0]};
  assign when_TrapPlugin_l348 = (&{TrapPlugin_logic_harts_0_trap_fsm_atsPorts_invalidated,TrapPlugin_logic_harts_0_trap_fsm_resetToRunConditions_0});
  always @(*) begin
    MmuPlugin_logic_refill_stateNext = MmuPlugin_logic_refill_stateReg;
    case(MmuPlugin_logic_refill_stateReg)
      MmuPlugin_logic_refill_enumDef_IDLE : begin
        if(MmuPlugin_logic_refill_arbiter_io_output_valid) begin
          MmuPlugin_logic_refill_stateNext = MmuPlugin_logic_refill_enumDef_CMD_1;
        end
      end
      MmuPlugin_logic_refill_enumDef_CMD_0 : begin
        if(when_MmuPlugin_l454) begin
          if(MmuPlugin_logic_accessBus_cmd_ready) begin
            MmuPlugin_logic_refill_stateNext = MmuPlugin_logic_refill_enumDef_RSP_0;
          end
        end
      end
      MmuPlugin_logic_refill_enumDef_CMD_1 : begin
        if(when_MmuPlugin_l454_1) begin
          if(MmuPlugin_logic_accessBus_cmd_ready) begin
            MmuPlugin_logic_refill_stateNext = MmuPlugin_logic_refill_enumDef_RSP_1;
          end
        end
      end
      MmuPlugin_logic_refill_enumDef_RSP_0 : begin
        if(MmuPlugin_logic_refill_load_rsp_valid) begin
          if(MmuPlugin_logic_refill_load_rsp_payload_redo) begin
            MmuPlugin_logic_refill_stateNext = MmuPlugin_logic_refill_enumDef_CMD_0;
          end else begin
            MmuPlugin_logic_refill_stateNext = MmuPlugin_logic_refill_enumDef_IDLE;
          end
        end
      end
      MmuPlugin_logic_refill_enumDef_RSP_1 : begin
        if(MmuPlugin_logic_refill_load_rsp_valid) begin
          if(MmuPlugin_logic_refill_load_rsp_payload_redo) begin
            MmuPlugin_logic_refill_stateNext = MmuPlugin_logic_refill_enumDef_CMD_1;
          end else begin
            if(when_MmuPlugin_l471) begin
              MmuPlugin_logic_refill_stateNext = MmuPlugin_logic_refill_enumDef_IDLE;
            end else begin
              MmuPlugin_logic_refill_stateNext = MmuPlugin_logic_refill_enumDef_CMD_0;
            end
          end
        end
      end
      default : begin
      end
    endcase
    if(MmuPlugin_logic_refill_wantStart) begin
      MmuPlugin_logic_refill_stateNext = MmuPlugin_logic_refill_enumDef_IDLE;
    end
    if(MmuPlugin_logic_refill_wantKill) begin
      MmuPlugin_logic_refill_stateNext = MmuPlugin_logic_refill_enumDef_BOOT;
    end
  end

  assign when_MmuPlugin_l454 = (1'b1 && (MmuPlugin_logic_refill_cacheRefillAny == 1'b0));
  assign when_MmuPlugin_l454_1 = (1'b1 && (MmuPlugin_logic_refill_cacheRefillAny == 1'b0));
  assign when_MmuPlugin_l463 = (! MmuPlugin_logic_refill_load_leaf);
  assign when_MmuPlugin_l439 = (MmuPlugin_logic_refill_fetch_0_pageFault || MmuPlugin_logic_refill_fetch_0_accessFault);
  assign _zz_54 = MmuPlugin_logic_refill_portOhReg[0];
  assign when_MmuPlugin_l439_1 = (MmuPlugin_logic_refill_fetch_0_pageFault || MmuPlugin_logic_refill_fetch_0_accessFault);
  assign when_MmuPlugin_l471 = (MmuPlugin_logic_refill_load_leaf || MmuPlugin_logic_refill_load_exception);
  assign when_MmuPlugin_l439_2 = (MmuPlugin_logic_refill_fetch_1_pageFault || MmuPlugin_logic_refill_fetch_1_accessFault);
  assign when_MmuPlugin_l439_3 = (MmuPlugin_logic_refill_fetch_1_pageFault || MmuPlugin_logic_refill_fetch_1_accessFault);
  always @(*) begin
    CsrAccessPlugin_logic_fsm_stateNext = CsrAccessPlugin_logic_fsm_stateReg;
    case(CsrAccessPlugin_logic_fsm_stateReg)
      CsrAccessPlugin_logic_fsm_enumDef_READ : begin
        if(when_CsrAccessPlugin_l308) begin
          CsrAccessPlugin_logic_fsm_stateNext = CsrAccessPlugin_logic_fsm_enumDef_WRITE;
        end
      end
      CsrAccessPlugin_logic_fsm_enumDef_WRITE : begin
        if(when_CsrAccessPlugin_l338) begin
          CsrAccessPlugin_logic_fsm_stateNext = CsrAccessPlugin_logic_fsm_enumDef_COMPLETION;
        end
      end
      CsrAccessPlugin_logic_fsm_enumDef_COMPLETION : begin
        if(toplevel_execute_ctrl2_down_isReady) begin
          CsrAccessPlugin_logic_fsm_stateNext = CsrAccessPlugin_logic_fsm_enumDef_IDLE;
        end
      end
      default : begin
        if(CsrAccessPlugin_logic_fsm_inject_onDecodeDo) begin
          if(when_CsrAccessPlugin_l224) begin
            CsrAccessPlugin_logic_fsm_stateNext = CsrAccessPlugin_logic_fsm_enumDef_READ;
          end
          if(CsrAccessPlugin_logic_fsm_inject_sampled) begin
            if(!CsrAccessPlugin_logic_fsm_inject_trapReg) begin
              CsrAccessPlugin_logic_fsm_stateNext = CsrAccessPlugin_logic_fsm_enumDef_READ;
            end
          end
        end
      end
    endcase
    if(CsrAccessPlugin_logic_fsm_wantKill) begin
      CsrAccessPlugin_logic_fsm_stateNext = CsrAccessPlugin_logic_fsm_enumDef_IDLE;
    end
  end

  assign when_CsrAccessPlugin_l308 = (! CsrAccessPlugin_bus_read_halt);
  assign when_CsrAccessPlugin_l338 = (! CsrAccessPlugin_bus_write_halt);
  assign when_CsrAccessPlugin_l224 = ((! CsrAccessPlugin_logic_fsm_inject_trap) && (! CsrAccessPlugin_bus_decode_trap));
  always @(posedge clk_cpu or posedge reset_cpu) begin
    if(reset_cpu) begin
      MmuPlugin_logic_satp_mode <= 1'b0;
      MmuPlugin_logic_satp_ppn <= 20'h0;
      MmuPlugin_logic_status_mxr <= 1'b0;
      MmuPlugin_logic_status_sum <= 1'b0;
      MmuPlugin_logic_status_mprv <= 1'b0;
      early0_MulPlugin_logic_writeback_buffer_valid <= 1'b0;
      early0_DivPlugin_logic_processing_cmdSent <= 1'b0;
      early0_DivPlugin_logic_processing_relaxer_hadRequest <= 1'b0;
      early0_DivPlugin_logic_processing_unscheduleRequest <= 1'b0;
      AlignerPlugin_logic_feeder_harts_0_dopId <= 10'h0;
      AlignerPlugin_logic_buffer_mask <= 4'b0000;
      AlignerPlugin_logic_buffer_last <= 4'b0000;
      AlignerPlugin_logic_buffer_trap <= 1'b0;
      FetchL1Plugin_logic_invalidate_counter <= 7'h0;
      FetchL1Plugin_logic_invalidate_firstEver <= 1'b1;
      FetchL1Plugin_logic_refill_slots_0_valid <= 1'b0;
      FetchL1Plugin_logic_refill_slots_0_cmdSent <= 1'b1;
      FetchL1Plugin_logic_refill_pushCounter <= 32'h0;
      FetchL1Plugin_logic_refill_onRsp_wordIndex <= 3'b000;
      FetchL1Plugin_logic_refill_onRsp_firstCycle <= 1'b1;
      FetchL1Plugin_logic_ctrl_plruLogic_buffer_regNext_valid <= 1'b0;
      FetchL1Plugin_logic_ctrl_trapSent <= 1'b0;
      FetchL1Plugin_logic_ctrl_firstCycle <= 1'b1;
      FetchL1Plugin_logic_initializer_counter <= 10'h0;
      PrivilegedPlugin_logic_harts_0_privilege <= 2'b11;
      PrivilegedPlugin_logic_harts_0_m_status_mie <= 1'b0;
      PrivilegedPlugin_logic_harts_0_m_status_mpie <= 1'b0;
      PrivilegedPlugin_logic_harts_0_m_status_mpp <= 2'b00;
      PrivilegedPlugin_logic_harts_0_m_status_fs <= 2'b00;
      PrivilegedPlugin_logic_harts_0_m_status_tsr <= 1'b0;
      PrivilegedPlugin_logic_harts_0_m_status_tvm <= 1'b0;
      PrivilegedPlugin_logic_harts_0_m_status_tw <= 1'b0;
      PrivilegedPlugin_logic_harts_0_m_cause_interrupt <= 1'b0;
      PrivilegedPlugin_logic_harts_0_m_cause_code <= 4'b0000;
      PrivilegedPlugin_logic_harts_0_m_ip_meip <= 1'b0;
      PrivilegedPlugin_logic_harts_0_m_ip_mtip <= 1'b0;
      PrivilegedPlugin_logic_harts_0_m_ip_msip <= 1'b0;
      PrivilegedPlugin_logic_harts_0_m_ie_meie <= 1'b0;
      PrivilegedPlugin_logic_harts_0_m_ie_mtie <= 1'b0;
      PrivilegedPlugin_logic_harts_0_m_ie_msie <= 1'b0;
      PrivilegedPlugin_logic_harts_0_m_edeleg_iam <= 1'b0;
      PrivilegedPlugin_logic_harts_0_m_edeleg_bp <= 1'b0;
      PrivilegedPlugin_logic_harts_0_m_edeleg_eu <= 1'b0;
      PrivilegedPlugin_logic_harts_0_m_edeleg_es <= 1'b0;
      PrivilegedPlugin_logic_harts_0_m_edeleg_ipf <= 1'b0;
      PrivilegedPlugin_logic_harts_0_m_edeleg_lpf <= 1'b0;
      PrivilegedPlugin_logic_harts_0_m_edeleg_spf <= 1'b0;
      PrivilegedPlugin_logic_harts_0_m_ideleg_st <= 1'b0;
      PrivilegedPlugin_logic_harts_0_m_ideleg_se <= 1'b0;
      PrivilegedPlugin_logic_harts_0_m_ideleg_ss <= 1'b0;
      PrivilegedPlugin_logic_harts_0_s_cause_interrupt <= 1'b0;
      PrivilegedPlugin_logic_harts_0_s_cause_code <= 4'b0000;
      PrivilegedPlugin_logic_harts_0_s_status_sie <= 1'b0;
      PrivilegedPlugin_logic_harts_0_s_status_spie <= 1'b0;
      PrivilegedPlugin_logic_harts_0_s_status_spp <= 1'b0;
      PrivilegedPlugin_logic_harts_0_s_ip_seipSoft <= 1'b0;
      PrivilegedPlugin_logic_harts_0_s_ip_stip <= 1'b0;
      PrivilegedPlugin_logic_harts_0_s_ip_ssip <= 1'b0;
      PrivilegedPlugin_logic_harts_0_s_ie_seie <= 1'b0;
      PrivilegedPlugin_logic_harts_0_s_ie_stie <= 1'b0;
      PrivilegedPlugin_logic_harts_0_s_ie_ssie <= 1'b0;
      BtbPlugin_logic_ras_ptr_push <= 2'b00;
      BtbPlugin_logic_ras_ptr_pop <= 2'b11;
      toplevel_decode_ctrls_0_up_LANE_SEL_0_regNext <= 1'b0;
      toplevel_decode_ctrls_0_up_LANE_SEL_1_regNext <= 1'b0;
      late0_BranchPlugin_logic_jumpLogic_learn_rValid <= 1'b0;
      late1_BranchPlugin_logic_jumpLogic_learn_rValid <= 1'b0;
      GSharePlugin_logic_initializer_counter <= 13'h0;
      DecoderPlugin_logic_harts_0_uopId <= 16'h0;
      DecoderPlugin_logic_interrupt_buffered <= 1'b0;
      toplevel_decode_ctrls_1_up_LANE_SEL_0_regNext <= 1'b0;
      toplevel_decode_ctrls_1_up_LANE_SEL_1_regNext <= 1'b0;
      CsrRamPlugin_csrMapper_fired <= 1'b0;
      DispatchPlugin_logic_slots_0_ctx_valid <= 1'b0;
      DispatchPlugin_logic_feeds_0_sent <= 1'b0;
      DispatchPlugin_logic_feeds_1_sent <= 1'b0;
      toplevel_decode_ctrls_1_up_LANE_SEL_0_regNext_1 <= 1'b0;
      toplevel_decode_ctrls_1_up_LANE_SEL_1_regNext_1 <= 1'b0;
      toplevel_execute_ctrl0_down_LANE_SEL_lane0_regNext <= 1'b0;
      toplevel_execute_ctrl0_down_LANE_SEL_lane1_regNext <= 1'b0;
      toplevel_execute_ctrl2_down_LANE_SEL_lane0_regNext <= 1'b0;
      toplevel_execute_ctrl2_down_LANE_SEL_lane1_regNext <= 1'b0;
      BtbPlugin_logic_applyIt_correctionSent <= 1'b0;
      BtbPlugin_logic_initializer_counter <= 9'h0;
      toplevel_decode_ctrls_1_up_LANE_SEL_0 <= 1'b0;
      toplevel_decode_ctrls_1_up_LANE_SEL_1 <= 1'b0;
      LsuL1Plugin_logic_refill_slots_0_valid <= 1'b0;
      LsuL1Plugin_logic_refill_slots_0_loaded <= 1'b1;
      LsuL1Plugin_logic_refill_pushCounter <= 32'h0;
      LsuL1Plugin_logic_refill_read_arbiter_lock <= 1'b0;
      LsuL1Plugin_logic_refill_read_wordIndex <= 3'b000;
      LsuL1Plugin_logic_refill_read_hadError <= 1'b0;
      LsuL1Plugin_logic_writeback_slots_0_valid <= 1'b0;
      LsuL1Plugin_logic_writeback_slots_0_busy <= 1'b0;
      LsuL1Plugin_logic_writeback_read_arbiter_lock <= 1'b0;
      LsuL1Plugin_logic_writeback_read_wordIndex <= 3'b000;
      LsuL1Plugin_logic_writeback_read_slotReadLast_valid <= 1'b0;
      LsuL1Plugin_logic_writeback_write_arbiter_lock <= 1'b0;
      LsuL1Plugin_logic_writeback_write_wordIndex <= 3'b000;
      LsuL1Plugin_logic_writeback_write_bufferRead_rValid <= 1'b0;
      LsuL1Plugin_logic_ls_rb1_onBanks_0_busyReg <= 1'b0;
      LsuL1Plugin_logic_ls_rb1_onBanks_1_busyReg <= 1'b0;
      LsuL1Plugin_logic_ls_ctrl_hazardReg <= 1'b0;
      LsuL1Plugin_logic_ls_ctrl_flushHazardReg <= 1'b0;
      LsuL1Plugin_logic_initializer_counter <= 7'h0;
      LsuL1Plugin_logic_initializerMem_counter <= 10'h0;
      LsuPlugin_logic_onAddress0_ls_storeId <= 12'h0;
      LsuPlugin_logic_onAddress0_access_waiter_valid <= 1'b0;
      toplevel_execute_ctrl3_up_LsuL1_SEL_lane0 <= 1'b0;
      toplevel_execute_ctrl4_up_LsuL1_SEL_lane0 <= 1'b0;
      LsuPlugin_logic_onCtrl_io_tooEarly <= 1'b0;
      LsuPlugin_logic_onCtrl_io_allowIt <= 1'b0;
      LsuPlugin_logic_onCtrl_io_doItReg <= 1'b0;
      LsuPlugin_logic_onCtrl_io_cmdSent <= 1'b0;
      LsuPlugin_logic_bus_rsp_toStream_rValid <= 1'b0;
      LsuPlugin_logic_onCtrl_rva_nc_reserved <= 1'b0;
      LsuPlugin_logic_onCtrl_hartRegulation_valid <= 1'b0;
      LsuL1Plugin_logic_bus_toTilelink_nonCoherent_onA_lock <= 1'b0;
      LsuL1Plugin_logic_bus_toTilelink_nonCoherent_onA_beat <= 3'b000;
      TrapPlugin_logic_harts_0_interrupt_validBuffer <= 1'b0;
      TrapPlugin_logic_harts_0_trap_fsm_atsPorts_invalidated <= 1'b0;
      TrapPlugin_logic_harts_0_trap_fsm_trapEnterDebug <= 1'b0;
      FetchL1Plugin_logic_translationStorage_logic_sl_0_allocId_value <= 1'b0;
      LsuPlugin_logic_translationStorage_logic_sl_0_allocId_value <= 1'b0;
      MmuPlugin_logic_refill_cacheRefillAny <= 1'b0;
      MmuPlugin_logic_refill_load_rsp_valid <= 1'b0;
      MmuPlugin_logic_invalidate_busy <= 1'b0;
      LsuTileLinkPlugin_logic_bridge_pendings_0_valid <= 1'b0;
      PcPlugin_logic_harts_0_self_id <= 10'h0;
      PcPlugin_logic_harts_0_self_increment <= 1'b0;
      PcPlugin_logic_harts_0_self_fault <= 1'b0;
      PcPlugin_logic_harts_0_self_state <= 32'h40000000;
      PcPlugin_logic_harts_0_holdReg <= 1'b1;
      CsrAccessPlugin_logic_fsm_inject_unfreeze <= 1'b0;
      CsrAccessPlugin_logic_fsm_inject_flushReg <= 1'b0;
      CsrAccessPlugin_logic_fsm_inject_sampled <= 1'b0;
      HistoryPlugin_logic_onFetch_value <= 12'h0;
      CsrRamPlugin_logic_readLogic_ohReg <= 2'b00;
      CsrRamPlugin_logic_readLogic_busy <= 1'b0;
      CsrRamPlugin_logic_flush_counter <= 4'b0000;
      toplevel_execute_ctrl1_up_LANE_SEL_lane0 <= 1'b0;
      toplevel_execute_ctrl2_up_LANE_SEL_lane0 <= 1'b0;
      toplevel_execute_ctrl3_up_LANE_SEL_lane0 <= 1'b0;
      toplevel_execute_ctrl4_up_LANE_SEL_lane0 <= 1'b0;
      toplevel_execute_ctrl5_up_LANE_SEL_lane0 <= 1'b0;
      toplevel_execute_ctrl1_up_LANE_SEL_lane1 <= 1'b0;
      toplevel_execute_ctrl2_up_LANE_SEL_lane1 <= 1'b0;
      toplevel_execute_ctrl3_up_LANE_SEL_lane1 <= 1'b0;
      toplevel_execute_ctrl4_up_LANE_SEL_lane1 <= 1'b0;
      toplevel_execute_ctrl5_up_LANE_SEL_lane1 <= 1'b0;
      integer_RegFilePlugin_logic_initalizer_counter <= 6'h0;
      _zz_WhiteboxerPlugin_logic_perf_executeFreezedCounter_2 <= 60'h0;
      _zz_WhiteboxerPlugin_logic_perf_dispatchHazardsCounter_2 <= 60'h0;
      _zz_WhiteboxerPlugin_logic_perf_candidatesCountCounters_0_2 <= 60'h0;
      _zz_WhiteboxerPlugin_logic_perf_candidatesCountCounters_1_2 <= 60'h0;
      _zz_WhiteboxerPlugin_logic_perf_candidatesCountCounters_2_2 <= 60'h0;
      _zz_WhiteboxerPlugin_logic_perf_candidatesCountCounters_3_2 <= 60'h0;
      _zz_WhiteboxerPlugin_logic_perf_dispatchFeedCounters_0_2 <= 60'h0;
      _zz_WhiteboxerPlugin_logic_perf_dispatchFeedCounters_1_2 <= 60'h0;
      _zz_WhiteboxerPlugin_logic_perf_dispatchFeedCounters_2_2 <= 60'h0;
      fetch_logic_ctrls_1_up_valid <= 1'b0;
      fetch_logic_ctrls_2_up_valid <= 1'b0;
      toplevel_decode_ctrls_1_up_valid <= 1'b0;
      LsuPlugin_logic_flusher_stateReg <= LsuPlugin_logic_flusher_enumDef_IDLE;
      TrapPlugin_logic_harts_0_trap_fsm_stateReg <= TrapPlugin_logic_harts_0_trap_fsm_enumDef_RESET;
      MmuPlugin_logic_refill_stateReg <= MmuPlugin_logic_refill_enumDef_BOOT;
      CsrAccessPlugin_logic_fsm_stateReg <= CsrAccessPlugin_logic_fsm_enumDef_IDLE;
    end else begin
      early0_MulPlugin_logic_writeback_buffer_valid <= 1'b0;
      if(when_MulPlugin_l195) begin
        early0_MulPlugin_logic_writeback_buffer_valid <= 1'b1;
      end
      if(early0_DivPlugin_logic_processing_div_io_cmd_fire) begin
        early0_DivPlugin_logic_processing_cmdSent <= 1'b1;
      end
      if(toplevel_execute_ctrl2_down_isReady) begin
        early0_DivPlugin_logic_processing_cmdSent <= 1'b0;
      end
      early0_DivPlugin_logic_processing_relaxer_hadRequest <= (early0_DivPlugin_logic_processing_request && execute_freeze_valid);
      early0_DivPlugin_logic_processing_unscheduleRequest <= toplevel_execute_lane0_ctrls_2_upIsCancel;
      if(toplevel_execute_ctrl2_down_isReady) begin
        early0_DivPlugin_logic_processing_unscheduleRequest <= 1'b0;
      end
      if(when_AlignerPlugin_l173) begin
        AlignerPlugin_logic_feeder_harts_0_dopId <= (toplevel_decode_ctrls_0_down_Decode_DOP_ID_1 + 10'h001);
      end
      if(AlignerPlugin_logic_buffer_downFire) begin
        AlignerPlugin_logic_buffer_mask <= (AlignerPlugin_logic_buffer_mask & (~ AlignerPlugin_logic_buffer_usedMask[3 : 0]));
        AlignerPlugin_logic_buffer_last <= (AlignerPlugin_logic_buffer_last & (~ AlignerPlugin_logic_buffer_usedMask[3 : 0]));
      end
      if(when_AlignerPlugin_l259) begin
        AlignerPlugin_logic_buffer_mask <= (fetch_logic_ctrls_2_down_AlignerPlugin_logic_FETCH_MASK & (~ (AlignerPlugin_logic_buffer_downFire ? AlignerPlugin_logic_buffer_usedMask[7 : 4] : 4'b0000)));
        AlignerPlugin_logic_buffer_trap <= fetch_logic_ctrls_2_down_TRAP;
        AlignerPlugin_logic_buffer_last <= fetch_logic_ctrls_2_down_AlignerPlugin_logic_FETCH_LAST;
      end
      if(FetchL1Plugin_logic_invalidate_done) begin
        FetchL1Plugin_logic_invalidate_firstEver <= 1'b0;
      end
      if(when_FetchL1Plugin_l220) begin
        FetchL1Plugin_logic_invalidate_counter <= FetchL1Plugin_logic_invalidate_counterIncr;
      end
      if(when_FetchL1Plugin_l227) begin
        FetchL1Plugin_logic_invalidate_counter <= 7'h0;
      end
      if(when_FetchL1Plugin_l271) begin
        if(_zz_when) begin
          FetchL1Plugin_logic_refill_slots_0_valid <= 1'b1;
          FetchL1Plugin_logic_refill_slots_0_cmdSent <= 1'b0;
        end
        FetchL1Plugin_logic_refill_pushCounter <= (FetchL1Plugin_logic_refill_pushCounter + 32'h00000001);
      end
      if(FetchL1Plugin_logic_bus_cmd_ready) begin
        if(FetchL1Plugin_logic_refill_onCmd_oh[0]) begin
          FetchL1Plugin_logic_refill_slots_0_cmdSent <= 1'b1;
        end
      end
      if(FetchL1Plugin_logic_bus_rsp_fire) begin
        FetchL1Plugin_logic_refill_onRsp_firstCycle <= 1'b0;
      end
      if(FetchL1Plugin_logic_bus_rsp_valid) begin
        FetchL1Plugin_logic_refill_onRsp_wordIndex <= (FetchL1Plugin_logic_refill_onRsp_wordIndex + 3'b001);
        if(when_FetchL1Plugin_l350) begin
          FetchL1Plugin_logic_refill_onRsp_firstCycle <= 1'b1;
          FetchL1Plugin_logic_refill_slots_0_valid <= 1'b0;
        end
      end
      FetchL1Plugin_logic_ctrl_plruLogic_buffer_regNext_valid <= FetchL1Plugin_logic_ctrl_plruLogic_buffer_valid;
      if(FetchL1Plugin_logic_trapPort_valid) begin
        FetchL1Plugin_logic_ctrl_trapSent <= 1'b1;
      end
      if(fetch_logic_ctrls_2_up_isCancel) begin
        FetchL1Plugin_logic_ctrl_trapSent <= 1'b0;
      end
      if(fetch_logic_ctrls_2_up_isValid) begin
        FetchL1Plugin_logic_ctrl_firstCycle <= 1'b0;
      end
      if(when_FetchL1Plugin_l550) begin
        FetchL1Plugin_logic_ctrl_firstCycle <= 1'b1;
      end
      `ifndef SYNTHESIS
        `ifdef FORMAL
          assert((! ((|FetchL1Plugin_logic_refill_slots_0_valid) && (! FetchL1Plugin_logic_invalidate_done)))); // FetchL1Plugin.scala:L565
        `else
          if(!(! ((|FetchL1Plugin_logic_refill_slots_0_valid) && (! FetchL1Plugin_logic_invalidate_done)))) begin
            $display("FAILURE "); // FetchL1Plugin.scala:L565
            $finish;
          end
        `endif
      `endif
      if(FetchL1Plugin_logic_initializer_busy) begin
        FetchL1Plugin_logic_initializer_counter <= (FetchL1Plugin_logic_initializer_counter + 10'h001);
      end
      PrivilegedPlugin_logic_harts_0_m_ip_meip <= PrivilegedPlugin_logic_harts_0_int_m_external;
      PrivilegedPlugin_logic_harts_0_m_ip_mtip <= PrivilegedPlugin_logic_harts_0_int_m_timer;
      PrivilegedPlugin_logic_harts_0_m_ip_msip <= PrivilegedPlugin_logic_harts_0_int_m_software;
      BtbPlugin_logic_ras_ptr_push <= (_zz_BtbPlugin_logic_ras_ptr_push - _zz_BtbPlugin_logic_ras_ptr_push_3);
      toplevel_decode_ctrls_0_up_LANE_SEL_0_regNext <= toplevel_decode_ctrls_0_up_LANE_SEL_0;
      if(when_CtrlLaneApi_l46) begin
        toplevel_decode_ctrls_0_up_LANE_SEL_0_regNext <= 1'b0;
      end
      toplevel_decode_ctrls_0_up_LANE_SEL_1_regNext <= toplevel_decode_ctrls_0_up_LANE_SEL_1;
      if(when_CtrlLaneApi_l46_1) begin
        toplevel_decode_ctrls_0_up_LANE_SEL_1_regNext <= 1'b0;
      end
      if(PrivilegedPlugin_logic_harts_0_xretAwayFromMachine) begin
        MmuPlugin_logic_status_mprv <= 1'b0;
      end
      if(late0_BranchPlugin_logic_jumpLogic_learn_ready) begin
        late0_BranchPlugin_logic_jumpLogic_learn_rValid <= late0_BranchPlugin_logic_jumpLogic_learn_valid;
      end
      if(late1_BranchPlugin_logic_jumpLogic_learn_ready) begin
        late1_BranchPlugin_logic_jumpLogic_learn_rValid <= late1_BranchPlugin_logic_jumpLogic_learn_valid;
      end
      if(GSharePlugin_logic_initializer_busy) begin
        GSharePlugin_logic_initializer_counter <= (GSharePlugin_logic_initializer_counter + 13'h0001);
      end
      if(when_DecoderPlugin_l135) begin
        DecoderPlugin_logic_harts_0_uopId <= (DecoderPlugin_logic_harts_0_uopId + 16'h0002);
      end
      if(when_DecoderPlugin_l143) begin
        DecoderPlugin_logic_interrupt_buffered <= DecoderPlugin_logic_interrupt_async;
      end
      toplevel_decode_ctrls_1_up_LANE_SEL_0_regNext <= toplevel_decode_ctrls_1_up_LANE_SEL_0;
      if(when_CtrlLaneApi_l46_2) begin
        toplevel_decode_ctrls_1_up_LANE_SEL_0_regNext <= 1'b0;
      end
      toplevel_decode_ctrls_1_up_LANE_SEL_1_regNext <= toplevel_decode_ctrls_1_up_LANE_SEL_1;
      if(when_CtrlLaneApi_l46_3) begin
        toplevel_decode_ctrls_1_up_LANE_SEL_1_regNext <= 1'b0;
      end
      if(when_CsrRamPlugin_l84) begin
        CsrRamPlugin_csrMapper_fired <= 1'b1;
      end
      if(CsrAccessPlugin_bus_write_moving) begin
        CsrRamPlugin_csrMapper_fired <= 1'b0;
      end
      if(DispatchPlugin_logic_feeds_0_sending) begin
        DispatchPlugin_logic_feeds_0_sent <= 1'b1;
      end
      if(toplevel_decode_ctrls_1_up_isMoving) begin
        DispatchPlugin_logic_feeds_0_sent <= 1'b0;
      end
      if(DispatchPlugin_logic_feeds_1_sending) begin
        DispatchPlugin_logic_feeds_1_sent <= 1'b1;
      end
      if(toplevel_decode_ctrls_1_up_isMoving) begin
        DispatchPlugin_logic_feeds_1_sent <= 1'b0;
      end
      if(when_DispatchPlugin_l368) begin
        DispatchPlugin_logic_slots_0_ctx_valid <= 1'b0;
      end
      toplevel_decode_ctrls_1_up_LANE_SEL_0_regNext_1 <= toplevel_decode_ctrls_1_up_LANE_SEL_0;
      if(when_CtrlLaneApi_l46_4) begin
        toplevel_decode_ctrls_1_up_LANE_SEL_0_regNext_1 <= 1'b0;
      end
      toplevel_decode_ctrls_1_up_LANE_SEL_1_regNext_1 <= toplevel_decode_ctrls_1_up_LANE_SEL_1;
      if(when_CtrlLaneApi_l46_5) begin
        toplevel_decode_ctrls_1_up_LANE_SEL_1_regNext_1 <= 1'b0;
      end
      toplevel_execute_ctrl0_down_LANE_SEL_lane0_regNext <= toplevel_execute_ctrl0_down_LANE_SEL_lane0;
      if(when_CtrlLaneApi_l46_6) begin
        toplevel_execute_ctrl0_down_LANE_SEL_lane0_regNext <= 1'b0;
      end
      toplevel_execute_ctrl0_down_LANE_SEL_lane1_regNext <= toplevel_execute_ctrl0_down_LANE_SEL_lane1;
      if(when_CtrlLaneApi_l46_7) begin
        toplevel_execute_ctrl0_down_LANE_SEL_lane1_regNext <= 1'b0;
      end
      toplevel_execute_ctrl2_down_LANE_SEL_lane0_regNext <= toplevel_execute_ctrl2_down_LANE_SEL_lane0;
      if(when_CtrlLaneApi_l46_8) begin
        toplevel_execute_ctrl2_down_LANE_SEL_lane0_regNext <= 1'b0;
      end
      toplevel_execute_ctrl2_down_LANE_SEL_lane1_regNext <= toplevel_execute_ctrl2_down_LANE_SEL_lane1;
      if(when_CtrlLaneApi_l46_9) begin
        toplevel_execute_ctrl2_down_LANE_SEL_lane1_regNext <= 1'b0;
      end
      `ifndef SYNTHESIS
        `ifdef FORMAL
          assert((! (fetch_logic_ctrls_1_up_isValid && fetch_logic_ctrls_1_down_BtbPlugin_logic_readCmd_HAZARDS[0]))); // BtbPlugin.scala:L187
        `else
          if(!(! (fetch_logic_ctrls_1_up_isValid && fetch_logic_ctrls_1_down_BtbPlugin_logic_readCmd_HAZARDS[0]))) begin
            $display("FAILURE "); // BtbPlugin.scala:L187
            $finish;
          end
        `endif
      `endif
      `ifndef SYNTHESIS
        `ifdef FORMAL
          assert((! (fetch_logic_ctrls_1_up_isValid && fetch_logic_ctrls_1_down_BtbPlugin_logic_readCmd_HAZARDS[1]))); // BtbPlugin.scala:L187
        `else
          if(!(! (fetch_logic_ctrls_1_up_isValid && fetch_logic_ctrls_1_down_BtbPlugin_logic_readCmd_HAZARDS[1]))) begin
            $display("FAILURE "); // BtbPlugin.scala:L187
            $finish;
          end
        `endif
      `endif
      if(fetch_logic_ctrls_2_up_isValid) begin
        BtbPlugin_logic_applyIt_correctionSent <= 1'b1;
      end
      if(when_BtbPlugin_l205) begin
        BtbPlugin_logic_applyIt_correctionSent <= 1'b0;
      end
      if(BtbPlugin_logic_initializer_busy) begin
        BtbPlugin_logic_initializer_counter <= (BtbPlugin_logic_initializer_counter + 9'h001);
      end
      if(AlignerPlugin_logic_buffer_flushIt) begin
        AlignerPlugin_logic_buffer_mask <= 4'b0000;
        AlignerPlugin_logic_buffer_last <= 4'b0000;
      end
      if(DispatchPlugin_logic_slotsFeeds_doIt) begin
        DispatchPlugin_logic_slots_0_ctx_valid <= _zz_DispatchPlugin_logic_slots_0_ctx_valid_4[0];
      end
      if(LsuL1Plugin_logic_refill_slots_0_loadedSet) begin
        LsuL1Plugin_logic_refill_slots_0_loaded <= 1'b1;
      end
      if(LsuL1Plugin_logic_refill_slots_0_fire) begin
        LsuL1Plugin_logic_refill_slots_0_valid <= 1'b0;
      end
      if(LsuL1Plugin_logic_refill_push_valid) begin
        LsuL1Plugin_logic_refill_pushCounter <= (LsuL1Plugin_logic_refill_pushCounter + 32'h00000001);
      end
      if(LsuL1Plugin_logic_refill_push_valid) begin
        if(when_LsuL1Plugin_l358) begin
          LsuL1Plugin_logic_refill_slots_0_valid <= 1'b1;
          LsuL1Plugin_logic_refill_slots_0_loaded <= 1'b0;
        end
      end
      LsuL1Plugin_logic_refill_read_arbiter_lock <= LsuL1Plugin_logic_refill_read_arbiter_oh;
      if(LsuL1Plugin_logic_bus_read_cmd_fire) begin
        LsuL1Plugin_logic_refill_read_arbiter_lock <= 1'b0;
      end
      if(LsuL1Plugin_logic_bus_read_rsp_valid) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(LsuL1Plugin_logic_refill_read_writeReservation_win); // LsuL1Plugin.scala:L408
          `else
            if(!LsuL1Plugin_logic_refill_read_writeReservation_win) begin
              $display("FAILURE "); // LsuL1Plugin.scala:L408
              $finish;
            end
          `endif
        `endif
      end
      if(when_LsuL1Plugin_l434) begin
        LsuL1Plugin_logic_refill_read_hadError <= 1'b1;
      end
      if(LsuL1Plugin_logic_bus_read_rsp_valid) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(LsuL1Plugin_logic_refill_read_reservation_win); // LsuL1Plugin.scala:L442
          `else
            if(!LsuL1Plugin_logic_refill_read_reservation_win) begin
              $display("FAILURE "); // LsuL1Plugin.scala:L442
              $finish;
            end
          `endif
        `endif
        if(LsuL1Plugin_logic_refill_read_rspWithData) begin
          LsuL1Plugin_logic_refill_read_wordIndex <= (LsuL1Plugin_logic_refill_read_wordIndex + 3'b001);
        end
        if(when_LsuL1Plugin_l446) begin
          LsuL1Plugin_logic_refill_read_hadError <= 1'b0;
        end
      end
      if(LsuL1Plugin_logic_writeback_slots_0_fire) begin
        LsuL1Plugin_logic_writeback_slots_0_valid <= 1'b0;
      end
      if(LsuL1Plugin_logic_writeback_slots_0_fire) begin
        LsuL1Plugin_logic_writeback_slots_0_busy <= 1'b0;
      end
      if(when_LsuL1Plugin_l509) begin
        LsuL1Plugin_logic_writeback_slots_0_valid <= 1'b0;
      end
      if(LsuL1Plugin_logic_writeback_push_valid) begin
        if(when_LsuL1Plugin_l532) begin
          LsuL1Plugin_logic_writeback_slots_0_valid <= 1'b1;
          LsuL1Plugin_logic_writeback_slots_0_busy <= 1'b1;
        end
      end
      LsuL1Plugin_logic_writeback_read_arbiter_lock <= LsuL1Plugin_logic_writeback_read_arbiter_oh;
      LsuL1Plugin_logic_writeback_read_wordIndex <= (LsuL1Plugin_logic_writeback_read_wordIndex + _zz_LsuL1Plugin_logic_writeback_read_wordIndex);
      if(when_LsuL1Plugin_l577) begin
        LsuL1Plugin_logic_writeback_read_arbiter_lock <= 1'b0;
      end
      LsuL1Plugin_logic_writeback_read_slotReadLast_valid <= LsuL1Plugin_logic_writeback_read_slotRead_valid;
      LsuL1Plugin_logic_writeback_write_arbiter_lock <= LsuL1Plugin_logic_writeback_write_arbiter_oh;
      LsuL1Plugin_logic_writeback_write_wordIndex <= (LsuL1Plugin_logic_writeback_write_wordIndex + _zz_LsuL1Plugin_logic_writeback_write_wordIndex);
      if(when_LsuL1Plugin_l651) begin
        LsuL1Plugin_logic_writeback_write_arbiter_lock <= 1'b0;
      end
      if(LsuL1Plugin_logic_writeback_write_bufferRead_ready) begin
        LsuL1Plugin_logic_writeback_write_bufferRead_rValid <= LsuL1Plugin_logic_writeback_write_bufferRead_valid;
      end
      if(LsuL1Plugin_logic_banks_0_usedByWriteback) begin
        LsuL1Plugin_logic_ls_rb1_onBanks_0_busyReg <= 1'b1;
      end
      if(when_LsuL1Plugin_l706) begin
        LsuL1Plugin_logic_ls_rb1_onBanks_0_busyReg <= 1'b0;
      end
      if(LsuL1Plugin_logic_banks_1_usedByWriteback) begin
        LsuL1Plugin_logic_ls_rb1_onBanks_1_busyReg <= 1'b1;
      end
      if(when_LsuL1Plugin_l706_1) begin
        LsuL1Plugin_logic_ls_rb1_onBanks_1_busyReg <= 1'b0;
      end
      LsuL1Plugin_logic_ls_ctrl_hazardReg <= (toplevel_execute_ctrl4_down_LsuL1_HAZARD_lane0 && execute_freeze_valid);
      LsuL1Plugin_logic_ls_ctrl_flushHazardReg <= (toplevel_execute_ctrl4_down_LsuL1_FLUSH_HAZARD_lane0 && execute_freeze_valid);
      if(toplevel_execute_ctrl4_down_LsuL1_SEL_lane0) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert((_zz_55 <= 2'b01)); // LsuL1Plugin.scala:L855
          `else
            if(!(_zz_55 <= 2'b01)) begin
              $display("FAILURE Multiple way hit ???"); // LsuL1Plugin.scala:L855
              $finish;
            end
          `endif
        `endif
      end
      if(when_LsuL1Plugin_l876) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert((_zz_57 < 2'b10)); // LsuL1Plugin.scala:L877
          `else
            if(!(_zz_57 < 2'b10)) begin
              $display("FAILURE "); // LsuL1Plugin.scala:L877
              $finish;
            end
          `endif
        `endif
      end
      if(when_LsuL1Plugin_l1160) begin
        LsuL1Plugin_logic_initializer_counter <= (LsuL1Plugin_logic_initializer_counter + 7'h01);
      end
      if(LsuL1Plugin_logic_initializerMem_busy) begin
        LsuL1Plugin_logic_initializerMem_counter <= (LsuL1Plugin_logic_initializerMem_counter + 10'h001);
      end
      LsuPlugin_logic_onAddress0_ls_storeId <= (LsuPlugin_logic_onAddress0_ls_storeId + _zz_LsuPlugin_logic_onAddress0_ls_storeId);
      if(when_LsuPlugin_l200) begin
        LsuPlugin_logic_onAddress0_access_waiter_valid <= 1'b0;
      end
      LsuPlugin_logic_onCtrl_io_tooEarly <= 1'b1;
      if(execute_freeze_valid) begin
        LsuPlugin_logic_onCtrl_io_tooEarly <= 1'b0;
      end
      LsuPlugin_logic_onCtrl_io_allowIt <= 1'b0;
      if(when_LsuPlugin_l491) begin
        LsuPlugin_logic_onCtrl_io_allowIt <= 1'b1;
      end
      LsuPlugin_logic_onCtrl_io_doItReg <= LsuPlugin_logic_onCtrl_io_doIt;
      if(LsuPlugin_logic_bus_cmd_fire) begin
        LsuPlugin_logic_onCtrl_io_cmdSent <= 1'b1;
      end
      if(when_LsuPlugin_l495) begin
        LsuPlugin_logic_onCtrl_io_cmdSent <= 1'b0;
      end
      if(LsuPlugin_logic_bus_rsp_toStream_valid) begin
        LsuPlugin_logic_bus_rsp_toStream_rValid <= 1'b1;
      end
      if(LsuPlugin_logic_onCtrl_io_rsp_fire) begin
        LsuPlugin_logic_bus_rsp_toStream_rValid <= 1'b0;
      end
      if(when_LsuPlugin_l573) begin
        if(toplevel_execute_ctrl4_down_LsuL1_STORE_lane0) begin
          LsuPlugin_logic_onCtrl_rva_nc_reserved <= 1'b0;
        end
      end
      if(when_LsuPlugin_l585) begin
        LsuPlugin_logic_onCtrl_rva_nc_reserved <= 1'b0;
      end
      if(LsuPlugin_logic_onCtrl_rva_nc_capture) begin
        LsuPlugin_logic_onCtrl_rva_nc_reserved <= (! LsuPlugin_logic_onCtrl_rva_nc_reserved);
      end
      if(when_LsuPlugin_l796) begin
        if(when_LsuPlugin_l204) begin
          LsuPlugin_logic_onAddress0_access_waiter_valid <= 1'b1;
        end
      end
      if(when_LsuPlugin_l200_1) begin
        LsuPlugin_logic_onCtrl_hartRegulation_valid <= 1'b0;
      end
      if(when_LsuPlugin_l803) begin
        if(when_LsuPlugin_l204_1) begin
          LsuPlugin_logic_onCtrl_hartRegulation_valid <= 1'b1;
        end
      end
      if(LsuL1TileLinkPlugin_logic_down_a_valid) begin
        LsuL1Plugin_logic_bus_toTilelink_nonCoherent_onA_lock <= 1'b1;
      end
      if(LsuL1TileLinkPlugin_logic_down_a_fire) begin
        LsuL1Plugin_logic_bus_toTilelink_nonCoherent_onA_beat <= (LsuL1Plugin_logic_bus_toTilelink_nonCoherent_onA_beat + 3'b001);
        if(LsuL1TileLinkPlugin_logic_down_a_tracker_last) begin
          LsuL1Plugin_logic_bus_toTilelink_nonCoherent_onA_beat <= 3'b000;
        end
      end
      if(when_LsuL1Bus_l402) begin
        LsuL1Plugin_logic_bus_toTilelink_nonCoherent_onA_lock <= 1'b0;
      end
      TrapPlugin_logic_harts_0_interrupt_validBuffer <= TrapPlugin_logic_harts_0_interrupt_valid;
      if(TrapPlugin_logic_harts_0_trap_fsm_atsPorts_invalidate_cmd_fire) begin
        TrapPlugin_logic_harts_0_trap_fsm_atsPorts_invalidated <= 1'b1;
      end
      FetchL1Plugin_logic_translationStorage_logic_sl_0_allocId_value <= FetchL1Plugin_logic_translationStorage_logic_sl_0_allocId_valueNext;
      LsuPlugin_logic_translationStorage_logic_sl_0_allocId_value <= LsuPlugin_logic_translationStorage_logic_sl_0_allocId_valueNext;
      MmuPlugin_logic_refill_cacheRefillAny <= ((MmuPlugin_logic_refill_cacheRefillAny || MmuPlugin_logic_refill_cacheRefillAnySet) && (! 1'b0));
      MmuPlugin_logic_refill_load_rsp_valid <= MmuPlugin_logic_accessBus_rsp_valid;
      if(when_MmuPlugin_l496) begin
        if(MmuPlugin_logic_invalidate_arbiter_io_output_valid) begin
          MmuPlugin_logic_invalidate_busy <= 1'b1;
        end
      end else begin
        if(when_MmuPlugin_l510) begin
          MmuPlugin_logic_invalidate_busy <= 1'b0;
        end
      end
      if(LsuTileLinkPlugin_logic_bridge_down_d_fire) begin
        LsuTileLinkPlugin_logic_bridge_pendings_0_valid <= 1'b0;
      end
      if(LsuTileLinkPlugin_logic_bridge_down_a_fire) begin
        LsuTileLinkPlugin_logic_bridge_pendings_0_valid <= 1'b1;
      end
      PcPlugin_logic_harts_0_holdReg <= PcPlugin_logic_harts_0_holdComb;
      PcPlugin_logic_harts_0_self_state <= PcPlugin_logic_harts_0_output_payload_pc;
      PcPlugin_logic_harts_0_self_fault <= PcPlugin_logic_harts_0_output_payload_fault;
      PcPlugin_logic_harts_0_self_increment <= 1'b0;
      if(PcPlugin_logic_harts_0_output_fire) begin
        PcPlugin_logic_harts_0_self_increment <= 1'b1;
        PcPlugin_logic_harts_0_self_state[2 : 1] <= 2'b00;
      end
      if(fetch_logic_ctrls_0_up_isFiring) begin
        PcPlugin_logic_harts_0_self_id <= (PcPlugin_logic_harts_0_self_id + 10'h001);
      end
      `ifndef SYNTHESIS
        `ifdef FORMAL
          assert((! ((toplevel_execute_ctrl2_up_LANE_SEL_lane0 && toplevel_execute_ctrl2_down_CsrAccessPlugin_SEL_lane0) && toplevel_execute_lane0_ctrls_2_upIsCancel))); // CsrAccessPlugin.scala:L136
        `else
          if(!(! ((toplevel_execute_ctrl2_up_LANE_SEL_lane0 && toplevel_execute_ctrl2_down_CsrAccessPlugin_SEL_lane0) && toplevel_execute_lane0_ctrls_2_upIsCancel))) begin
            $display("FAILURE CsrAccessPlugin saw forbidden select && cancel request"); // CsrAccessPlugin.scala:L136
            $finish;
          end
        `endif
      `endif
      CsrAccessPlugin_logic_fsm_inject_unfreeze <= 1'b0;
      if(CsrAccessPlugin_logic_flushPort_valid) begin
        CsrAccessPlugin_logic_fsm_inject_flushReg <= 1'b1;
      end
      if(when_CsrAccessPlugin_l209) begin
        CsrAccessPlugin_logic_fsm_inject_flushReg <= 1'b0;
      end
      CsrAccessPlugin_logic_fsm_inject_sampled <= execute_freeze_valid;
      if(when_CsrAccessPlugin_l359) begin
        PrivilegedPlugin_logic_harts_0_m_status_mpie <= CsrAccessPlugin_bus_write_bits[7];
        PrivilegedPlugin_logic_harts_0_m_status_mie <= CsrAccessPlugin_bus_write_bits[3];
        if(when_CsrService_l166) begin
          case(switch_PrivilegedPlugin_l540)
            2'b11 : begin
              PrivilegedPlugin_logic_harts_0_m_status_mpp <= 2'b11;
            end
            2'b01 : begin
              PrivilegedPlugin_logic_harts_0_m_status_mpp <= 2'b01;
            end
            2'b00 : begin
              PrivilegedPlugin_logic_harts_0_m_status_mpp <= 2'b00;
            end
            default : begin
            end
          endcase
        end
        PrivilegedPlugin_logic_harts_0_m_status_fs <= CsrAccessPlugin_bus_write_bits[14 : 13];
        PrivilegedPlugin_logic_harts_0_m_status_tsr <= CsrAccessPlugin_bus_write_bits[22];
        PrivilegedPlugin_logic_harts_0_m_status_tvm <= CsrAccessPlugin_bus_write_bits[20];
        PrivilegedPlugin_logic_harts_0_m_status_tw <= CsrAccessPlugin_bus_write_bits[21];
        PrivilegedPlugin_logic_harts_0_s_status_spp <= CsrAccessPlugin_bus_write_bits[8 : 8];
        PrivilegedPlugin_logic_harts_0_s_status_spie <= CsrAccessPlugin_bus_write_bits[5];
        PrivilegedPlugin_logic_harts_0_s_status_sie <= CsrAccessPlugin_bus_write_bits[1];
        MmuPlugin_logic_status_mxr <= CsrAccessPlugin_bus_write_bits[19];
        MmuPlugin_logic_status_sum <= CsrAccessPlugin_bus_write_bits[18];
        MmuPlugin_logic_status_mprv <= CsrAccessPlugin_bus_write_bits[17];
      end
      if(when_CsrAccessPlugin_l359_1) begin
        PrivilegedPlugin_logic_harts_0_m_cause_interrupt <= CsrAccessPlugin_bus_write_bits[31];
        PrivilegedPlugin_logic_harts_0_m_cause_code <= CsrAccessPlugin_bus_write_bits[3 : 0];
      end
      if(when_CsrAccessPlugin_l359_2) begin
        PrivilegedPlugin_logic_harts_0_s_ip_seipSoft <= CsrAccessPlugin_bus_write_bits[9];
        PrivilegedPlugin_logic_harts_0_s_ip_stip <= CsrAccessPlugin_bus_write_bits[5];
        PrivilegedPlugin_logic_harts_0_s_ip_ssip <= CsrAccessPlugin_bus_write_bits[1];
      end
      if(when_CsrAccessPlugin_l359_3) begin
        PrivilegedPlugin_logic_harts_0_m_ie_meie <= CsrAccessPlugin_bus_write_bits[11];
        PrivilegedPlugin_logic_harts_0_m_ie_mtie <= CsrAccessPlugin_bus_write_bits[7];
        PrivilegedPlugin_logic_harts_0_m_ie_msie <= CsrAccessPlugin_bus_write_bits[3];
        PrivilegedPlugin_logic_harts_0_s_ie_seie <= CsrAccessPlugin_bus_write_bits[9];
        PrivilegedPlugin_logic_harts_0_s_ie_stie <= CsrAccessPlugin_bus_write_bits[5];
        PrivilegedPlugin_logic_harts_0_s_ie_ssie <= CsrAccessPlugin_bus_write_bits[1];
      end
      if(when_CsrAccessPlugin_l359_4) begin
        PrivilegedPlugin_logic_harts_0_m_edeleg_iam <= CsrAccessPlugin_bus_write_bits[0];
        PrivilegedPlugin_logic_harts_0_m_edeleg_bp <= CsrAccessPlugin_bus_write_bits[3];
        PrivilegedPlugin_logic_harts_0_m_edeleg_eu <= CsrAccessPlugin_bus_write_bits[8];
        PrivilegedPlugin_logic_harts_0_m_edeleg_es <= CsrAccessPlugin_bus_write_bits[9];
        PrivilegedPlugin_logic_harts_0_m_edeleg_ipf <= CsrAccessPlugin_bus_write_bits[12];
        PrivilegedPlugin_logic_harts_0_m_edeleg_lpf <= CsrAccessPlugin_bus_write_bits[13];
        PrivilegedPlugin_logic_harts_0_m_edeleg_spf <= CsrAccessPlugin_bus_write_bits[15];
      end
      if(when_CsrAccessPlugin_l359_5) begin
        PrivilegedPlugin_logic_harts_0_m_ideleg_se <= CsrAccessPlugin_bus_write_bits[9];
        PrivilegedPlugin_logic_harts_0_m_ideleg_st <= CsrAccessPlugin_bus_write_bits[5];
        PrivilegedPlugin_logic_harts_0_m_ideleg_ss <= CsrAccessPlugin_bus_write_bits[1];
      end
      if(when_CsrAccessPlugin_l359_6) begin
        PrivilegedPlugin_logic_harts_0_s_cause_interrupt <= CsrAccessPlugin_bus_write_bits[31];
        PrivilegedPlugin_logic_harts_0_s_cause_code <= CsrAccessPlugin_bus_write_bits[3 : 0];
      end
      if(when_CsrAccessPlugin_l359_7) begin
        PrivilegedPlugin_logic_harts_0_s_status_spp <= CsrAccessPlugin_bus_write_bits[8 : 8];
        PrivilegedPlugin_logic_harts_0_s_status_spie <= CsrAccessPlugin_bus_write_bits[5];
        PrivilegedPlugin_logic_harts_0_s_status_sie <= CsrAccessPlugin_bus_write_bits[1];
        PrivilegedPlugin_logic_harts_0_m_status_fs <= CsrAccessPlugin_bus_write_bits[14 : 13];
        MmuPlugin_logic_status_mxr <= CsrAccessPlugin_bus_write_bits[19];
        MmuPlugin_logic_status_sum <= CsrAccessPlugin_bus_write_bits[18];
      end
      if(when_CsrAccessPlugin_l359_8) begin
        if(when_CsrService_l166) begin
          if(PrivilegedPlugin_logic_harts_0_m_ideleg_se) begin
            PrivilegedPlugin_logic_harts_0_s_ie_seie <= CsrAccessPlugin_bus_write_bits[9];
          end
        end
        if(when_CsrService_l166) begin
          if(PrivilegedPlugin_logic_harts_0_m_ideleg_st) begin
            PrivilegedPlugin_logic_harts_0_s_ie_stie <= CsrAccessPlugin_bus_write_bits[5];
          end
        end
        if(when_CsrService_l166) begin
          if(PrivilegedPlugin_logic_harts_0_m_ideleg_ss) begin
            PrivilegedPlugin_logic_harts_0_s_ie_ssie <= CsrAccessPlugin_bus_write_bits[1];
          end
        end
      end
      if(when_CsrAccessPlugin_l359_9) begin
        if(when_CsrService_l166) begin
          if(PrivilegedPlugin_logic_harts_0_m_ideleg_ss) begin
            PrivilegedPlugin_logic_harts_0_s_ip_ssip <= CsrAccessPlugin_bus_write_bits[1];
          end
        end
      end
      if(when_CsrAccessPlugin_l366) begin
        if(when_CsrAccessPlugin_l359_10) begin
          MmuPlugin_logic_satp_mode <= CsrAccessPlugin_bus_write_bits[31 : 31];
          MmuPlugin_logic_satp_ppn <= CsrAccessPlugin_bus_write_bits[19 : 0];
        end
      end
      HistoryPlugin_logic_onFetch_value <= HistoryPlugin_logic_onFetch_valueNext;
      CsrRamPlugin_logic_readLogic_ohReg <= (CsrRamPlugin_logic_readLogic_port_cmd_valid ? CsrRamPlugin_logic_readLogic_oh : 2'b00);
      CsrRamPlugin_logic_readLogic_busy <= CsrRamPlugin_logic_readLogic_port_cmd_valid;
      CsrRamPlugin_logic_flush_counter <= (CsrRamPlugin_logic_flush_counter + _zz_CsrRamPlugin_logic_flush_counter);
      if(when_RegFilePlugin_l127) begin
        integer_RegFilePlugin_logic_initalizer_counter <= (integer_RegFilePlugin_logic_initalizer_counter + 6'h01);
      end
      _zz_WhiteboxerPlugin_logic_perf_executeFreezedCounter_2 <= _zz_WhiteboxerPlugin_logic_perf_executeFreezedCounter_1;
      _zz_WhiteboxerPlugin_logic_perf_dispatchHazardsCounter_2 <= _zz_WhiteboxerPlugin_logic_perf_dispatchHazardsCounter_1;
      _zz_WhiteboxerPlugin_logic_perf_candidatesCountCounters_0_2 <= _zz_WhiteboxerPlugin_logic_perf_candidatesCountCounters_0_1;
      _zz_WhiteboxerPlugin_logic_perf_candidatesCountCounters_1_2 <= _zz_WhiteboxerPlugin_logic_perf_candidatesCountCounters_1_1;
      _zz_WhiteboxerPlugin_logic_perf_candidatesCountCounters_2_2 <= _zz_WhiteboxerPlugin_logic_perf_candidatesCountCounters_2_1;
      _zz_WhiteboxerPlugin_logic_perf_candidatesCountCounters_3_2 <= _zz_WhiteboxerPlugin_logic_perf_candidatesCountCounters_3_1;
      _zz_WhiteboxerPlugin_logic_perf_dispatchFeedCounters_0_2 <= _zz_WhiteboxerPlugin_logic_perf_dispatchFeedCounters_0_1;
      _zz_WhiteboxerPlugin_logic_perf_dispatchFeedCounters_1_2 <= _zz_WhiteboxerPlugin_logic_perf_dispatchFeedCounters_1_1;
      _zz_WhiteboxerPlugin_logic_perf_dispatchFeedCounters_2_2 <= _zz_WhiteboxerPlugin_logic_perf_dispatchFeedCounters_2_1;
      if(fetch_logic_ctrls_1_up_forgetOne) begin
        fetch_logic_ctrls_1_up_valid <= 1'b0;
      end
      if(fetch_logic_ctrls_0_down_isReady) begin
        fetch_logic_ctrls_1_up_valid <= fetch_logic_ctrls_0_down_isValid;
      end
      if(fetch_logic_ctrls_2_up_forgetOne) begin
        fetch_logic_ctrls_2_up_valid <= 1'b0;
      end
      if(fetch_logic_ctrls_1_down_isReady) begin
        fetch_logic_ctrls_2_up_valid <= fetch_logic_ctrls_1_down_isValid;
      end
      if(toplevel_decode_ctrls_0_down_isReady) begin
        toplevel_decode_ctrls_1_up_valid <= toplevel_decode_ctrls_0_down_isValid;
      end
      if(toplevel_decode_ctrls_0_down_isReady) begin
        toplevel_decode_ctrls_1_up_LANE_SEL_0 <= toplevel_decode_ctrls_0_down_LANE_SEL_0;
        toplevel_decode_ctrls_1_up_LANE_SEL_1 <= toplevel_decode_ctrls_0_down_LANE_SEL_1;
      end
      if(when_DecodePipelinePlugin_l68) begin
        toplevel_decode_ctrls_1_up_LANE_SEL_0 <= 1'b0;
      end
      if(when_DecodePipelinePlugin_l68_1) begin
        toplevel_decode_ctrls_1_up_LANE_SEL_1 <= 1'b0;
      end
      if(toplevel_execute_ctrl0_down_isReady) begin
        toplevel_execute_ctrl1_up_LANE_SEL_lane0 <= toplevel_execute_ctrl0_down_LANE_SEL_lane0;
        toplevel_execute_ctrl1_up_LANE_SEL_lane1 <= toplevel_execute_ctrl0_down_LANE_SEL_lane1;
      end
      if(toplevel_execute_ctrl1_down_isReady) begin
        toplevel_execute_ctrl2_up_LANE_SEL_lane0 <= toplevel_execute_ctrl1_down_LANE_SEL_lane0;
        toplevel_execute_ctrl2_up_LANE_SEL_lane1 <= toplevel_execute_ctrl1_down_LANE_SEL_lane1;
      end
      if(toplevel_execute_ctrl2_down_isReady) begin
        toplevel_execute_ctrl3_up_LANE_SEL_lane0 <= toplevel_execute_ctrl2_down_LANE_SEL_lane0;
        toplevel_execute_ctrl3_up_LANE_SEL_lane1 <= toplevel_execute_ctrl2_down_LANE_SEL_lane1;
        toplevel_execute_ctrl3_up_LsuL1_SEL_lane0 <= toplevel_execute_ctrl2_down_LsuL1_SEL_lane0;
      end
      if(toplevel_execute_ctrl3_down_isReady) begin
        toplevel_execute_ctrl4_up_LANE_SEL_lane0 <= toplevel_execute_ctrl3_down_LANE_SEL_lane0;
        toplevel_execute_ctrl4_up_LANE_SEL_lane1 <= toplevel_execute_ctrl3_down_LANE_SEL_lane1;
        toplevel_execute_ctrl4_up_LsuL1_SEL_lane0 <= toplevel_execute_ctrl3_down_LsuL1_SEL_lane0;
      end
      if(toplevel_execute_ctrl4_down_isReady) begin
        toplevel_execute_ctrl5_up_LANE_SEL_lane0 <= toplevel_execute_ctrl4_down_LANE_SEL_lane0;
        toplevel_execute_ctrl5_up_LANE_SEL_lane1 <= toplevel_execute_ctrl4_down_LANE_SEL_lane1;
      end
      LsuPlugin_logic_flusher_stateReg <= LsuPlugin_logic_flusher_stateNext;
      TrapPlugin_logic_harts_0_trap_fsm_stateReg <= TrapPlugin_logic_harts_0_trap_fsm_stateNext;
      case(TrapPlugin_logic_harts_0_trap_fsm_stateReg)
        TrapPlugin_logic_harts_0_trap_fsm_enumDef_RUNNING : begin
        end
        TrapPlugin_logic_harts_0_trap_fsm_enumDef_PROCESS_1 : begin
          TrapPlugin_logic_harts_0_trap_fsm_trapEnterDebug <= 1'b0;
          if(!when_TrapPlugin_l393) begin
            case(TrapPlugin_logic_harts_0_trap_pending_state_code)
              4'b0000 : begin
                `ifndef SYNTHESIS
                  `ifdef FORMAL
                    assert((! TrapPlugin_logic_harts_0_trap_fsm_buffer_i_valid)); // TrapPlugin.scala:L415
                  `else
                    if(!(! TrapPlugin_logic_harts_0_trap_fsm_buffer_i_valid)) begin
                      $display("FAILURE "); // TrapPlugin.scala:L415
                      $finish;
                    end
                  `endif
                `endif
              end
              4'b0001 : begin
              end
              4'b0010 : begin
              end
              4'b0100 : begin
              end
              4'b0101 : begin
              end
              4'b1000 : begin
              end
              4'b0110 : begin
              end
              4'b0111 : begin
              end
              default : begin
                `ifndef SYNTHESIS
                  `ifdef FORMAL
                    assert(1'b0); // TrapPlugin.scala:L466
                  `else
                    if(!1'b0) begin
                      $display("FAILURE Unexpected trap reason"); // TrapPlugin.scala:L466
                      $finish;
                    end
                  `endif
                `endif
              end
            endcase
          end
        end
        TrapPlugin_logic_harts_0_trap_fsm_enumDef_TRAP_EPC : begin
        end
        TrapPlugin_logic_harts_0_trap_fsm_enumDef_TRAP_TVAL : begin
        end
        TrapPlugin_logic_harts_0_trap_fsm_enumDef_TRAP_TVEC : begin
        end
        TrapPlugin_logic_harts_0_trap_fsm_enumDef_TRAP_APPLY : begin
          PrivilegedPlugin_logic_harts_0_privilege <= TrapPlugin_logic_harts_0_trap_fsm_buffer_trap_targetPrivilege;
          case(TrapPlugin_logic_harts_0_trap_fsm_buffer_trap_targetPrivilege)
            2'b11 : begin
              PrivilegedPlugin_logic_harts_0_m_status_mie <= 1'b0;
              PrivilegedPlugin_logic_harts_0_m_status_mpie <= PrivilegedPlugin_logic_harts_0_m_status_mie;
              PrivilegedPlugin_logic_harts_0_m_status_mpp <= PrivilegedPlugin_logic_harts_0_privilege;
              PrivilegedPlugin_logic_harts_0_m_cause_code <= TrapPlugin_logic_harts_0_trap_fsm_buffer_trap_code;
              PrivilegedPlugin_logic_harts_0_m_cause_interrupt <= TrapPlugin_logic_harts_0_trap_fsm_buffer_trap_interrupt;
            end
            2'b01 : begin
              PrivilegedPlugin_logic_harts_0_s_status_sie <= 1'b0;
              PrivilegedPlugin_logic_harts_0_s_status_spie <= PrivilegedPlugin_logic_harts_0_s_status_sie;
              PrivilegedPlugin_logic_harts_0_s_status_spp <= PrivilegedPlugin_logic_harts_0_privilege[0 : 0];
              PrivilegedPlugin_logic_harts_0_s_cause_code <= TrapPlugin_logic_harts_0_trap_fsm_buffer_trap_code;
              PrivilegedPlugin_logic_harts_0_s_cause_interrupt <= TrapPlugin_logic_harts_0_trap_fsm_buffer_trap_interrupt;
            end
            default : begin
            end
          endcase
        end
        TrapPlugin_logic_harts_0_trap_fsm_enumDef_XRET_EPC : begin
        end
        TrapPlugin_logic_harts_0_trap_fsm_enumDef_XRET_APPLY : begin
          PrivilegedPlugin_logic_harts_0_privilege <= TrapPlugin_logic_harts_0_trap_pending_xret_targetPrivilege;
          case(switch_TrapPlugin_l638)
            2'b11 : begin
              PrivilegedPlugin_logic_harts_0_m_status_mpp <= 2'b00;
              PrivilegedPlugin_logic_harts_0_m_status_mie <= PrivilegedPlugin_logic_harts_0_m_status_mpie;
              PrivilegedPlugin_logic_harts_0_m_status_mpie <= 1'b1;
            end
            2'b01 : begin
              PrivilegedPlugin_logic_harts_0_s_status_spp <= 1'b0;
              PrivilegedPlugin_logic_harts_0_s_status_sie <= PrivilegedPlugin_logic_harts_0_s_status_spie;
              PrivilegedPlugin_logic_harts_0_s_status_spie <= 1'b1;
            end
            default : begin
            end
          endcase
        end
        TrapPlugin_logic_harts_0_trap_fsm_enumDef_ATS_RSP : begin
        end
        TrapPlugin_logic_harts_0_trap_fsm_enumDef_JUMP : begin
        end
        TrapPlugin_logic_harts_0_trap_fsm_enumDef_LSU_FLUSH : begin
        end
        TrapPlugin_logic_harts_0_trap_fsm_enumDef_FETCH_FLUSH : begin
        end
        default : begin
        end
      endcase
      MmuPlugin_logic_refill_stateReg <= MmuPlugin_logic_refill_stateNext;
      CsrAccessPlugin_logic_fsm_stateReg <= CsrAccessPlugin_logic_fsm_stateNext;
      case(CsrAccessPlugin_logic_fsm_stateReg)
        CsrAccessPlugin_logic_fsm_enumDef_READ : begin
        end
        CsrAccessPlugin_logic_fsm_enumDef_WRITE : begin
        end
        CsrAccessPlugin_logic_fsm_enumDef_COMPLETION : begin
        end
        default : begin
          if(CsrAccessPlugin_logic_fsm_inject_onDecodeDo) begin
            if(CsrAccessPlugin_logic_fsm_inject_sampled) begin
              if(CsrAccessPlugin_logic_fsm_inject_trapReg) begin
                CsrAccessPlugin_logic_fsm_inject_unfreeze <= execute_freeze_valid;
              end
            end
          end
        end
      endcase
      case(CsrAccessPlugin_logic_fsm_stateNext)
        CsrAccessPlugin_logic_fsm_enumDef_READ : begin
        end
        CsrAccessPlugin_logic_fsm_enumDef_WRITE : begin
        end
        CsrAccessPlugin_logic_fsm_enumDef_COMPLETION : begin
          CsrAccessPlugin_logic_fsm_inject_unfreeze <= 1'b1;
        end
        default : begin
        end
      endcase
      BtbPlugin_logic_ras_ptr_pop <= BtbPlugin_logic_ras_ptr_pop_aheadValue;
    end
  end

  always @(posedge clk_cpu) begin
    early0_MulPlugin_logic_writeback_buffer_data <= toplevel_execute_ctrl4_down_early0_MulPlugin_logic_steps_1_adders_0_lane0[63 : 32];
    early0_DivPlugin_logic_processing_divRevertResult <= ((toplevel_execute_ctrl2_down_RsUnsignedPlugin_RS1_REVERT_lane0 ^ (toplevel_execute_ctrl2_down_RsUnsignedPlugin_RS2_REVERT_lane0 && (! toplevel_execute_ctrl2_down_DivPlugin_REM_lane0))) && (! (((toplevel_execute_ctrl2_down_RsUnsignedPlugin_RS2_FORMATED_lane0 == 32'h0) && toplevel_execute_ctrl2_down_RsUnsignedPlugin_RS2_SIGNED_lane0) && (! toplevel_execute_ctrl2_down_DivPlugin_REM_lane0))));
    early0_DivPlugin_logic_processing_a_delay_1 <= early0_DivPlugin_logic_processing_a;
    early0_DivPlugin_logic_processing_b_delay_1 <= early0_DivPlugin_logic_processing_b;
    if(when_AlignerPlugin_l259) begin
      AlignerPlugin_logic_buffer_data <= fetch_logic_ctrls_2_down_Fetch_WORD;
      AlignerPlugin_logic_buffer_pc <= fetch_logic_ctrls_2_down_Fetch_WORD_PC;
      AlignerPlugin_logic_buffer_hm_Fetch_ID <= fetch_logic_ctrls_2_down_Fetch_ID;
      AlignerPlugin_logic_buffer_hm_GSharePlugin_GSHARE_COUNTER_0 <= fetch_logic_ctrls_2_down_GSharePlugin_GSHARE_COUNTER_0;
      AlignerPlugin_logic_buffer_hm_GSharePlugin_GSHARE_COUNTER_1 <= fetch_logic_ctrls_2_down_GSharePlugin_GSHARE_COUNTER_1;
      AlignerPlugin_logic_buffer_hm_GSharePlugin_GSHARE_COUNTER_2 <= fetch_logic_ctrls_2_down_GSharePlugin_GSHARE_COUNTER_2;
      AlignerPlugin_logic_buffer_hm_GSharePlugin_GSHARE_COUNTER_3 <= fetch_logic_ctrls_2_down_GSharePlugin_GSHARE_COUNTER_3;
      AlignerPlugin_logic_buffer_hm_Prediction_BRANCH_HISTORY <= fetch_logic_ctrls_2_down_Prediction_BRANCH_HISTORY;
      AlignerPlugin_logic_buffer_hm_Prediction_WORD_SLICES_BRANCH <= fetch_logic_ctrls_2_down_Prediction_WORD_SLICES_BRANCH;
      AlignerPlugin_logic_buffer_hm_Prediction_WORD_SLICES_TAKEN <= fetch_logic_ctrls_2_down_Prediction_WORD_SLICES_TAKEN;
      AlignerPlugin_logic_buffer_hm_Prediction_WORD_JUMP_PC <= fetch_logic_ctrls_2_down_Prediction_WORD_JUMP_PC;
      AlignerPlugin_logic_buffer_hm_Prediction_WORD_JUMPED <= fetch_logic_ctrls_2_down_Prediction_WORD_JUMPED;
      AlignerPlugin_logic_buffer_hm_Prediction_WORD_JUMP_SLICE <= fetch_logic_ctrls_2_down_Prediction_WORD_JUMP_SLICE;
    end
    if(when_FetchL1Plugin_l271) begin
      if(_zz_when) begin
        FetchL1Plugin_logic_refill_slots_0_address <= FetchL1Plugin_logic_refill_start_address;
        FetchL1Plugin_logic_refill_slots_0_isIo <= FetchL1Plugin_logic_refill_start_isIo;
        FetchL1Plugin_logic_refill_slots_0_wayToAllocate <= FetchL1Plugin_logic_refill_start_wayToAllocate;
        FetchL1Plugin_logic_refill_slots_0_priority <= FetchL1Plugin_logic_refill_slots_0_valid;
      end
    end
    FetchL1Plugin_logic_ctrl_plruLogic_buffer_regNext_payload_address <= FetchL1Plugin_logic_ctrl_plruLogic_buffer_payload_address;
    FetchL1Plugin_logic_ctrl_plruLogic_buffer_regNext_payload_data_0 <= FetchL1Plugin_logic_ctrl_plruLogic_buffer_payload_data_0;
    PrivilegedPlugin_logic_harts_0_s_ip_seipInput <= PrivilegedPlugin_logic_harts_0_int_s_external;
    if(BtbPlugin_logic_ras_readIt) begin
      BtbPlugin_logic_ras_read <= BtbPlugin_logic_ras_mem_stack_spinal_port0;
    end
    if(late0_BranchPlugin_logic_jumpLogic_learn_ready) begin
      late0_BranchPlugin_logic_jumpLogic_learn_rData_pcOnLastSlice <= late0_BranchPlugin_logic_jumpLogic_learn_payload_pcOnLastSlice;
      late0_BranchPlugin_logic_jumpLogic_learn_rData_pcTarget <= late0_BranchPlugin_logic_jumpLogic_learn_payload_pcTarget;
      late0_BranchPlugin_logic_jumpLogic_learn_rData_taken <= late0_BranchPlugin_logic_jumpLogic_learn_payload_taken;
      late0_BranchPlugin_logic_jumpLogic_learn_rData_isBranch <= late0_BranchPlugin_logic_jumpLogic_learn_payload_isBranch;
      late0_BranchPlugin_logic_jumpLogic_learn_rData_isPush <= late0_BranchPlugin_logic_jumpLogic_learn_payload_isPush;
      late0_BranchPlugin_logic_jumpLogic_learn_rData_isPop <= late0_BranchPlugin_logic_jumpLogic_learn_payload_isPop;
      late0_BranchPlugin_logic_jumpLogic_learn_rData_wasWrong <= late0_BranchPlugin_logic_jumpLogic_learn_payload_wasWrong;
      late0_BranchPlugin_logic_jumpLogic_learn_rData_badPredictedTarget <= late0_BranchPlugin_logic_jumpLogic_learn_payload_badPredictedTarget;
      late0_BranchPlugin_logic_jumpLogic_learn_rData_history <= late0_BranchPlugin_logic_jumpLogic_learn_payload_history;
      late0_BranchPlugin_logic_jumpLogic_learn_rData_uopId <= late0_BranchPlugin_logic_jumpLogic_learn_payload_uopId;
      late0_BranchPlugin_logic_jumpLogic_learn_rData_ctx_GSharePlugin_GSHARE_COUNTER_0 <= late0_BranchPlugin_logic_jumpLogic_learn_payload_ctx_GSharePlugin_GSHARE_COUNTER_0;
      late0_BranchPlugin_logic_jumpLogic_learn_rData_ctx_GSharePlugin_GSHARE_COUNTER_1 <= late0_BranchPlugin_logic_jumpLogic_learn_payload_ctx_GSharePlugin_GSHARE_COUNTER_1;
      late0_BranchPlugin_logic_jumpLogic_learn_rData_ctx_GSharePlugin_GSHARE_COUNTER_2 <= late0_BranchPlugin_logic_jumpLogic_learn_payload_ctx_GSharePlugin_GSHARE_COUNTER_2;
      late0_BranchPlugin_logic_jumpLogic_learn_rData_ctx_GSharePlugin_GSHARE_COUNTER_3 <= late0_BranchPlugin_logic_jumpLogic_learn_payload_ctx_GSharePlugin_GSHARE_COUNTER_3;
    end
    if(late1_BranchPlugin_logic_jumpLogic_learn_ready) begin
      late1_BranchPlugin_logic_jumpLogic_learn_rData_pcOnLastSlice <= late1_BranchPlugin_logic_jumpLogic_learn_payload_pcOnLastSlice;
      late1_BranchPlugin_logic_jumpLogic_learn_rData_pcTarget <= late1_BranchPlugin_logic_jumpLogic_learn_payload_pcTarget;
      late1_BranchPlugin_logic_jumpLogic_learn_rData_taken <= late1_BranchPlugin_logic_jumpLogic_learn_payload_taken;
      late1_BranchPlugin_logic_jumpLogic_learn_rData_isBranch <= late1_BranchPlugin_logic_jumpLogic_learn_payload_isBranch;
      late1_BranchPlugin_logic_jumpLogic_learn_rData_isPush <= late1_BranchPlugin_logic_jumpLogic_learn_payload_isPush;
      late1_BranchPlugin_logic_jumpLogic_learn_rData_isPop <= late1_BranchPlugin_logic_jumpLogic_learn_payload_isPop;
      late1_BranchPlugin_logic_jumpLogic_learn_rData_wasWrong <= late1_BranchPlugin_logic_jumpLogic_learn_payload_wasWrong;
      late1_BranchPlugin_logic_jumpLogic_learn_rData_badPredictedTarget <= late1_BranchPlugin_logic_jumpLogic_learn_payload_badPredictedTarget;
      late1_BranchPlugin_logic_jumpLogic_learn_rData_history <= late1_BranchPlugin_logic_jumpLogic_learn_payload_history;
      late1_BranchPlugin_logic_jumpLogic_learn_rData_uopId <= late1_BranchPlugin_logic_jumpLogic_learn_payload_uopId;
      late1_BranchPlugin_logic_jumpLogic_learn_rData_ctx_GSharePlugin_GSHARE_COUNTER_0 <= late1_BranchPlugin_logic_jumpLogic_learn_payload_ctx_GSharePlugin_GSHARE_COUNTER_0;
      late1_BranchPlugin_logic_jumpLogic_learn_rData_ctx_GSharePlugin_GSHARE_COUNTER_1 <= late1_BranchPlugin_logic_jumpLogic_learn_payload_ctx_GSharePlugin_GSHARE_COUNTER_1;
      late1_BranchPlugin_logic_jumpLogic_learn_rData_ctx_GSharePlugin_GSHARE_COUNTER_2 <= late1_BranchPlugin_logic_jumpLogic_learn_payload_ctx_GSharePlugin_GSHARE_COUNTER_2;
      late1_BranchPlugin_logic_jumpLogic_learn_rData_ctx_GSharePlugin_GSHARE_COUNTER_3 <= late1_BranchPlugin_logic_jumpLogic_learn_payload_ctx_GSharePlugin_GSHARE_COUNTER_3;
    end
    if(DispatchPlugin_logic_slotsFeeds_doIt) begin
      DispatchPlugin_logic_slots_0_ctx_laneLayerHits <= _zz_DispatchPlugin_logic_slots_0_ctx_valid_4[4 : 1];
      DispatchPlugin_logic_slots_0_ctx_uop <= _zz_DispatchPlugin_logic_slots_0_ctx_valid_4[36 : 5];
      DispatchPlugin_logic_slots_0_ctx_hm_Prediction_ALIGNED_JUMPED <= _zz_DispatchPlugin_logic_slots_0_ctx_hm_Prediction_ALIGNED_JUMPED[0];
      DispatchPlugin_logic_slots_0_ctx_hm_Prediction_ALIGNED_JUMPED_PC <= _zz_DispatchPlugin_logic_slots_0_ctx_hm_Prediction_ALIGNED_JUMPED[32 : 1];
      DispatchPlugin_logic_slots_0_ctx_hm_Prediction_ALIGNED_SLICES_TAKEN <= _zz_DispatchPlugin_logic_slots_0_ctx_hm_Prediction_ALIGNED_JUMPED[36 : 33];
      DispatchPlugin_logic_slots_0_ctx_hm_Prediction_ALIGNED_SLICES_BRANCH <= _zz_DispatchPlugin_logic_slots_0_ctx_hm_Prediction_ALIGNED_JUMPED[40 : 37];
      DispatchPlugin_logic_slots_0_ctx_hm_GSharePlugin_GSHARE_COUNTER_0 <= _zz_DispatchPlugin_logic_slots_0_ctx_hm_GSharePlugin_GSHARE_COUNTER_0[1 : 0];
      DispatchPlugin_logic_slots_0_ctx_hm_GSharePlugin_GSHARE_COUNTER_1 <= _zz_DispatchPlugin_logic_slots_0_ctx_hm_GSharePlugin_GSHARE_COUNTER_0[3 : 2];
      DispatchPlugin_logic_slots_0_ctx_hm_GSharePlugin_GSHARE_COUNTER_2 <= _zz_DispatchPlugin_logic_slots_0_ctx_hm_GSharePlugin_GSHARE_COUNTER_0[5 : 4];
      DispatchPlugin_logic_slots_0_ctx_hm_GSharePlugin_GSHARE_COUNTER_3 <= _zz_DispatchPlugin_logic_slots_0_ctx_hm_GSharePlugin_GSHARE_COUNTER_0[7 : 6];
      DispatchPlugin_logic_slots_0_ctx_hm_Prediction_BRANCH_HISTORY <= _zz_DispatchPlugin_logic_slots_0_ctx_hm_Prediction_ALIGNED_JUMPED[60 : 49];
      DispatchPlugin_logic_slots_0_ctx_hm_DispatchPlugin_FENCE_OLDER <= _zz_DispatchPlugin_logic_slots_0_ctx_hm_Prediction_ALIGNED_JUMPED[61];
      DispatchPlugin_logic_slots_0_ctx_hm_DispatchPlugin_MAY_FLUSH <= _zz_DispatchPlugin_logic_slots_0_ctx_hm_Prediction_ALIGNED_JUMPED[62];
      DispatchPlugin_logic_slots_0_ctx_hm_DispatchPlugin_DONT_FLUSH <= _zz_DispatchPlugin_logic_slots_0_ctx_hm_Prediction_ALIGNED_JUMPED[63];
      DispatchPlugin_logic_slots_0_ctx_hm_DispatchPlugin_DONT_FLUSH_FROM_LANES <= _zz_DispatchPlugin_logic_slots_0_ctx_hm_Prediction_ALIGNED_JUMPED[64];
      DispatchPlugin_logic_slots_0_ctx_hm_Decode_INSTRUCTION_SLICE_COUNT <= _zz_DispatchPlugin_logic_slots_0_ctx_hm_Prediction_ALIGNED_JUMPED[65 : 65];
      DispatchPlugin_logic_slots_0_ctx_hm_DONT_FLUSH_PRECISE_3 <= _zz_DispatchPlugin_logic_slots_0_ctx_hm_Prediction_ALIGNED_JUMPED[66];
      DispatchPlugin_logic_slots_0_ctx_hm_DONT_FLUSH_PRECISE_4 <= _zz_DispatchPlugin_logic_slots_0_ctx_hm_Prediction_ALIGNED_JUMPED[67];
      DispatchPlugin_logic_slots_0_ctx_hm_PC <= _zz_DispatchPlugin_logic_slots_0_ctx_hm_Prediction_ALIGNED_JUMPED[99 : 68];
      DispatchPlugin_logic_slots_0_ctx_hm_TRAP <= _zz_DispatchPlugin_logic_slots_0_ctx_hm_Prediction_ALIGNED_JUMPED[100];
      DispatchPlugin_logic_slots_0_ctx_hm_Decode_UOP_ID <= _zz_DispatchPlugin_logic_slots_0_ctx_hm_Prediction_ALIGNED_JUMPED[116 : 101];
      DispatchPlugin_logic_slots_0_ctx_hm_RS1_ENABLE <= _zz_DispatchPlugin_logic_slots_0_ctx_hm_Prediction_ALIGNED_JUMPED[117];
      DispatchPlugin_logic_slots_0_ctx_hm_RS1_PHYS <= _zz_DispatchPlugin_logic_slots_0_ctx_hm_Prediction_ALIGNED_JUMPED[122 : 118];
      DispatchPlugin_logic_slots_0_ctx_hm_RS2_ENABLE <= _zz_DispatchPlugin_logic_slots_0_ctx_hm_Prediction_ALIGNED_JUMPED[123];
      DispatchPlugin_logic_slots_0_ctx_hm_RS2_PHYS <= _zz_DispatchPlugin_logic_slots_0_ctx_hm_Prediction_ALIGNED_JUMPED[128 : 124];
      DispatchPlugin_logic_slots_0_ctx_hm_RD_ENABLE <= _zz_DispatchPlugin_logic_slots_0_ctx_hm_Prediction_ALIGNED_JUMPED[129];
      DispatchPlugin_logic_slots_0_ctx_hm_RD_PHYS <= _zz_DispatchPlugin_logic_slots_0_ctx_hm_Prediction_ALIGNED_JUMPED[134 : 130];
      DispatchPlugin_logic_slots_0_ctx_hm_DispatchPlugin_logic_hcs_0_onRs_0_ENABLES_0 <= _zz_DispatchPlugin_logic_slots_0_ctx_hm_Prediction_ALIGNED_JUMPED[135];
      DispatchPlugin_logic_slots_0_ctx_hm_DispatchPlugin_logic_hcs_0_onRs_1_ENABLES_0 <= _zz_DispatchPlugin_logic_slots_0_ctx_hm_Prediction_ALIGNED_JUMPED[136];
      DispatchPlugin_logic_slots_0_ctx_hm_DispatchPlugin_logic_hcs_1_onRs_0_ENABLES_0 <= _zz_DispatchPlugin_logic_slots_0_ctx_hm_Prediction_ALIGNED_JUMPED[137];
      DispatchPlugin_logic_slots_0_ctx_hm_DispatchPlugin_logic_hcs_1_onRs_1_ENABLES_0 <= _zz_DispatchPlugin_logic_slots_0_ctx_hm_Prediction_ALIGNED_JUMPED[138];
      DispatchPlugin_logic_slots_0_ctx_hm_DispatchPlugin_logic_hcs_1_onRs_1_ENABLES_1 <= _zz_DispatchPlugin_logic_slots_0_ctx_hm_Prediction_ALIGNED_JUMPED[139];
      DispatchPlugin_logic_slots_0_ctx_hm_DispatchPlugin_logic_hcs_2_onRs_0_ENABLES_0 <= _zz_DispatchPlugin_logic_slots_0_ctx_hm_Prediction_ALIGNED_JUMPED[140];
      DispatchPlugin_logic_slots_0_ctx_hm_DispatchPlugin_logic_hcs_2_onRs_1_ENABLES_0 <= _zz_DispatchPlugin_logic_slots_0_ctx_hm_Prediction_ALIGNED_JUMPED[141];
      DispatchPlugin_logic_slots_0_ctx_hm_DispatchPlugin_logic_hcs_3_onRs_0_ENABLES_0 <= _zz_DispatchPlugin_logic_slots_0_ctx_hm_Prediction_ALIGNED_JUMPED[142];
      DispatchPlugin_logic_slots_0_ctx_hm_DispatchPlugin_logic_hcs_3_onRs_1_ENABLES_0 <= _zz_DispatchPlugin_logic_slots_0_ctx_hm_Prediction_ALIGNED_JUMPED[143];
    end
    LsuL1Plugin_logic_refill_slots_0_loadedCounter <= (LsuL1Plugin_logic_refill_slots_0_loadedCounter + ((LsuL1Plugin_logic_refill_slots_0_loaded && (! LsuL1Plugin_logic_refill_slots_0_loadedDone)) && (! execute_freeze_valid)));
    if(LsuL1Plugin_logic_refill_push_valid) begin
      if(when_LsuL1Plugin_l358) begin
        LsuL1Plugin_logic_refill_slots_0_address <= LsuL1Plugin_logic_refill_push_payload_address;
        LsuL1Plugin_logic_refill_slots_0_way <= LsuL1Plugin_logic_refill_push_payload_way;
        LsuL1Plugin_logic_refill_slots_0_cmdSent <= 1'b0;
        LsuL1Plugin_logic_refill_slots_0_loadedCounter <= 1'b0;
        LsuL1Plugin_logic_refill_slots_0_victim <= LsuL1Plugin_logic_refill_push_payload_victim;
        LsuL1Plugin_logic_refill_slots_0_dirty <= LsuL1Plugin_logic_refill_push_payload_dirty;
      end
    end
    if(LsuL1Plugin_logic_refill_read_arbiter_oh[0]) begin
      if(LsuL1Plugin_logic_bus_read_cmd_ready) begin
        LsuL1Plugin_logic_refill_slots_0_cmdSent <= 1'b1;
      end
    end
    LsuL1Plugin_logic_writeback_slots_0_timer_counter <= (LsuL1Plugin_logic_writeback_slots_0_timer_counter + ((! LsuL1Plugin_logic_writeback_slots_0_timer_done) && (! execute_freeze_valid)));
    if(LsuL1Plugin_logic_writeback_push_valid) begin
      if(when_LsuL1Plugin_l532) begin
        LsuL1Plugin_logic_writeback_slots_0_address <= LsuL1Plugin_logic_writeback_push_payload_address;
        LsuL1Plugin_logic_writeback_slots_0_way <= LsuL1Plugin_logic_writeback_push_payload_way;
        LsuL1Plugin_logic_writeback_slots_0_timer_counter <= 1'b0;
        LsuL1Plugin_logic_writeback_slots_0_writeCmdDone <= 1'b0;
        LsuL1Plugin_logic_writeback_slots_0_readCmdDone <= 1'b0;
        LsuL1Plugin_logic_writeback_slots_0_readRspDone <= 1'b0;
        LsuL1Plugin_logic_writeback_slots_0_victimBufferReady <= 1'b0;
      end
    end
    if(when_LsuL1Plugin_l577) begin
      if(LsuL1Plugin_logic_writeback_read_arbiter_oh[0]) begin
        LsuL1Plugin_logic_writeback_slots_0_readCmdDone <= 1'b1;
      end
    end
    if(LsuL1Plugin_logic_writeback_read_slotRead_valid) begin
      LsuL1Plugin_logic_refill_slots_0_victim[0] <= 1'b0;
    end
    LsuL1Plugin_logic_writeback_read_slotReadLast_payload_last <= LsuL1Plugin_logic_writeback_read_slotRead_payload_last;
    LsuL1Plugin_logic_writeback_read_slotReadLast_payload_wordIndex <= LsuL1Plugin_logic_writeback_read_slotRead_payload_wordIndex;
    LsuL1Plugin_logic_writeback_read_slotReadLast_payload_way <= LsuL1Plugin_logic_writeback_read_slotRead_payload_way;
    if(LsuL1Plugin_logic_writeback_read_slotReadLast_valid) begin
      LsuL1Plugin_logic_writeback_slots_0_victimBufferReady <= 1'b1;
      if(LsuL1Plugin_logic_writeback_read_slotReadLast_payload_last) begin
        LsuL1Plugin_logic_writeback_slots_0_readRspDone <= 1'b1;
      end
    end
    if(when_LsuL1Plugin_l651) begin
      if(LsuL1Plugin_logic_writeback_write_arbiter_oh[0]) begin
        LsuL1Plugin_logic_writeback_slots_0_writeCmdDone <= 1'b1;
      end
    end
    if(LsuL1Plugin_logic_writeback_write_bufferRead_ready) begin
      LsuL1Plugin_logic_writeback_write_bufferRead_rData_address <= LsuL1Plugin_logic_writeback_write_bufferRead_payload_address;
      LsuL1Plugin_logic_writeback_write_bufferRead_rData_last <= LsuL1Plugin_logic_writeback_write_bufferRead_payload_last;
    end
    if(LsuPlugin_logic_onAddress0_flush_port_fire) begin
      LsuPlugin_logic_flusher_cmdCounter <= (LsuPlugin_logic_flusher_cmdCounter + 7'h01);
    end
    if(LsuPlugin_logic_bus_rsp_toStream_ready) begin
      LsuPlugin_logic_bus_rsp_toStream_rData_error <= LsuPlugin_logic_bus_rsp_toStream_payload_error;
      LsuPlugin_logic_bus_rsp_toStream_rData_data <= LsuPlugin_logic_bus_rsp_toStream_payload_data;
    end
    LsuPlugin_logic_onCtrl_rva_srcBuffer <= toplevel_execute_ctrl4_down_LsuPlugin_logic_onCtrl_loadData_RESULT_lane0;
    LsuPlugin_logic_onCtrl_rva_aluBuffer <= LsuPlugin_logic_onCtrl_rva_alu_result;
    _zz_LsuPlugin_logic_onCtrl_rva_delay_0 <= (! execute_freeze_valid);
    _zz_LsuPlugin_logic_onCtrl_rva_delay_1 <= _zz_LsuPlugin_logic_onCtrl_rva_delay_0;
    if(!when_LsuPlugin_l585) begin
      LsuPlugin_logic_onCtrl_rva_nc_age <= (LsuPlugin_logic_onCtrl_rva_nc_age + _zz_LsuPlugin_logic_onCtrl_rva_nc_age);
    end
    if(LsuPlugin_logic_onCtrl_rva_nc_capture) begin
      LsuPlugin_logic_onCtrl_rva_nc_address <= toplevel_execute_ctrl4_down_LsuL1_PHYSICAL_ADDRESS_lane0;
      LsuPlugin_logic_onCtrl_rva_nc_age <= 6'h0;
    end
    if(when_LsuPlugin_l761) begin
      LsuPlugin_logic_flusher_cmdCounter <= {1'd0, _zz_LsuPlugin_logic_flusher_cmdCounter};
    end
    if(when_LsuPlugin_l796) begin
      if(when_LsuPlugin_l204) begin
        LsuPlugin_logic_onAddress0_access_waiter_refill <= toplevel_execute_ctrl4_down_LsuL1_WAIT_REFILL_lane0;
      end
    end
    if(when_LsuPlugin_l803) begin
      if(when_LsuPlugin_l204_1) begin
        LsuPlugin_logic_onCtrl_hartRegulation_refill <= toplevel_execute_ctrl4_down_LsuL1_WAIT_REFILL_lane0;
      end
    end
    LsuL1Plugin_logic_bus_toTilelink_nonCoherent_onA_selReg <= LsuL1Plugin_logic_bus_toTilelink_nonCoherent_onA_sel;
    if(TrapPlugin_logic_harts_0_trap_pending_arbiter_down_valid) begin
      TrapPlugin_logic_harts_0_trap_pending_state_exception <= TrapPlugin_logic_harts_0_trap_pending_arbiter_down_payload_exception;
      TrapPlugin_logic_harts_0_trap_pending_state_tval <= TrapPlugin_logic_harts_0_trap_pending_arbiter_down_payload_tval;
      TrapPlugin_logic_harts_0_trap_pending_state_code <= TrapPlugin_logic_harts_0_trap_pending_arbiter_down_payload_code;
      TrapPlugin_logic_harts_0_trap_pending_state_arg <= TrapPlugin_logic_harts_0_trap_pending_arbiter_down_payload_arg;
    end
    if(TrapPlugin_logic_harts_0_trap_trigger_valid) begin
      TrapPlugin_logic_harts_0_trap_pending_pc <= ((_zz_TrapPlugin_logic_harts_0_trap_pending_pc ? toplevel_execute_ctrl4_down_PC_lane0 : 32'h0) | (_zz_TrapPlugin_logic_harts_0_trap_pending_pc_1 ? toplevel_execute_ctrl4_down_PC_lane1 : 32'h0));
      TrapPlugin_logic_harts_0_trap_pending_history <= ((_zz_TrapPlugin_logic_harts_0_trap_pending_pc ? toplevel_execute_ctrl4_down_Prediction_BRANCH_HISTORY_lane0 : 12'h0) | (_zz_TrapPlugin_logic_harts_0_trap_pending_pc_1 ? toplevel_execute_ctrl4_down_Prediction_BRANCH_HISTORY_lane1 : 12'h0));
      TrapPlugin_logic_harts_0_trap_pending_slices <= (_zz_TrapPlugin_logic_harts_0_trap_pending_slices + 2'b01);
    end
    if(TrapPlugin_logic_harts_0_trap_fsm_buffer_sampleIt) begin
      TrapPlugin_logic_harts_0_trap_fsm_buffer_i_valid <= TrapPlugin_logic_harts_0_interrupt_valid;
    end
    if(TrapPlugin_logic_harts_0_trap_fsm_buffer_sampleIt) begin
      TrapPlugin_logic_harts_0_trap_fsm_buffer_i_code <= TrapPlugin_logic_harts_0_interrupt_code;
    end
    if(TrapPlugin_logic_harts_0_trap_fsm_buffer_sampleIt) begin
      TrapPlugin_logic_harts_0_trap_fsm_buffer_i_targetPrivilege <= TrapPlugin_logic_harts_0_interrupt_targetPrivilege;
    end
    TrapPlugin_logic_harts_0_trap_fsm_jumpTarget <= (TrapPlugin_logic_harts_0_trap_pending_pc + _zz_TrapPlugin_logic_harts_0_trap_fsm_jumpTarget);
    if(when_TrapPlugin_l539) begin
      TrapPlugin_logic_harts_0_trap_fsm_readed <= TrapPlugin_logic_harts_0_crsPorts_read_data;
    end
    MmuPlugin_logic_refill_load_rsp_payload_data <= MmuPlugin_logic_accessBus_rsp_payload_data;
    MmuPlugin_logic_refill_load_rsp_payload_error <= MmuPlugin_logic_accessBus_rsp_payload_error;
    MmuPlugin_logic_refill_load_rsp_payload_redo <= MmuPlugin_logic_accessBus_rsp_payload_redo;
    MmuPlugin_logic_refill_load_rsp_payload_waitAny <= MmuPlugin_logic_accessBus_rsp_payload_waitAny;
    if(when_MmuPlugin_l496) begin
      MmuPlugin_logic_invalidate_counter <= 6'h0;
    end else begin
      MmuPlugin_logic_invalidate_counter <= (MmuPlugin_logic_invalidate_counter + 6'h01);
    end
    if(LsuTileLinkPlugin_logic_bridge_down_a_fire) begin
      LsuTileLinkPlugin_logic_bridge_pendings_0_hash <= LsuTileLinkPlugin_logic_bridge_cmdHash;
      LsuTileLinkPlugin_logic_bridge_pendings_0_mask <= LsuPlugin_logic_bus_cmd_payload_mask;
      LsuTileLinkPlugin_logic_bridge_pendings_0_io <= LsuPlugin_logic_bus_cmd_payload_io;
    end
    CsrAccessPlugin_logic_fsm_regs_read <= ((toplevel_execute_ctrl2_down_CsrAccessPlugin_SEL_lane0 && (! CsrAccessPlugin_logic_fsm_inject_trap)) && CsrAccessPlugin_logic_fsm_inject_csrRead);
    CsrAccessPlugin_logic_fsm_regs_write <= ((toplevel_execute_ctrl2_down_CsrAccessPlugin_SEL_lane0 && (! CsrAccessPlugin_logic_fsm_inject_trap)) && CsrAccessPlugin_logic_fsm_inject_csrWrite);
    CsrAccessPlugin_logic_fsm_inject_trapReg <= CsrAccessPlugin_logic_fsm_inject_trap;
    CsrAccessPlugin_logic_fsm_inject_busTrapReg <= CsrAccessPlugin_bus_decode_trap;
    CsrAccessPlugin_logic_fsm_inject_busTrapCodeReg <= CsrAccessPlugin_bus_decode_trapCode;
    CsrAccessPlugin_logic_fsm_regs_onWriteBits <= CsrAccessPlugin_logic_fsm_writeLogic_alu_result;
    if(fetch_logic_ctrls_0_down_isReady) begin
      fetch_logic_ctrls_1_up_Fetch_WORD_PC <= fetch_logic_ctrls_0_down_Fetch_WORD_PC;
      fetch_logic_ctrls_1_up_Fetch_PC_FAULT <= fetch_logic_ctrls_0_down_Fetch_PC_FAULT;
      fetch_logic_ctrls_1_up_Fetch_ID <= fetch_logic_ctrls_0_down_Fetch_ID;
      _zz_1 <= 1'b0;
      fetch_logic_ctrls_1_up_FetchL1Plugin_logic_cmd_PLRU_BYPASS_VALID <= fetch_logic_ctrls_0_down_FetchL1Plugin_logic_cmd_PLRU_BYPASS_VALID;
      fetch_logic_ctrls_1_up_FetchL1Plugin_logic_cmd_PLRU_BYPASS_DATA_0 <= fetch_logic_ctrls_0_down_FetchL1Plugin_logic_cmd_PLRU_BYPASS_DATA_0;
      fetch_logic_ctrls_1_up_FetchL1Plugin_logic_cmd_TAGS_UPDATE <= fetch_logic_ctrls_0_down_FetchL1Plugin_logic_cmd_TAGS_UPDATE;
      fetch_logic_ctrls_1_up_FetchL1Plugin_logic_cmd_TAGS_UPDATE_ADDRESS <= fetch_logic_ctrls_0_down_FetchL1Plugin_logic_cmd_TAGS_UPDATE_ADDRESS;
      fetch_logic_ctrls_1_up_GSharePlugin_logic_HASH <= fetch_logic_ctrls_0_down_GSharePlugin_logic_HASH;
      fetch_logic_ctrls_1_up_Prediction_BRANCH_HISTORY <= fetch_logic_ctrls_0_down_Prediction_BRANCH_HISTORY;
      fetch_logic_ctrls_1_up_GSharePlugin_logic_BYPASS_valid <= fetch_logic_ctrls_0_down_GSharePlugin_logic_BYPASS_valid;
      fetch_logic_ctrls_1_up_GSharePlugin_logic_BYPASS_payload_address <= fetch_logic_ctrls_0_down_GSharePlugin_logic_BYPASS_payload_address;
      fetch_logic_ctrls_1_up_GSharePlugin_logic_BYPASS_payload_data_0 <= fetch_logic_ctrls_0_down_GSharePlugin_logic_BYPASS_payload_data_0;
      fetch_logic_ctrls_1_up_GSharePlugin_logic_BYPASS_payload_data_1 <= fetch_logic_ctrls_0_down_GSharePlugin_logic_BYPASS_payload_data_1;
      fetch_logic_ctrls_1_up_GSharePlugin_logic_BYPASS_payload_data_2 <= fetch_logic_ctrls_0_down_GSharePlugin_logic_BYPASS_payload_data_2;
      fetch_logic_ctrls_1_up_GSharePlugin_logic_BYPASS_payload_data_3 <= fetch_logic_ctrls_0_down_GSharePlugin_logic_BYPASS_payload_data_3;
      fetch_logic_ctrls_1_up_BtbPlugin_logic_readCmd_HAZARDS <= fetch_logic_ctrls_0_down_BtbPlugin_logic_readCmd_HAZARDS;
    end
    if(fetch_logic_ctrls_1_down_isReady) begin
      fetch_logic_ctrls_2_up_Fetch_WORD_PC <= fetch_logic_ctrls_1_down_Fetch_WORD_PC;
      fetch_logic_ctrls_2_up_Fetch_PC_FAULT <= fetch_logic_ctrls_1_down_Fetch_PC_FAULT;
      fetch_logic_ctrls_2_up_Fetch_ID <= fetch_logic_ctrls_1_down_Fetch_ID;
      fetch_logic_ctrls_2_up_Prediction_BRANCH_HISTORY <= fetch_logic_ctrls_1_down_Prediction_BRANCH_HISTORY;
      fetch_logic_ctrls_2_up_FetchL1Plugin_logic_WAYS_TAGS_0_loaded <= fetch_logic_ctrls_1_down_FetchL1Plugin_logic_WAYS_TAGS_0_loaded;
      fetch_logic_ctrls_2_up_FetchL1Plugin_logic_WAYS_TAGS_0_error <= fetch_logic_ctrls_1_down_FetchL1Plugin_logic_WAYS_TAGS_0_error;
      fetch_logic_ctrls_2_up_FetchL1Plugin_logic_WAYS_TAGS_0_address <= fetch_logic_ctrls_1_down_FetchL1Plugin_logic_WAYS_TAGS_0_address;
      fetch_logic_ctrls_2_up_FetchL1Plugin_logic_WAYS_TAGS_1_loaded <= fetch_logic_ctrls_1_down_FetchL1Plugin_logic_WAYS_TAGS_1_loaded;
      fetch_logic_ctrls_2_up_FetchL1Plugin_logic_WAYS_TAGS_1_error <= fetch_logic_ctrls_1_down_FetchL1Plugin_logic_WAYS_TAGS_1_error;
      fetch_logic_ctrls_2_up_FetchL1Plugin_logic_WAYS_TAGS_1_address <= fetch_logic_ctrls_1_down_FetchL1Plugin_logic_WAYS_TAGS_1_address;
      fetch_logic_ctrls_2_up_FetchL1Plugin_logic_PLRU_BYPASSED_0 <= fetch_logic_ctrls_1_down_FetchL1Plugin_logic_PLRU_BYPASSED_0;
      fetch_logic_ctrls_2_up_FetchL1Plugin_logic_BANKS_MUXES_0 <= fetch_logic_ctrls_1_down_FetchL1Plugin_logic_BANKS_MUXES_0;
      fetch_logic_ctrls_2_up_FetchL1Plugin_logic_BANKS_MUXES_1 <= fetch_logic_ctrls_1_down_FetchL1Plugin_logic_BANKS_MUXES_1;
      fetch_logic_ctrls_2_up_FetchL1Plugin_logic_HAZARD <= fetch_logic_ctrls_1_down_FetchL1Plugin_logic_HAZARD;
      fetch_logic_ctrls_2_up_FetchL1Plugin_logic_WAYS_HITS_0 <= fetch_logic_ctrls_1_down_FetchL1Plugin_logic_WAYS_HITS_0;
      fetch_logic_ctrls_2_up_FetchL1Plugin_logic_WAYS_HITS_1 <= fetch_logic_ctrls_1_down_FetchL1Plugin_logic_WAYS_HITS_1;
      fetch_logic_ctrls_2_up_MMU_BYPASS_TRANSLATION <= fetch_logic_ctrls_1_down_MMU_BYPASS_TRANSLATION;
      fetch_logic_ctrls_2_up_FetchL1Plugin_logic_WAYS_HIT <= fetch_logic_ctrls_1_down_FetchL1Plugin_logic_WAYS_HIT;
      fetch_logic_ctrls_2_up_GSharePlugin_GSHARE_COUNTER_0 <= fetch_logic_ctrls_1_down_GSharePlugin_GSHARE_COUNTER_0;
      fetch_logic_ctrls_2_up_GSharePlugin_GSHARE_COUNTER_1 <= fetch_logic_ctrls_1_down_GSharePlugin_GSHARE_COUNTER_1;
      fetch_logic_ctrls_2_up_GSharePlugin_GSHARE_COUNTER_2 <= fetch_logic_ctrls_1_down_GSharePlugin_GSHARE_COUNTER_2;
      fetch_logic_ctrls_2_up_GSharePlugin_GSHARE_COUNTER_3 <= fetch_logic_ctrls_1_down_GSharePlugin_GSHARE_COUNTER_3;
      fetch_logic_ctrls_2_up_BtbPlugin_logic_chunksLogic_0_readRsp_ENTRY_hash <= fetch_logic_ctrls_1_down_BtbPlugin_logic_chunksLogic_0_readRsp_ENTRY_hash;
      fetch_logic_ctrls_2_up_BtbPlugin_logic_chunksLogic_0_readRsp_ENTRY_sliceLow <= fetch_logic_ctrls_1_down_BtbPlugin_logic_chunksLogic_0_readRsp_ENTRY_sliceLow;
      fetch_logic_ctrls_2_up_BtbPlugin_logic_chunksLogic_0_readRsp_ENTRY_pcTarget <= fetch_logic_ctrls_1_down_BtbPlugin_logic_chunksLogic_0_readRsp_ENTRY_pcTarget;
      fetch_logic_ctrls_2_up_BtbPlugin_logic_chunksLogic_0_readRsp_ENTRY_isBranch <= fetch_logic_ctrls_1_down_BtbPlugin_logic_chunksLogic_0_readRsp_ENTRY_isBranch;
      fetch_logic_ctrls_2_up_BtbPlugin_logic_chunksLogic_0_readRsp_ENTRY_isPush <= fetch_logic_ctrls_1_down_BtbPlugin_logic_chunksLogic_0_readRsp_ENTRY_isPush;
      fetch_logic_ctrls_2_up_BtbPlugin_logic_chunksLogic_0_readRsp_ENTRY_isPop <= fetch_logic_ctrls_1_down_BtbPlugin_logic_chunksLogic_0_readRsp_ENTRY_isPop;
      fetch_logic_ctrls_2_up_BtbPlugin_logic_chunksLogic_0_hitCalc_HIT <= fetch_logic_ctrls_1_down_BtbPlugin_logic_chunksLogic_0_hitCalc_HIT;
      fetch_logic_ctrls_2_up_BtbPlugin_logic_chunksLogic_1_readRsp_ENTRY_hash <= fetch_logic_ctrls_1_down_BtbPlugin_logic_chunksLogic_1_readRsp_ENTRY_hash;
      fetch_logic_ctrls_2_up_BtbPlugin_logic_chunksLogic_1_readRsp_ENTRY_sliceLow <= fetch_logic_ctrls_1_down_BtbPlugin_logic_chunksLogic_1_readRsp_ENTRY_sliceLow;
      fetch_logic_ctrls_2_up_BtbPlugin_logic_chunksLogic_1_readRsp_ENTRY_pcTarget <= fetch_logic_ctrls_1_down_BtbPlugin_logic_chunksLogic_1_readRsp_ENTRY_pcTarget;
      fetch_logic_ctrls_2_up_BtbPlugin_logic_chunksLogic_1_readRsp_ENTRY_isBranch <= fetch_logic_ctrls_1_down_BtbPlugin_logic_chunksLogic_1_readRsp_ENTRY_isBranch;
      fetch_logic_ctrls_2_up_BtbPlugin_logic_chunksLogic_1_readRsp_ENTRY_isPush <= fetch_logic_ctrls_1_down_BtbPlugin_logic_chunksLogic_1_readRsp_ENTRY_isPush;
      fetch_logic_ctrls_2_up_BtbPlugin_logic_chunksLogic_1_readRsp_ENTRY_isPop <= fetch_logic_ctrls_1_down_BtbPlugin_logic_chunksLogic_1_readRsp_ENTRY_isPop;
      fetch_logic_ctrls_2_up_BtbPlugin_logic_chunksLogic_1_hitCalc_HIT <= fetch_logic_ctrls_1_down_BtbPlugin_logic_chunksLogic_1_hitCalc_HIT;
      fetch_logic_ctrls_2_up_MMU_HAZARD <= fetch_logic_ctrls_1_down_MMU_HAZARD;
      fetch_logic_ctrls_2_up_MMU_REFILL <= fetch_logic_ctrls_1_down_MMU_REFILL;
      fetch_logic_ctrls_2_up_MMU_TRANSLATED <= fetch_logic_ctrls_1_down_MMU_TRANSLATED;
      fetch_logic_ctrls_2_up_MMU_ALLOW_EXECUTE <= fetch_logic_ctrls_1_down_MMU_ALLOW_EXECUTE;
      fetch_logic_ctrls_2_up_MMU_PAGE_FAULT <= fetch_logic_ctrls_1_down_MMU_PAGE_FAULT;
      fetch_logic_ctrls_2_up_MMU_ACCESS_FAULT <= fetch_logic_ctrls_1_down_MMU_ACCESS_FAULT;
    end
    if(toplevel_decode_ctrls_0_down_isReady) begin
      toplevel_decode_ctrls_1_up_Decode_INSTRUCTION_0 <= toplevel_decode_ctrls_0_down_Decode_INSTRUCTION_0;
      toplevel_decode_ctrls_1_up_Decode_DECOMPRESSION_FAULT_0 <= toplevel_decode_ctrls_0_down_Decode_DECOMPRESSION_FAULT_0;
      toplevel_decode_ctrls_1_up_Decode_INSTRUCTION_RAW_0 <= toplevel_decode_ctrls_0_down_Decode_INSTRUCTION_RAW_0;
      toplevel_decode_ctrls_1_up_Decode_INSTRUCTION_SLICE_COUNT_0 <= toplevel_decode_ctrls_0_down_Decode_INSTRUCTION_SLICE_COUNT_0;
      toplevel_decode_ctrls_1_up_PC_0 <= toplevel_decode_ctrls_0_down_PC_0;
      toplevel_decode_ctrls_1_up_Decode_DOP_ID_0 <= toplevel_decode_ctrls_0_down_Decode_DOP_ID_0;
      toplevel_decode_ctrls_1_up_GSharePlugin_GSHARE_COUNTER_0_0 <= toplevel_decode_ctrls_0_down_GSharePlugin_GSHARE_COUNTER_0_0;
      toplevel_decode_ctrls_1_up_GSharePlugin_GSHARE_COUNTER_0_1 <= toplevel_decode_ctrls_0_down_GSharePlugin_GSHARE_COUNTER_0_1;
      toplevel_decode_ctrls_1_up_GSharePlugin_GSHARE_COUNTER_0_2 <= toplevel_decode_ctrls_0_down_GSharePlugin_GSHARE_COUNTER_0_2;
      toplevel_decode_ctrls_1_up_GSharePlugin_GSHARE_COUNTER_0_3 <= toplevel_decode_ctrls_0_down_GSharePlugin_GSHARE_COUNTER_0_3;
      toplevel_decode_ctrls_1_up_Prediction_BRANCH_HISTORY_0 <= toplevel_decode_ctrls_0_down_Prediction_BRANCH_HISTORY_0;
      toplevel_decode_ctrls_1_up_TRAP_0 <= toplevel_decode_ctrls_0_down_TRAP_0;
      toplevel_decode_ctrls_1_up_Prediction_ALIGNED_JUMPED_0 <= toplevel_decode_ctrls_0_down_Prediction_ALIGNED_JUMPED_0;
      toplevel_decode_ctrls_1_up_Prediction_ALIGNED_JUMPED_PC_0 <= toplevel_decode_ctrls_0_down_Prediction_ALIGNED_JUMPED_PC_0;
      toplevel_decode_ctrls_1_up_Prediction_ALIGNED_SLICES_BRANCH_0 <= toplevel_decode_ctrls_0_down_Prediction_ALIGNED_SLICES_BRANCH_0;
      toplevel_decode_ctrls_1_up_Prediction_ALIGNED_SLICES_TAKEN_0 <= toplevel_decode_ctrls_0_down_Prediction_ALIGNED_SLICES_TAKEN_0;
      toplevel_decode_ctrls_1_up_Prediction_ALIGN_REDO_0 <= toplevel_decode_ctrls_0_down_Prediction_ALIGN_REDO_0;
      toplevel_decode_ctrls_1_up_Decode_INSTRUCTION_1 <= toplevel_decode_ctrls_0_down_Decode_INSTRUCTION_1;
      toplevel_decode_ctrls_1_up_Decode_DECOMPRESSION_FAULT_1 <= toplevel_decode_ctrls_0_down_Decode_DECOMPRESSION_FAULT_1;
      toplevel_decode_ctrls_1_up_Decode_INSTRUCTION_RAW_1 <= toplevel_decode_ctrls_0_down_Decode_INSTRUCTION_RAW_1;
      toplevel_decode_ctrls_1_up_Decode_INSTRUCTION_SLICE_COUNT_1 <= toplevel_decode_ctrls_0_down_Decode_INSTRUCTION_SLICE_COUNT_1;
      toplevel_decode_ctrls_1_up_PC_1 <= toplevel_decode_ctrls_0_down_PC_1;
      toplevel_decode_ctrls_1_up_Decode_DOP_ID_1 <= toplevel_decode_ctrls_0_down_Decode_DOP_ID_1;
      toplevel_decode_ctrls_1_up_GSharePlugin_GSHARE_COUNTER_1_0 <= toplevel_decode_ctrls_0_down_GSharePlugin_GSHARE_COUNTER_1_0;
      toplevel_decode_ctrls_1_up_GSharePlugin_GSHARE_COUNTER_1_1 <= toplevel_decode_ctrls_0_down_GSharePlugin_GSHARE_COUNTER_1_1;
      toplevel_decode_ctrls_1_up_GSharePlugin_GSHARE_COUNTER_1_2 <= toplevel_decode_ctrls_0_down_GSharePlugin_GSHARE_COUNTER_1_2;
      toplevel_decode_ctrls_1_up_GSharePlugin_GSHARE_COUNTER_1_3 <= toplevel_decode_ctrls_0_down_GSharePlugin_GSHARE_COUNTER_1_3;
      toplevel_decode_ctrls_1_up_Prediction_BRANCH_HISTORY_1 <= toplevel_decode_ctrls_0_down_Prediction_BRANCH_HISTORY_1;
      toplevel_decode_ctrls_1_up_TRAP_1 <= toplevel_decode_ctrls_0_down_TRAP_1;
      toplevel_decode_ctrls_1_up_Prediction_ALIGNED_JUMPED_1 <= toplevel_decode_ctrls_0_down_Prediction_ALIGNED_JUMPED_1;
      toplevel_decode_ctrls_1_up_Prediction_ALIGNED_JUMPED_PC_1 <= toplevel_decode_ctrls_0_down_Prediction_ALIGNED_JUMPED_PC_1;
      toplevel_decode_ctrls_1_up_Prediction_ALIGNED_SLICES_BRANCH_1 <= toplevel_decode_ctrls_0_down_Prediction_ALIGNED_SLICES_BRANCH_1;
      toplevel_decode_ctrls_1_up_Prediction_ALIGNED_SLICES_TAKEN_1 <= toplevel_decode_ctrls_0_down_Prediction_ALIGNED_SLICES_TAKEN_1;
      toplevel_decode_ctrls_1_up_Prediction_ALIGN_REDO_1 <= toplevel_decode_ctrls_0_down_Prediction_ALIGN_REDO_1;
    end
    if(toplevel_execute_ctrl0_down_isReady) begin
      toplevel_execute_ctrl1_up_Decode_UOP_lane0 <= toplevel_execute_ctrl0_down_Decode_UOP_lane0;
      toplevel_execute_ctrl1_up_Prediction_ALIGNED_JUMPED_lane0 <= toplevel_execute_ctrl0_down_Prediction_ALIGNED_JUMPED_lane0;
      toplevel_execute_ctrl1_up_Prediction_ALIGNED_JUMPED_PC_lane0 <= toplevel_execute_ctrl0_down_Prediction_ALIGNED_JUMPED_PC_lane0;
      toplevel_execute_ctrl1_up_Prediction_ALIGNED_SLICES_TAKEN_lane0 <= toplevel_execute_ctrl0_down_Prediction_ALIGNED_SLICES_TAKEN_lane0;
      toplevel_execute_ctrl1_up_Prediction_ALIGNED_SLICES_BRANCH_lane0 <= toplevel_execute_ctrl0_down_Prediction_ALIGNED_SLICES_BRANCH_lane0;
      toplevel_execute_ctrl1_up_GSharePlugin_GSHARE_COUNTER_lane0_0 <= toplevel_execute_ctrl0_down_GSharePlugin_GSHARE_COUNTER_lane0_0;
      toplevel_execute_ctrl1_up_GSharePlugin_GSHARE_COUNTER_lane0_1 <= toplevel_execute_ctrl0_down_GSharePlugin_GSHARE_COUNTER_lane0_1;
      toplevel_execute_ctrl1_up_GSharePlugin_GSHARE_COUNTER_lane0_2 <= toplevel_execute_ctrl0_down_GSharePlugin_GSHARE_COUNTER_lane0_2;
      toplevel_execute_ctrl1_up_GSharePlugin_GSHARE_COUNTER_lane0_3 <= toplevel_execute_ctrl0_down_GSharePlugin_GSHARE_COUNTER_lane0_3;
      toplevel_execute_ctrl1_up_Prediction_BRANCH_HISTORY_lane0 <= toplevel_execute_ctrl0_down_Prediction_BRANCH_HISTORY_lane0;
      toplevel_execute_ctrl1_up_Decode_INSTRUCTION_SLICE_COUNT_lane0 <= toplevel_execute_ctrl0_down_Decode_INSTRUCTION_SLICE_COUNT_lane0;
      toplevel_execute_ctrl1_up_PC_lane0 <= toplevel_execute_ctrl0_down_PC_lane0;
      toplevel_execute_ctrl1_up_TRAP_lane0 <= toplevel_execute_ctrl0_down_TRAP_lane0;
      toplevel_execute_ctrl1_up_Decode_UOP_ID_lane0 <= toplevel_execute_ctrl0_down_Decode_UOP_ID_lane0;
      toplevel_execute_ctrl1_up_RS1_PHYS_lane0 <= toplevel_execute_ctrl0_down_RS1_PHYS_lane0;
      toplevel_execute_ctrl1_up_RS2_PHYS_lane0 <= toplevel_execute_ctrl0_down_RS2_PHYS_lane0;
      toplevel_execute_ctrl1_up_RD_ENABLE_lane0 <= toplevel_execute_ctrl0_down_RD_ENABLE_lane0;
      toplevel_execute_ctrl1_up_RD_PHYS_lane0 <= toplevel_execute_ctrl0_down_RD_PHYS_lane0;
      toplevel_execute_ctrl1_up_LANE_AGE_lane0 <= toplevel_execute_ctrl0_down_LANE_AGE_lane0;
      toplevel_execute_ctrl1_up_COMPLETED_lane0 <= toplevel_execute_ctrl0_down_COMPLETED_lane0;
      toplevel_execute_ctrl1_up_execute_lane0_LAYER_SEL_lane0 <= toplevel_execute_ctrl0_down_execute_lane0_LAYER_SEL_lane0;
      toplevel_execute_ctrl1_up_Decode_UOP_lane1 <= toplevel_execute_ctrl0_down_Decode_UOP_lane1;
      toplevel_execute_ctrl1_up_Prediction_ALIGNED_JUMPED_lane1 <= toplevel_execute_ctrl0_down_Prediction_ALIGNED_JUMPED_lane1;
      toplevel_execute_ctrl1_up_Prediction_ALIGNED_JUMPED_PC_lane1 <= toplevel_execute_ctrl0_down_Prediction_ALIGNED_JUMPED_PC_lane1;
      toplevel_execute_ctrl1_up_Prediction_ALIGNED_SLICES_TAKEN_lane1 <= toplevel_execute_ctrl0_down_Prediction_ALIGNED_SLICES_TAKEN_lane1;
      toplevel_execute_ctrl1_up_Prediction_ALIGNED_SLICES_BRANCH_lane1 <= toplevel_execute_ctrl0_down_Prediction_ALIGNED_SLICES_BRANCH_lane1;
      toplevel_execute_ctrl1_up_GSharePlugin_GSHARE_COUNTER_lane1_0 <= toplevel_execute_ctrl0_down_GSharePlugin_GSHARE_COUNTER_lane1_0;
      toplevel_execute_ctrl1_up_GSharePlugin_GSHARE_COUNTER_lane1_1 <= toplevel_execute_ctrl0_down_GSharePlugin_GSHARE_COUNTER_lane1_1;
      toplevel_execute_ctrl1_up_GSharePlugin_GSHARE_COUNTER_lane1_2 <= toplevel_execute_ctrl0_down_GSharePlugin_GSHARE_COUNTER_lane1_2;
      toplevel_execute_ctrl1_up_GSharePlugin_GSHARE_COUNTER_lane1_3 <= toplevel_execute_ctrl0_down_GSharePlugin_GSHARE_COUNTER_lane1_3;
      toplevel_execute_ctrl1_up_Prediction_BRANCH_HISTORY_lane1 <= toplevel_execute_ctrl0_down_Prediction_BRANCH_HISTORY_lane1;
      toplevel_execute_ctrl1_up_Decode_INSTRUCTION_SLICE_COUNT_lane1 <= toplevel_execute_ctrl0_down_Decode_INSTRUCTION_SLICE_COUNT_lane1;
      toplevel_execute_ctrl1_up_PC_lane1 <= toplevel_execute_ctrl0_down_PC_lane1;
      toplevel_execute_ctrl1_up_TRAP_lane1 <= toplevel_execute_ctrl0_down_TRAP_lane1;
      toplevel_execute_ctrl1_up_Decode_UOP_ID_lane1 <= toplevel_execute_ctrl0_down_Decode_UOP_ID_lane1;
      toplevel_execute_ctrl1_up_RS1_PHYS_lane1 <= toplevel_execute_ctrl0_down_RS1_PHYS_lane1;
      toplevel_execute_ctrl1_up_RS2_PHYS_lane1 <= toplevel_execute_ctrl0_down_RS2_PHYS_lane1;
      toplevel_execute_ctrl1_up_RD_ENABLE_lane1 <= toplevel_execute_ctrl0_down_RD_ENABLE_lane1;
      toplevel_execute_ctrl1_up_RD_PHYS_lane1 <= toplevel_execute_ctrl0_down_RD_PHYS_lane1;
      toplevel_execute_ctrl1_up_LANE_AGE_lane1 <= toplevel_execute_ctrl0_down_LANE_AGE_lane1;
      toplevel_execute_ctrl1_up_COMPLETED_lane1 <= toplevel_execute_ctrl0_down_COMPLETED_lane1;
      toplevel_execute_ctrl1_up_execute_lane1_LAYER_SEL_lane1 <= toplevel_execute_ctrl0_down_execute_lane1_LAYER_SEL_lane1;
      toplevel_execute_ctrl1_up_AguPlugin_SIZE_lane0 <= toplevel_execute_ctrl0_down_AguPlugin_SIZE_lane0;
    end
    if(toplevel_execute_ctrl1_down_isReady) begin
      toplevel_execute_ctrl2_up_Decode_UOP_lane0 <= toplevel_execute_ctrl1_down_Decode_UOP_lane0;
      toplevel_execute_ctrl2_up_Prediction_ALIGNED_JUMPED_lane0 <= toplevel_execute_ctrl1_down_Prediction_ALIGNED_JUMPED_lane0;
      toplevel_execute_ctrl2_up_Prediction_ALIGNED_JUMPED_PC_lane0 <= toplevel_execute_ctrl1_down_Prediction_ALIGNED_JUMPED_PC_lane0;
      toplevel_execute_ctrl2_up_Prediction_ALIGNED_SLICES_TAKEN_lane0 <= toplevel_execute_ctrl1_down_Prediction_ALIGNED_SLICES_TAKEN_lane0;
      toplevel_execute_ctrl2_up_Prediction_ALIGNED_SLICES_BRANCH_lane0 <= toplevel_execute_ctrl1_down_Prediction_ALIGNED_SLICES_BRANCH_lane0;
      toplevel_execute_ctrl2_up_GSharePlugin_GSHARE_COUNTER_lane0_0 <= toplevel_execute_ctrl1_down_GSharePlugin_GSHARE_COUNTER_lane0_0;
      toplevel_execute_ctrl2_up_GSharePlugin_GSHARE_COUNTER_lane0_1 <= toplevel_execute_ctrl1_down_GSharePlugin_GSHARE_COUNTER_lane0_1;
      toplevel_execute_ctrl2_up_GSharePlugin_GSHARE_COUNTER_lane0_2 <= toplevel_execute_ctrl1_down_GSharePlugin_GSHARE_COUNTER_lane0_2;
      toplevel_execute_ctrl2_up_GSharePlugin_GSHARE_COUNTER_lane0_3 <= toplevel_execute_ctrl1_down_GSharePlugin_GSHARE_COUNTER_lane0_3;
      toplevel_execute_ctrl2_up_Prediction_BRANCH_HISTORY_lane0 <= toplevel_execute_ctrl1_down_Prediction_BRANCH_HISTORY_lane0;
      toplevel_execute_ctrl2_up_Decode_INSTRUCTION_SLICE_COUNT_lane0 <= toplevel_execute_ctrl1_down_Decode_INSTRUCTION_SLICE_COUNT_lane0;
      toplevel_execute_ctrl2_up_PC_lane0 <= toplevel_execute_ctrl1_down_PC_lane0;
      toplevel_execute_ctrl2_up_TRAP_lane0 <= toplevel_execute_ctrl1_down_TRAP_lane0;
      toplevel_execute_ctrl2_up_Decode_UOP_ID_lane0 <= toplevel_execute_ctrl1_down_Decode_UOP_ID_lane0;
      toplevel_execute_ctrl2_up_RS1_PHYS_lane0 <= toplevel_execute_ctrl1_down_RS1_PHYS_lane0;
      toplevel_execute_ctrl2_up_RS2_PHYS_lane0 <= toplevel_execute_ctrl1_down_RS2_PHYS_lane0;
      toplevel_execute_ctrl2_up_RD_ENABLE_lane0 <= toplevel_execute_ctrl1_down_RD_ENABLE_lane0;
      toplevel_execute_ctrl2_up_RD_PHYS_lane0 <= toplevel_execute_ctrl1_down_RD_PHYS_lane0;
      toplevel_execute_ctrl2_up_LANE_AGE_lane0 <= toplevel_execute_ctrl1_down_LANE_AGE_lane0;
      toplevel_execute_ctrl2_up_COMPLETED_lane0 <= toplevel_execute_ctrl1_down_COMPLETED_lane0;
      toplevel_execute_ctrl2_up_Decode_UOP_lane1 <= toplevel_execute_ctrl1_down_Decode_UOP_lane1;
      toplevel_execute_ctrl2_up_Prediction_ALIGNED_JUMPED_lane1 <= toplevel_execute_ctrl1_down_Prediction_ALIGNED_JUMPED_lane1;
      toplevel_execute_ctrl2_up_Prediction_ALIGNED_JUMPED_PC_lane1 <= toplevel_execute_ctrl1_down_Prediction_ALIGNED_JUMPED_PC_lane1;
      toplevel_execute_ctrl2_up_Prediction_ALIGNED_SLICES_TAKEN_lane1 <= toplevel_execute_ctrl1_down_Prediction_ALIGNED_SLICES_TAKEN_lane1;
      toplevel_execute_ctrl2_up_Prediction_ALIGNED_SLICES_BRANCH_lane1 <= toplevel_execute_ctrl1_down_Prediction_ALIGNED_SLICES_BRANCH_lane1;
      toplevel_execute_ctrl2_up_GSharePlugin_GSHARE_COUNTER_lane1_0 <= toplevel_execute_ctrl1_down_GSharePlugin_GSHARE_COUNTER_lane1_0;
      toplevel_execute_ctrl2_up_GSharePlugin_GSHARE_COUNTER_lane1_1 <= toplevel_execute_ctrl1_down_GSharePlugin_GSHARE_COUNTER_lane1_1;
      toplevel_execute_ctrl2_up_GSharePlugin_GSHARE_COUNTER_lane1_2 <= toplevel_execute_ctrl1_down_GSharePlugin_GSHARE_COUNTER_lane1_2;
      toplevel_execute_ctrl2_up_GSharePlugin_GSHARE_COUNTER_lane1_3 <= toplevel_execute_ctrl1_down_GSharePlugin_GSHARE_COUNTER_lane1_3;
      toplevel_execute_ctrl2_up_Prediction_BRANCH_HISTORY_lane1 <= toplevel_execute_ctrl1_down_Prediction_BRANCH_HISTORY_lane1;
      toplevel_execute_ctrl2_up_Decode_INSTRUCTION_SLICE_COUNT_lane1 <= toplevel_execute_ctrl1_down_Decode_INSTRUCTION_SLICE_COUNT_lane1;
      toplevel_execute_ctrl2_up_PC_lane1 <= toplevel_execute_ctrl1_down_PC_lane1;
      toplevel_execute_ctrl2_up_TRAP_lane1 <= toplevel_execute_ctrl1_down_TRAP_lane1;
      toplevel_execute_ctrl2_up_Decode_UOP_ID_lane1 <= toplevel_execute_ctrl1_down_Decode_UOP_ID_lane1;
      toplevel_execute_ctrl2_up_RS1_PHYS_lane1 <= toplevel_execute_ctrl1_down_RS1_PHYS_lane1;
      toplevel_execute_ctrl2_up_RS2_PHYS_lane1 <= toplevel_execute_ctrl1_down_RS2_PHYS_lane1;
      toplevel_execute_ctrl2_up_RD_ENABLE_lane1 <= toplevel_execute_ctrl1_down_RD_ENABLE_lane1;
      toplevel_execute_ctrl2_up_RD_PHYS_lane1 <= toplevel_execute_ctrl1_down_RD_PHYS_lane1;
      toplevel_execute_ctrl2_up_LANE_AGE_lane1 <= toplevel_execute_ctrl1_down_LANE_AGE_lane1;
      toplevel_execute_ctrl2_up_COMPLETED_lane1 <= toplevel_execute_ctrl1_down_COMPLETED_lane1;
      toplevel_execute_ctrl2_up_AguPlugin_SIZE_lane0 <= toplevel_execute_ctrl1_down_AguPlugin_SIZE_lane0;
      toplevel_execute_ctrl2_up_early0_SrcPlugin_SRC1_lane0 <= toplevel_execute_ctrl1_down_early0_SrcPlugin_SRC1_lane0;
      toplevel_execute_ctrl2_up_integer_RS1_lane0 <= toplevel_execute_ctrl1_down_integer_RS1_lane0;
      toplevel_execute_ctrl2_up_early0_SrcPlugin_SRC2_lane0 <= toplevel_execute_ctrl1_down_early0_SrcPlugin_SRC2_lane0;
      toplevel_execute_ctrl2_up_integer_RS2_lane0 <= toplevel_execute_ctrl1_down_integer_RS2_lane0;
      toplevel_execute_ctrl2_up_early1_SrcPlugin_SRC1_lane1 <= toplevel_execute_ctrl1_down_early1_SrcPlugin_SRC1_lane1;
      toplevel_execute_ctrl2_up_integer_RS1_lane1 <= toplevel_execute_ctrl1_down_integer_RS1_lane1;
      toplevel_execute_ctrl2_up_early1_SrcPlugin_SRC2_lane1 <= toplevel_execute_ctrl1_down_early1_SrcPlugin_SRC2_lane1;
      toplevel_execute_ctrl2_up_integer_RS2_lane1 <= toplevel_execute_ctrl1_down_integer_RS2_lane1;
      toplevel_execute_ctrl2_up_MAY_FLUSH_PRECISE_3_lane0 <= toplevel_execute_ctrl1_down_MAY_FLUSH_PRECISE_3_lane0;
      toplevel_execute_ctrl2_up_MAY_FLUSH_PRECISE_3_lane1 <= toplevel_execute_ctrl1_down_MAY_FLUSH_PRECISE_3_lane1;
      toplevel_execute_ctrl2_up_early0_IntAluPlugin_SEL_lane0 <= toplevel_execute_ctrl1_down_early0_IntAluPlugin_SEL_lane0;
      toplevel_execute_ctrl2_up_early0_BarrelShifterPlugin_SEL_lane0 <= toplevel_execute_ctrl1_down_early0_BarrelShifterPlugin_SEL_lane0;
      toplevel_execute_ctrl2_up_early0_BranchPlugin_SEL_lane0 <= toplevel_execute_ctrl1_down_early0_BranchPlugin_SEL_lane0;
      toplevel_execute_ctrl2_up_early0_MulPlugin_SEL_lane0 <= toplevel_execute_ctrl1_down_early0_MulPlugin_SEL_lane0;
      toplevel_execute_ctrl2_up_early0_DivPlugin_SEL_lane0 <= toplevel_execute_ctrl1_down_early0_DivPlugin_SEL_lane0;
      toplevel_execute_ctrl2_up_early0_EnvPlugin_SEL_lane0 <= toplevel_execute_ctrl1_down_early0_EnvPlugin_SEL_lane0;
      toplevel_execute_ctrl2_up_late0_IntAluPlugin_SEL_lane0 <= toplevel_execute_ctrl1_down_late0_IntAluPlugin_SEL_lane0;
      toplevel_execute_ctrl2_up_late0_BarrelShifterPlugin_SEL_lane0 <= toplevel_execute_ctrl1_down_late0_BarrelShifterPlugin_SEL_lane0;
      toplevel_execute_ctrl2_up_late0_BranchPlugin_SEL_lane0 <= toplevel_execute_ctrl1_down_late0_BranchPlugin_SEL_lane0;
      toplevel_execute_ctrl2_up_MulPlugin_HIGH_lane0 <= toplevel_execute_ctrl1_down_MulPlugin_HIGH_lane0;
      toplevel_execute_ctrl2_up_CsrAccessPlugin_SEL_lane0 <= toplevel_execute_ctrl1_down_CsrAccessPlugin_SEL_lane0;
      toplevel_execute_ctrl2_up_AguPlugin_SEL_lane0 <= toplevel_execute_ctrl1_down_AguPlugin_SEL_lane0;
      toplevel_execute_ctrl2_up_LsuPlugin_logic_FENCE_lane0 <= toplevel_execute_ctrl1_down_LsuPlugin_logic_FENCE_lane0;
      toplevel_execute_ctrl2_up_lane0_integer_WriteBackPlugin_SEL_lane0 <= toplevel_execute_ctrl1_down_lane0_integer_WriteBackPlugin_SEL_lane0;
      toplevel_execute_ctrl2_up_COMPLETION_AT_2_lane0 <= toplevel_execute_ctrl1_down_COMPLETION_AT_2_lane0;
      toplevel_execute_ctrl2_up_COMPLETION_AT_3_lane0 <= toplevel_execute_ctrl1_down_COMPLETION_AT_3_lane0;
      toplevel_execute_ctrl2_up_COMPLETION_AT_4_lane0 <= toplevel_execute_ctrl1_down_COMPLETION_AT_4_lane0;
      toplevel_execute_ctrl2_up_execute_lane0_logic_completions_onCtrl_0_ENABLE_lane0 <= toplevel_execute_ctrl1_down_execute_lane0_logic_completions_onCtrl_0_ENABLE_lane0;
      toplevel_execute_ctrl2_up_execute_lane0_logic_completions_onCtrl_1_ENABLE_lane0 <= toplevel_execute_ctrl1_down_execute_lane0_logic_completions_onCtrl_1_ENABLE_lane0;
      toplevel_execute_ctrl2_up_execute_lane0_logic_completions_onCtrl_2_ENABLE_lane0 <= toplevel_execute_ctrl1_down_execute_lane0_logic_completions_onCtrl_2_ENABLE_lane0;
      toplevel_execute_ctrl2_up_early0_IntAluPlugin_ALU_ADD_SUB_lane0 <= toplevel_execute_ctrl1_down_early0_IntAluPlugin_ALU_ADD_SUB_lane0;
      toplevel_execute_ctrl2_up_early0_IntAluPlugin_ALU_SLTX_lane0 <= toplevel_execute_ctrl1_down_early0_IntAluPlugin_ALU_SLTX_lane0;
      toplevel_execute_ctrl2_up_early0_IntAluPlugin_ALU_BITWISE_CTRL_lane0 <= toplevel_execute_ctrl1_down_early0_IntAluPlugin_ALU_BITWISE_CTRL_lane0;
      toplevel_execute_ctrl2_up_SrcStageables_REVERT_lane0 <= toplevel_execute_ctrl1_down_SrcStageables_REVERT_lane0;
      toplevel_execute_ctrl2_up_SrcStageables_ZERO_lane0 <= toplevel_execute_ctrl1_down_SrcStageables_ZERO_lane0;
      toplevel_execute_ctrl2_up_lane0_IntFormatPlugin_logic_SIGNED_lane0 <= toplevel_execute_ctrl1_down_lane0_IntFormatPlugin_logic_SIGNED_lane0;
      toplevel_execute_ctrl2_up_lane0_IntFormatPlugin_logic_WIDTH_ID_lane0 <= toplevel_execute_ctrl1_down_lane0_IntFormatPlugin_logic_WIDTH_ID_lane0;
      toplevel_execute_ctrl2_up_BYPASSED_AT_3_lane0 <= toplevel_execute_ctrl1_down_BYPASSED_AT_3_lane0;
      toplevel_execute_ctrl2_up_SrcStageables_UNSIGNED_lane0 <= toplevel_execute_ctrl1_down_SrcStageables_UNSIGNED_lane0;
      toplevel_execute_ctrl2_up_BarrelShifterPlugin_LEFT_lane0 <= toplevel_execute_ctrl1_down_BarrelShifterPlugin_LEFT_lane0;
      toplevel_execute_ctrl2_up_BarrelShifterPlugin_SIGNED_lane0 <= toplevel_execute_ctrl1_down_BarrelShifterPlugin_SIGNED_lane0;
      toplevel_execute_ctrl2_up_BranchPlugin_BRANCH_CTRL_lane0 <= toplevel_execute_ctrl1_down_BranchPlugin_BRANCH_CTRL_lane0;
      toplevel_execute_ctrl2_up_RsUnsignedPlugin_RS1_SIGNED_lane0 <= toplevel_execute_ctrl1_down_RsUnsignedPlugin_RS1_SIGNED_lane0;
      toplevel_execute_ctrl2_up_RsUnsignedPlugin_RS2_SIGNED_lane0 <= toplevel_execute_ctrl1_down_RsUnsignedPlugin_RS2_SIGNED_lane0;
      toplevel_execute_ctrl2_up_DivPlugin_REM_lane0 <= toplevel_execute_ctrl1_down_DivPlugin_REM_lane0;
      toplevel_execute_ctrl2_up_CsrAccessPlugin_CSR_IMM_lane0 <= toplevel_execute_ctrl1_down_CsrAccessPlugin_CSR_IMM_lane0;
      toplevel_execute_ctrl2_up_CsrAccessPlugin_CSR_MASK_lane0 <= toplevel_execute_ctrl1_down_CsrAccessPlugin_CSR_MASK_lane0;
      toplevel_execute_ctrl2_up_CsrAccessPlugin_CSR_CLEAR_lane0 <= toplevel_execute_ctrl1_down_CsrAccessPlugin_CSR_CLEAR_lane0;
      toplevel_execute_ctrl2_up_AguPlugin_LOAD_lane0 <= toplevel_execute_ctrl1_down_AguPlugin_LOAD_lane0;
      toplevel_execute_ctrl2_up_AguPlugin_STORE_lane0 <= toplevel_execute_ctrl1_down_AguPlugin_STORE_lane0;
      toplevel_execute_ctrl2_up_AguPlugin_ATOMIC_lane0 <= toplevel_execute_ctrl1_down_AguPlugin_ATOMIC_lane0;
      toplevel_execute_ctrl2_up_AguPlugin_FLOAT_lane0 <= toplevel_execute_ctrl1_down_AguPlugin_FLOAT_lane0;
      toplevel_execute_ctrl2_up_LsuPlugin_logic_LSU_PREFETCH_lane0 <= toplevel_execute_ctrl1_down_LsuPlugin_logic_LSU_PREFETCH_lane0;
      toplevel_execute_ctrl2_up_early0_EnvPlugin_OP_lane0 <= toplevel_execute_ctrl1_down_early0_EnvPlugin_OP_lane0;
      toplevel_execute_ctrl2_up_late0_IntAluPlugin_ALU_ADD_SUB_lane0 <= toplevel_execute_ctrl1_down_late0_IntAluPlugin_ALU_ADD_SUB_lane0;
      toplevel_execute_ctrl2_up_late0_IntAluPlugin_ALU_SLTX_lane0 <= toplevel_execute_ctrl1_down_late0_IntAluPlugin_ALU_SLTX_lane0;
      toplevel_execute_ctrl2_up_late0_IntAluPlugin_ALU_BITWISE_CTRL_lane0 <= toplevel_execute_ctrl1_down_late0_IntAluPlugin_ALU_BITWISE_CTRL_lane0;
      toplevel_execute_ctrl2_up_late0_SrcPlugin_logic_SRC1_CTRL_lane0 <= toplevel_execute_ctrl1_down_late0_SrcPlugin_logic_SRC1_CTRL_lane0;
      toplevel_execute_ctrl2_up_late0_SrcPlugin_logic_SRC2_CTRL_lane0 <= toplevel_execute_ctrl1_down_late0_SrcPlugin_logic_SRC2_CTRL_lane0;
      toplevel_execute_ctrl2_up_early1_IntAluPlugin_SEL_lane1 <= toplevel_execute_ctrl1_down_early1_IntAluPlugin_SEL_lane1;
      toplevel_execute_ctrl2_up_early1_BarrelShifterPlugin_SEL_lane1 <= toplevel_execute_ctrl1_down_early1_BarrelShifterPlugin_SEL_lane1;
      toplevel_execute_ctrl2_up_early1_BranchPlugin_SEL_lane1 <= toplevel_execute_ctrl1_down_early1_BranchPlugin_SEL_lane1;
      toplevel_execute_ctrl2_up_late1_IntAluPlugin_SEL_lane1 <= toplevel_execute_ctrl1_down_late1_IntAluPlugin_SEL_lane1;
      toplevel_execute_ctrl2_up_late1_BarrelShifterPlugin_SEL_lane1 <= toplevel_execute_ctrl1_down_late1_BarrelShifterPlugin_SEL_lane1;
      toplevel_execute_ctrl2_up_late1_BranchPlugin_SEL_lane1 <= toplevel_execute_ctrl1_down_late1_BranchPlugin_SEL_lane1;
      toplevel_execute_ctrl2_up_lane1_integer_WriteBackPlugin_SEL_lane1 <= toplevel_execute_ctrl1_down_lane1_integer_WriteBackPlugin_SEL_lane1;
      toplevel_execute_ctrl2_up_COMPLETION_AT_2_lane1 <= toplevel_execute_ctrl1_down_COMPLETION_AT_2_lane1;
      toplevel_execute_ctrl2_up_COMPLETION_AT_3_lane1 <= toplevel_execute_ctrl1_down_COMPLETION_AT_3_lane1;
      toplevel_execute_ctrl2_up_COMPLETION_AT_4_lane1 <= toplevel_execute_ctrl1_down_COMPLETION_AT_4_lane1;
      toplevel_execute_ctrl2_up_execute_lane1_logic_completions_onCtrl_0_ENABLE_lane1 <= toplevel_execute_ctrl1_down_execute_lane1_logic_completions_onCtrl_0_ENABLE_lane1;
      toplevel_execute_ctrl2_up_execute_lane1_logic_completions_onCtrl_1_ENABLE_lane1 <= toplevel_execute_ctrl1_down_execute_lane1_logic_completions_onCtrl_1_ENABLE_lane1;
      toplevel_execute_ctrl2_up_execute_lane1_logic_completions_onCtrl_2_ENABLE_lane1 <= toplevel_execute_ctrl1_down_execute_lane1_logic_completions_onCtrl_2_ENABLE_lane1;
      toplevel_execute_ctrl2_up_early1_IntAluPlugin_ALU_ADD_SUB_lane1 <= toplevel_execute_ctrl1_down_early1_IntAluPlugin_ALU_ADD_SUB_lane1;
      toplevel_execute_ctrl2_up_early1_IntAluPlugin_ALU_SLTX_lane1 <= toplevel_execute_ctrl1_down_early1_IntAluPlugin_ALU_SLTX_lane1;
      toplevel_execute_ctrl2_up_early1_IntAluPlugin_ALU_BITWISE_CTRL_lane1 <= toplevel_execute_ctrl1_down_early1_IntAluPlugin_ALU_BITWISE_CTRL_lane1;
      toplevel_execute_ctrl2_up_SrcStageables_REVERT_lane1 <= toplevel_execute_ctrl1_down_SrcStageables_REVERT_lane1;
      toplevel_execute_ctrl2_up_SrcStageables_ZERO_lane1 <= toplevel_execute_ctrl1_down_SrcStageables_ZERO_lane1;
      toplevel_execute_ctrl2_up_BYPASSED_AT_3_lane1 <= toplevel_execute_ctrl1_down_BYPASSED_AT_3_lane1;
      toplevel_execute_ctrl2_up_SrcStageables_UNSIGNED_lane1 <= toplevel_execute_ctrl1_down_SrcStageables_UNSIGNED_lane1;
      toplevel_execute_ctrl2_up_BarrelShifterPlugin_LEFT_lane1 <= toplevel_execute_ctrl1_down_BarrelShifterPlugin_LEFT_lane1;
      toplevel_execute_ctrl2_up_BarrelShifterPlugin_SIGNED_lane1 <= toplevel_execute_ctrl1_down_BarrelShifterPlugin_SIGNED_lane1;
      toplevel_execute_ctrl2_up_BranchPlugin_BRANCH_CTRL_lane1 <= toplevel_execute_ctrl1_down_BranchPlugin_BRANCH_CTRL_lane1;
      toplevel_execute_ctrl2_up_late1_IntAluPlugin_ALU_ADD_SUB_lane1 <= toplevel_execute_ctrl1_down_late1_IntAluPlugin_ALU_ADD_SUB_lane1;
      toplevel_execute_ctrl2_up_late1_IntAluPlugin_ALU_SLTX_lane1 <= toplevel_execute_ctrl1_down_late1_IntAluPlugin_ALU_SLTX_lane1;
      toplevel_execute_ctrl2_up_late1_IntAluPlugin_ALU_BITWISE_CTRL_lane1 <= toplevel_execute_ctrl1_down_late1_IntAluPlugin_ALU_BITWISE_CTRL_lane1;
      toplevel_execute_ctrl2_up_late1_SrcPlugin_logic_SRC1_CTRL_lane1 <= toplevel_execute_ctrl1_down_late1_SrcPlugin_logic_SRC1_CTRL_lane1;
      toplevel_execute_ctrl2_up_late1_SrcPlugin_logic_SRC2_CTRL_lane1 <= toplevel_execute_ctrl1_down_late1_SrcPlugin_logic_SRC2_CTRL_lane1;
    end
    if(toplevel_execute_ctrl2_down_isReady) begin
      toplevel_execute_ctrl3_up_Decode_UOP_lane0 <= toplevel_execute_ctrl2_down_Decode_UOP_lane0;
      toplevel_execute_ctrl3_up_Prediction_ALIGNED_JUMPED_lane0 <= toplevel_execute_ctrl2_down_Prediction_ALIGNED_JUMPED_lane0;
      toplevel_execute_ctrl3_up_Prediction_ALIGNED_JUMPED_PC_lane0 <= toplevel_execute_ctrl2_down_Prediction_ALIGNED_JUMPED_PC_lane0;
      toplevel_execute_ctrl3_up_Prediction_ALIGNED_SLICES_TAKEN_lane0 <= toplevel_execute_ctrl2_down_Prediction_ALIGNED_SLICES_TAKEN_lane0;
      toplevel_execute_ctrl3_up_Prediction_ALIGNED_SLICES_BRANCH_lane0 <= toplevel_execute_ctrl2_down_Prediction_ALIGNED_SLICES_BRANCH_lane0;
      toplevel_execute_ctrl3_up_GSharePlugin_GSHARE_COUNTER_lane0_0 <= toplevel_execute_ctrl2_down_GSharePlugin_GSHARE_COUNTER_lane0_0;
      toplevel_execute_ctrl3_up_GSharePlugin_GSHARE_COUNTER_lane0_1 <= toplevel_execute_ctrl2_down_GSharePlugin_GSHARE_COUNTER_lane0_1;
      toplevel_execute_ctrl3_up_GSharePlugin_GSHARE_COUNTER_lane0_2 <= toplevel_execute_ctrl2_down_GSharePlugin_GSHARE_COUNTER_lane0_2;
      toplevel_execute_ctrl3_up_GSharePlugin_GSHARE_COUNTER_lane0_3 <= toplevel_execute_ctrl2_down_GSharePlugin_GSHARE_COUNTER_lane0_3;
      toplevel_execute_ctrl3_up_Prediction_BRANCH_HISTORY_lane0 <= toplevel_execute_ctrl2_down_Prediction_BRANCH_HISTORY_lane0;
      toplevel_execute_ctrl3_up_Decode_INSTRUCTION_SLICE_COUNT_lane0 <= toplevel_execute_ctrl2_down_Decode_INSTRUCTION_SLICE_COUNT_lane0;
      toplevel_execute_ctrl3_up_PC_lane0 <= toplevel_execute_ctrl2_down_PC_lane0;
      toplevel_execute_ctrl3_up_TRAP_lane0 <= toplevel_execute_ctrl2_down_TRAP_lane0;
      toplevel_execute_ctrl3_up_Decode_UOP_ID_lane0 <= toplevel_execute_ctrl2_down_Decode_UOP_ID_lane0;
      toplevel_execute_ctrl3_up_RS1_PHYS_lane0 <= toplevel_execute_ctrl2_down_RS1_PHYS_lane0;
      toplevel_execute_ctrl3_up_RS2_PHYS_lane0 <= toplevel_execute_ctrl2_down_RS2_PHYS_lane0;
      toplevel_execute_ctrl3_up_RD_ENABLE_lane0 <= toplevel_execute_ctrl2_down_RD_ENABLE_lane0;
      toplevel_execute_ctrl3_up_RD_PHYS_lane0 <= toplevel_execute_ctrl2_down_RD_PHYS_lane0;
      toplevel_execute_ctrl3_up_LANE_AGE_lane0 <= toplevel_execute_ctrl2_down_LANE_AGE_lane0;
      toplevel_execute_ctrl3_up_COMPLETED_lane0 <= toplevel_execute_ctrl2_down_COMPLETED_lane0;
      toplevel_execute_ctrl3_up_Decode_UOP_lane1 <= toplevel_execute_ctrl2_down_Decode_UOP_lane1;
      toplevel_execute_ctrl3_up_Prediction_ALIGNED_JUMPED_lane1 <= toplevel_execute_ctrl2_down_Prediction_ALIGNED_JUMPED_lane1;
      toplevel_execute_ctrl3_up_Prediction_ALIGNED_JUMPED_PC_lane1 <= toplevel_execute_ctrl2_down_Prediction_ALIGNED_JUMPED_PC_lane1;
      toplevel_execute_ctrl3_up_Prediction_ALIGNED_SLICES_TAKEN_lane1 <= toplevel_execute_ctrl2_down_Prediction_ALIGNED_SLICES_TAKEN_lane1;
      toplevel_execute_ctrl3_up_Prediction_ALIGNED_SLICES_BRANCH_lane1 <= toplevel_execute_ctrl2_down_Prediction_ALIGNED_SLICES_BRANCH_lane1;
      toplevel_execute_ctrl3_up_GSharePlugin_GSHARE_COUNTER_lane1_0 <= toplevel_execute_ctrl2_down_GSharePlugin_GSHARE_COUNTER_lane1_0;
      toplevel_execute_ctrl3_up_GSharePlugin_GSHARE_COUNTER_lane1_1 <= toplevel_execute_ctrl2_down_GSharePlugin_GSHARE_COUNTER_lane1_1;
      toplevel_execute_ctrl3_up_GSharePlugin_GSHARE_COUNTER_lane1_2 <= toplevel_execute_ctrl2_down_GSharePlugin_GSHARE_COUNTER_lane1_2;
      toplevel_execute_ctrl3_up_GSharePlugin_GSHARE_COUNTER_lane1_3 <= toplevel_execute_ctrl2_down_GSharePlugin_GSHARE_COUNTER_lane1_3;
      toplevel_execute_ctrl3_up_Prediction_BRANCH_HISTORY_lane1 <= toplevel_execute_ctrl2_down_Prediction_BRANCH_HISTORY_lane1;
      toplevel_execute_ctrl3_up_Decode_INSTRUCTION_SLICE_COUNT_lane1 <= toplevel_execute_ctrl2_down_Decode_INSTRUCTION_SLICE_COUNT_lane1;
      toplevel_execute_ctrl3_up_PC_lane1 <= toplevel_execute_ctrl2_down_PC_lane1;
      toplevel_execute_ctrl3_up_TRAP_lane1 <= toplevel_execute_ctrl2_down_TRAP_lane1;
      toplevel_execute_ctrl3_up_Decode_UOP_ID_lane1 <= toplevel_execute_ctrl2_down_Decode_UOP_ID_lane1;
      toplevel_execute_ctrl3_up_RS1_PHYS_lane1 <= toplevel_execute_ctrl2_down_RS1_PHYS_lane1;
      toplevel_execute_ctrl3_up_RS2_PHYS_lane1 <= toplevel_execute_ctrl2_down_RS2_PHYS_lane1;
      toplevel_execute_ctrl3_up_RD_ENABLE_lane1 <= toplevel_execute_ctrl2_down_RD_ENABLE_lane1;
      toplevel_execute_ctrl3_up_RD_PHYS_lane1 <= toplevel_execute_ctrl2_down_RD_PHYS_lane1;
      toplevel_execute_ctrl3_up_LANE_AGE_lane1 <= toplevel_execute_ctrl2_down_LANE_AGE_lane1;
      toplevel_execute_ctrl3_up_COMPLETED_lane1 <= toplevel_execute_ctrl2_down_COMPLETED_lane1;
      toplevel_execute_ctrl3_up_AguPlugin_SIZE_lane0 <= toplevel_execute_ctrl2_down_AguPlugin_SIZE_lane0;
      toplevel_execute_ctrl3_up_integer_RS1_lane0 <= toplevel_execute_ctrl2_down_integer_RS1_lane0;
      toplevel_execute_ctrl3_up_integer_RS2_lane0 <= toplevel_execute_ctrl2_down_integer_RS2_lane0;
      toplevel_execute_ctrl3_up_integer_RS1_lane1 <= toplevel_execute_ctrl2_down_integer_RS1_lane1;
      toplevel_execute_ctrl3_up_integer_RS2_lane1 <= toplevel_execute_ctrl2_down_integer_RS2_lane1;
      toplevel_execute_ctrl3_up_early0_BarrelShifterPlugin_SEL_lane0 <= toplevel_execute_ctrl2_down_early0_BarrelShifterPlugin_SEL_lane0;
      toplevel_execute_ctrl3_up_early0_BranchPlugin_SEL_lane0 <= toplevel_execute_ctrl2_down_early0_BranchPlugin_SEL_lane0;
      toplevel_execute_ctrl3_up_early0_MulPlugin_SEL_lane0 <= toplevel_execute_ctrl2_down_early0_MulPlugin_SEL_lane0;
      toplevel_execute_ctrl3_up_early0_DivPlugin_SEL_lane0 <= toplevel_execute_ctrl2_down_early0_DivPlugin_SEL_lane0;
      toplevel_execute_ctrl3_up_late0_IntAluPlugin_SEL_lane0 <= toplevel_execute_ctrl2_down_late0_IntAluPlugin_SEL_lane0;
      toplevel_execute_ctrl3_up_late0_BarrelShifterPlugin_SEL_lane0 <= toplevel_execute_ctrl2_down_late0_BarrelShifterPlugin_SEL_lane0;
      toplevel_execute_ctrl3_up_late0_BranchPlugin_SEL_lane0 <= toplevel_execute_ctrl2_down_late0_BranchPlugin_SEL_lane0;
      toplevel_execute_ctrl3_up_MulPlugin_HIGH_lane0 <= toplevel_execute_ctrl2_down_MulPlugin_HIGH_lane0;
      toplevel_execute_ctrl3_up_CsrAccessPlugin_SEL_lane0 <= toplevel_execute_ctrl2_down_CsrAccessPlugin_SEL_lane0;
      toplevel_execute_ctrl3_up_AguPlugin_SEL_lane0 <= toplevel_execute_ctrl2_down_AguPlugin_SEL_lane0;
      toplevel_execute_ctrl3_up_LsuPlugin_logic_FENCE_lane0 <= toplevel_execute_ctrl2_down_LsuPlugin_logic_FENCE_lane0;
      toplevel_execute_ctrl3_up_lane0_integer_WriteBackPlugin_SEL_lane0 <= toplevel_execute_ctrl2_down_lane0_integer_WriteBackPlugin_SEL_lane0;
      toplevel_execute_ctrl3_up_COMPLETION_AT_3_lane0 <= toplevel_execute_ctrl2_down_COMPLETION_AT_3_lane0;
      toplevel_execute_ctrl3_up_COMPLETION_AT_4_lane0 <= toplevel_execute_ctrl2_down_COMPLETION_AT_4_lane0;
      toplevel_execute_ctrl3_up_execute_lane0_logic_completions_onCtrl_1_ENABLE_lane0 <= toplevel_execute_ctrl2_down_execute_lane0_logic_completions_onCtrl_1_ENABLE_lane0;
      toplevel_execute_ctrl3_up_execute_lane0_logic_completions_onCtrl_2_ENABLE_lane0 <= toplevel_execute_ctrl2_down_execute_lane0_logic_completions_onCtrl_2_ENABLE_lane0;
      toplevel_execute_ctrl3_up_SrcStageables_REVERT_lane0 <= toplevel_execute_ctrl2_down_SrcStageables_REVERT_lane0;
      toplevel_execute_ctrl3_up_SrcStageables_ZERO_lane0 <= toplevel_execute_ctrl2_down_SrcStageables_ZERO_lane0;
      toplevel_execute_ctrl3_up_lane0_IntFormatPlugin_logic_SIGNED_lane0 <= toplevel_execute_ctrl2_down_lane0_IntFormatPlugin_logic_SIGNED_lane0;
      toplevel_execute_ctrl3_up_lane0_IntFormatPlugin_logic_WIDTH_ID_lane0 <= toplevel_execute_ctrl2_down_lane0_IntFormatPlugin_logic_WIDTH_ID_lane0;
      toplevel_execute_ctrl3_up_SrcStageables_UNSIGNED_lane0 <= toplevel_execute_ctrl2_down_SrcStageables_UNSIGNED_lane0;
      toplevel_execute_ctrl3_up_BarrelShifterPlugin_LEFT_lane0 <= toplevel_execute_ctrl2_down_BarrelShifterPlugin_LEFT_lane0;
      toplevel_execute_ctrl3_up_BarrelShifterPlugin_SIGNED_lane0 <= toplevel_execute_ctrl2_down_BarrelShifterPlugin_SIGNED_lane0;
      toplevel_execute_ctrl3_up_BranchPlugin_BRANCH_CTRL_lane0 <= toplevel_execute_ctrl2_down_BranchPlugin_BRANCH_CTRL_lane0;
      toplevel_execute_ctrl3_up_AguPlugin_LOAD_lane0 <= toplevel_execute_ctrl2_down_AguPlugin_LOAD_lane0;
      toplevel_execute_ctrl3_up_AguPlugin_STORE_lane0 <= toplevel_execute_ctrl2_down_AguPlugin_STORE_lane0;
      toplevel_execute_ctrl3_up_AguPlugin_ATOMIC_lane0 <= toplevel_execute_ctrl2_down_AguPlugin_ATOMIC_lane0;
      toplevel_execute_ctrl3_up_AguPlugin_FLOAT_lane0 <= toplevel_execute_ctrl2_down_AguPlugin_FLOAT_lane0;
      toplevel_execute_ctrl3_up_LsuPlugin_logic_LSU_PREFETCH_lane0 <= toplevel_execute_ctrl2_down_LsuPlugin_logic_LSU_PREFETCH_lane0;
      toplevel_execute_ctrl3_up_late0_IntAluPlugin_ALU_ADD_SUB_lane0 <= toplevel_execute_ctrl2_down_late0_IntAluPlugin_ALU_ADD_SUB_lane0;
      toplevel_execute_ctrl3_up_late0_IntAluPlugin_ALU_SLTX_lane0 <= toplevel_execute_ctrl2_down_late0_IntAluPlugin_ALU_SLTX_lane0;
      toplevel_execute_ctrl3_up_late0_IntAluPlugin_ALU_BITWISE_CTRL_lane0 <= toplevel_execute_ctrl2_down_late0_IntAluPlugin_ALU_BITWISE_CTRL_lane0;
      toplevel_execute_ctrl3_up_late0_SrcPlugin_logic_SRC1_CTRL_lane0 <= toplevel_execute_ctrl2_down_late0_SrcPlugin_logic_SRC1_CTRL_lane0;
      toplevel_execute_ctrl3_up_late0_SrcPlugin_logic_SRC2_CTRL_lane0 <= toplevel_execute_ctrl2_down_late0_SrcPlugin_logic_SRC2_CTRL_lane0;
      toplevel_execute_ctrl3_up_early1_BarrelShifterPlugin_SEL_lane1 <= toplevel_execute_ctrl2_down_early1_BarrelShifterPlugin_SEL_lane1;
      toplevel_execute_ctrl3_up_early1_BranchPlugin_SEL_lane1 <= toplevel_execute_ctrl2_down_early1_BranchPlugin_SEL_lane1;
      toplevel_execute_ctrl3_up_late1_IntAluPlugin_SEL_lane1 <= toplevel_execute_ctrl2_down_late1_IntAluPlugin_SEL_lane1;
      toplevel_execute_ctrl3_up_late1_BarrelShifterPlugin_SEL_lane1 <= toplevel_execute_ctrl2_down_late1_BarrelShifterPlugin_SEL_lane1;
      toplevel_execute_ctrl3_up_late1_BranchPlugin_SEL_lane1 <= toplevel_execute_ctrl2_down_late1_BranchPlugin_SEL_lane1;
      toplevel_execute_ctrl3_up_lane1_integer_WriteBackPlugin_SEL_lane1 <= toplevel_execute_ctrl2_down_lane1_integer_WriteBackPlugin_SEL_lane1;
      toplevel_execute_ctrl3_up_COMPLETION_AT_3_lane1 <= toplevel_execute_ctrl2_down_COMPLETION_AT_3_lane1;
      toplevel_execute_ctrl3_up_COMPLETION_AT_4_lane1 <= toplevel_execute_ctrl2_down_COMPLETION_AT_4_lane1;
      toplevel_execute_ctrl3_up_execute_lane1_logic_completions_onCtrl_1_ENABLE_lane1 <= toplevel_execute_ctrl2_down_execute_lane1_logic_completions_onCtrl_1_ENABLE_lane1;
      toplevel_execute_ctrl3_up_execute_lane1_logic_completions_onCtrl_2_ENABLE_lane1 <= toplevel_execute_ctrl2_down_execute_lane1_logic_completions_onCtrl_2_ENABLE_lane1;
      toplevel_execute_ctrl3_up_SrcStageables_REVERT_lane1 <= toplevel_execute_ctrl2_down_SrcStageables_REVERT_lane1;
      toplevel_execute_ctrl3_up_SrcStageables_ZERO_lane1 <= toplevel_execute_ctrl2_down_SrcStageables_ZERO_lane1;
      toplevel_execute_ctrl3_up_SrcStageables_UNSIGNED_lane1 <= toplevel_execute_ctrl2_down_SrcStageables_UNSIGNED_lane1;
      toplevel_execute_ctrl3_up_BarrelShifterPlugin_LEFT_lane1 <= toplevel_execute_ctrl2_down_BarrelShifterPlugin_LEFT_lane1;
      toplevel_execute_ctrl3_up_BarrelShifterPlugin_SIGNED_lane1 <= toplevel_execute_ctrl2_down_BarrelShifterPlugin_SIGNED_lane1;
      toplevel_execute_ctrl3_up_BranchPlugin_BRANCH_CTRL_lane1 <= toplevel_execute_ctrl2_down_BranchPlugin_BRANCH_CTRL_lane1;
      toplevel_execute_ctrl3_up_late1_IntAluPlugin_ALU_ADD_SUB_lane1 <= toplevel_execute_ctrl2_down_late1_IntAluPlugin_ALU_ADD_SUB_lane1;
      toplevel_execute_ctrl3_up_late1_IntAluPlugin_ALU_SLTX_lane1 <= toplevel_execute_ctrl2_down_late1_IntAluPlugin_ALU_SLTX_lane1;
      toplevel_execute_ctrl3_up_late1_IntAluPlugin_ALU_BITWISE_CTRL_lane1 <= toplevel_execute_ctrl2_down_late1_IntAluPlugin_ALU_BITWISE_CTRL_lane1;
      toplevel_execute_ctrl3_up_late1_SrcPlugin_logic_SRC1_CTRL_lane1 <= toplevel_execute_ctrl2_down_late1_SrcPlugin_logic_SRC1_CTRL_lane1;
      toplevel_execute_ctrl3_up_late1_SrcPlugin_logic_SRC2_CTRL_lane1 <= toplevel_execute_ctrl2_down_late1_SrcPlugin_logic_SRC2_CTRL_lane1;
      toplevel_execute_ctrl3_up_COMMIT_lane0 <= toplevel_execute_ctrl2_down_COMMIT_lane0;
      toplevel_execute_ctrl3_up_COMMIT_lane1 <= toplevel_execute_ctrl2_down_COMMIT_lane1;
      toplevel_execute_ctrl3_up_early0_SrcPlugin_ADD_SUB_lane0 <= toplevel_execute_ctrl2_down_early0_SrcPlugin_ADD_SUB_lane0;
      toplevel_execute_ctrl3_up_early0_SrcPlugin_LESS_lane0 <= toplevel_execute_ctrl2_down_early0_SrcPlugin_LESS_lane0;
      toplevel_execute_ctrl3_up_early0_BarrelShifterPlugin_SHIFT_RESULT_lane0 <= toplevel_execute_ctrl2_down_early0_BarrelShifterPlugin_SHIFT_RESULT_lane0;
      toplevel_execute_ctrl3_up_MUL_SRC1_lane0 <= toplevel_execute_ctrl2_down_MUL_SRC1_lane0;
      toplevel_execute_ctrl3_up_MUL_SRC2_lane0 <= toplevel_execute_ctrl2_down_MUL_SRC2_lane0;
      toplevel_execute_ctrl3_up_DivPlugin_DIV_RESULT_lane0 <= toplevel_execute_ctrl2_down_DivPlugin_DIV_RESULT_lane0;
      toplevel_execute_ctrl3_up_early1_SrcPlugin_LESS_lane1 <= toplevel_execute_ctrl2_down_early1_SrcPlugin_LESS_lane1;
      toplevel_execute_ctrl3_up_early1_BarrelShifterPlugin_SHIFT_RESULT_lane1 <= toplevel_execute_ctrl2_down_early1_BarrelShifterPlugin_SHIFT_RESULT_lane1;
      toplevel_execute_ctrl3_up_early0_BranchPlugin_pcCalc_PC_TRUE_lane0 <= toplevel_execute_ctrl2_down_early0_BranchPlugin_pcCalc_PC_TRUE_lane0;
      toplevel_execute_ctrl3_up_early0_BranchPlugin_pcCalc_PC_FALSE_lane0 <= toplevel_execute_ctrl2_down_early0_BranchPlugin_pcCalc_PC_FALSE_lane0;
      toplevel_execute_ctrl3_up_early0_BranchPlugin_pcCalc_PC_LAST_SLICE_lane0 <= toplevel_execute_ctrl2_down_early0_BranchPlugin_pcCalc_PC_LAST_SLICE_lane0;
      toplevel_execute_ctrl3_up_early1_BranchPlugin_pcCalc_PC_TRUE_lane1 <= toplevel_execute_ctrl2_down_early1_BranchPlugin_pcCalc_PC_TRUE_lane1;
      toplevel_execute_ctrl3_up_early1_BranchPlugin_pcCalc_PC_FALSE_lane1 <= toplevel_execute_ctrl2_down_early1_BranchPlugin_pcCalc_PC_FALSE_lane1;
      toplevel_execute_ctrl3_up_early1_BranchPlugin_pcCalc_PC_LAST_SLICE_lane1 <= toplevel_execute_ctrl2_down_early1_BranchPlugin_pcCalc_PC_LAST_SLICE_lane1;
      toplevel_execute_ctrl3_up_early0_BranchPlugin_logic_alu_EQ_lane0 <= toplevel_execute_ctrl2_down_early0_BranchPlugin_logic_alu_EQ_lane0;
      toplevel_execute_ctrl3_up_early0_BranchPlugin_logic_alu_btb_BAD_TARGET_lane0 <= toplevel_execute_ctrl2_down_early0_BranchPlugin_logic_alu_btb_BAD_TARGET_lane0;
      toplevel_execute_ctrl3_up_early0_BranchPlugin_logic_alu_MSB_FAILED_lane0 <= toplevel_execute_ctrl2_down_early0_BranchPlugin_logic_alu_MSB_FAILED_lane0;
      toplevel_execute_ctrl3_up_early1_BranchPlugin_logic_alu_EQ_lane1 <= toplevel_execute_ctrl2_down_early1_BranchPlugin_logic_alu_EQ_lane1;
      toplevel_execute_ctrl3_up_early1_BranchPlugin_logic_alu_btb_BAD_TARGET_lane1 <= toplevel_execute_ctrl2_down_early1_BranchPlugin_logic_alu_btb_BAD_TARGET_lane1;
      toplevel_execute_ctrl3_up_early1_BranchPlugin_logic_alu_MSB_FAILED_lane1 <= toplevel_execute_ctrl2_down_early1_BranchPlugin_logic_alu_MSB_FAILED_lane1;
      toplevel_execute_ctrl3_up_lane0_integer_WriteBackPlugin_logic_DATA_lane0 <= toplevel_execute_ctrl2_down_lane0_integer_WriteBackPlugin_logic_DATA_lane0;
      toplevel_execute_ctrl3_up_lane1_integer_WriteBackPlugin_logic_DATA_lane1 <= toplevel_execute_ctrl2_down_lane1_integer_WriteBackPlugin_logic_DATA_lane1;
      toplevel_execute_ctrl3_up_LsuL1_MIXED_ADDRESS_lane0 <= toplevel_execute_ctrl2_down_LsuL1_MIXED_ADDRESS_lane0;
      toplevel_execute_ctrl3_up_LsuL1Plugin_logic_BANK_BUSY_lane0 <= toplevel_execute_ctrl2_down_LsuL1Plugin_logic_BANK_BUSY_lane0;
      toplevel_execute_ctrl3_up_LsuL1Plugin_logic_EVENT_WRITE_VALID_lane0 <= toplevel_execute_ctrl2_down_LsuL1Plugin_logic_EVENT_WRITE_VALID_lane0;
      toplevel_execute_ctrl3_up_LsuL1Plugin_logic_EVENT_WRITE_ADDRESS_lane0 <= toplevel_execute_ctrl2_down_LsuL1Plugin_logic_EVENT_WRITE_ADDRESS_lane0;
      toplevel_execute_ctrl3_up_LsuL1Plugin_logic_ls_rt0_SHARED_BYPASS_VALID_lane0 <= toplevel_execute_ctrl2_down_LsuL1Plugin_logic_ls_rt0_SHARED_BYPASS_VALID_lane0;
      toplevel_execute_ctrl3_up_LsuL1Plugin_logic_ls_rt0_SHARED_BYPASS_VALUE_lane0_plru_0 <= toplevel_execute_ctrl2_down_LsuL1Plugin_logic_ls_rt0_SHARED_BYPASS_VALUE_lane0_plru_0;
      toplevel_execute_ctrl3_up_LsuL1Plugin_logic_ls_rt0_SHARED_BYPASS_VALUE_lane0_dirty <= toplevel_execute_ctrl2_down_LsuL1Plugin_logic_ls_rt0_SHARED_BYPASS_VALUE_lane0_dirty;
      toplevel_execute_ctrl3_up_LsuL1Plugin_logic_EVENT_WRITE_DATA_lane0 <= toplevel_execute_ctrl2_down_LsuL1Plugin_logic_EVENT_WRITE_DATA_lane0;
      toplevel_execute_ctrl3_up_LsuL1Plugin_logic_EVENT_WRITE_MASK_lane0 <= toplevel_execute_ctrl2_down_LsuL1Plugin_logic_EVENT_WRITE_MASK_lane0;
      toplevel_execute_ctrl3_up_LsuPlugin_logic_FORCE_PHYSICAL_lane0 <= toplevel_execute_ctrl2_down_LsuPlugin_logic_FORCE_PHYSICAL_lane0;
      toplevel_execute_ctrl3_up_LsuPlugin_logic_FROM_ACCESS_lane0 <= toplevel_execute_ctrl2_down_LsuPlugin_logic_FROM_ACCESS_lane0;
      toplevel_execute_ctrl3_up_LsuL1_MASK_lane0 <= toplevel_execute_ctrl2_down_LsuL1_MASK_lane0;
      toplevel_execute_ctrl3_up_LsuL1_SIZE_lane0 <= toplevel_execute_ctrl2_down_LsuL1_SIZE_lane0;
      toplevel_execute_ctrl3_up_LsuL1_LOAD_lane0 <= toplevel_execute_ctrl2_down_LsuL1_LOAD_lane0;
      toplevel_execute_ctrl3_up_LsuL1_ATOMIC_lane0 <= toplevel_execute_ctrl2_down_LsuL1_ATOMIC_lane0;
      toplevel_execute_ctrl3_up_LsuL1_STORE_lane0 <= toplevel_execute_ctrl2_down_LsuL1_STORE_lane0;
      toplevel_execute_ctrl3_up_LsuL1_PREFETCH_lane0 <= toplevel_execute_ctrl2_down_LsuL1_PREFETCH_lane0;
      toplevel_execute_ctrl3_up_LsuL1_FLUSH_lane0 <= toplevel_execute_ctrl2_down_LsuL1_FLUSH_lane0;
      toplevel_execute_ctrl3_up_Decode_STORE_ID_lane0 <= toplevel_execute_ctrl2_down_Decode_STORE_ID_lane0;
      toplevel_execute_ctrl3_up_LsuPlugin_logic_FROM_LSU_lane0 <= toplevel_execute_ctrl2_down_LsuPlugin_logic_FROM_LSU_lane0;
      toplevel_execute_ctrl3_up_LsuPlugin_logic_FROM_PREFETCH_lane0 <= toplevel_execute_ctrl2_down_LsuPlugin_logic_FROM_PREFETCH_lane0;
    end
    if(toplevel_execute_ctrl3_down_isReady) begin
      toplevel_execute_ctrl4_up_Decode_UOP_lane0 <= toplevel_execute_ctrl3_down_Decode_UOP_lane0;
      toplevel_execute_ctrl4_up_Prediction_ALIGNED_JUMPED_lane0 <= toplevel_execute_ctrl3_down_Prediction_ALIGNED_JUMPED_lane0;
      toplevel_execute_ctrl4_up_Prediction_ALIGNED_JUMPED_PC_lane0 <= toplevel_execute_ctrl3_down_Prediction_ALIGNED_JUMPED_PC_lane0;
      toplevel_execute_ctrl4_up_Prediction_ALIGNED_SLICES_TAKEN_lane0 <= toplevel_execute_ctrl3_down_Prediction_ALIGNED_SLICES_TAKEN_lane0;
      toplevel_execute_ctrl4_up_Prediction_ALIGNED_SLICES_BRANCH_lane0 <= toplevel_execute_ctrl3_down_Prediction_ALIGNED_SLICES_BRANCH_lane0;
      toplevel_execute_ctrl4_up_GSharePlugin_GSHARE_COUNTER_lane0_0 <= toplevel_execute_ctrl3_down_GSharePlugin_GSHARE_COUNTER_lane0_0;
      toplevel_execute_ctrl4_up_GSharePlugin_GSHARE_COUNTER_lane0_1 <= toplevel_execute_ctrl3_down_GSharePlugin_GSHARE_COUNTER_lane0_1;
      toplevel_execute_ctrl4_up_GSharePlugin_GSHARE_COUNTER_lane0_2 <= toplevel_execute_ctrl3_down_GSharePlugin_GSHARE_COUNTER_lane0_2;
      toplevel_execute_ctrl4_up_GSharePlugin_GSHARE_COUNTER_lane0_3 <= toplevel_execute_ctrl3_down_GSharePlugin_GSHARE_COUNTER_lane0_3;
      toplevel_execute_ctrl4_up_Prediction_BRANCH_HISTORY_lane0 <= toplevel_execute_ctrl3_down_Prediction_BRANCH_HISTORY_lane0;
      toplevel_execute_ctrl4_up_Decode_INSTRUCTION_SLICE_COUNT_lane0 <= toplevel_execute_ctrl3_down_Decode_INSTRUCTION_SLICE_COUNT_lane0;
      toplevel_execute_ctrl4_up_PC_lane0 <= toplevel_execute_ctrl3_down_PC_lane0;
      toplevel_execute_ctrl4_up_TRAP_lane0 <= toplevel_execute_ctrl3_down_TRAP_lane0;
      toplevel_execute_ctrl4_up_Decode_UOP_ID_lane0 <= toplevel_execute_ctrl3_down_Decode_UOP_ID_lane0;
      toplevel_execute_ctrl4_up_RD_ENABLE_lane0 <= toplevel_execute_ctrl3_down_RD_ENABLE_lane0;
      toplevel_execute_ctrl4_up_RD_PHYS_lane0 <= toplevel_execute_ctrl3_down_RD_PHYS_lane0;
      toplevel_execute_ctrl4_up_LANE_AGE_lane0 <= toplevel_execute_ctrl3_down_LANE_AGE_lane0;
      toplevel_execute_ctrl4_up_COMPLETED_lane0 <= toplevel_execute_ctrl3_down_COMPLETED_lane0;
      toplevel_execute_ctrl4_up_Decode_UOP_lane1 <= toplevel_execute_ctrl3_down_Decode_UOP_lane1;
      toplevel_execute_ctrl4_up_Prediction_ALIGNED_JUMPED_lane1 <= toplevel_execute_ctrl3_down_Prediction_ALIGNED_JUMPED_lane1;
      toplevel_execute_ctrl4_up_Prediction_ALIGNED_JUMPED_PC_lane1 <= toplevel_execute_ctrl3_down_Prediction_ALIGNED_JUMPED_PC_lane1;
      toplevel_execute_ctrl4_up_Prediction_ALIGNED_SLICES_TAKEN_lane1 <= toplevel_execute_ctrl3_down_Prediction_ALIGNED_SLICES_TAKEN_lane1;
      toplevel_execute_ctrl4_up_Prediction_ALIGNED_SLICES_BRANCH_lane1 <= toplevel_execute_ctrl3_down_Prediction_ALIGNED_SLICES_BRANCH_lane1;
      toplevel_execute_ctrl4_up_GSharePlugin_GSHARE_COUNTER_lane1_0 <= toplevel_execute_ctrl3_down_GSharePlugin_GSHARE_COUNTER_lane1_0;
      toplevel_execute_ctrl4_up_GSharePlugin_GSHARE_COUNTER_lane1_1 <= toplevel_execute_ctrl3_down_GSharePlugin_GSHARE_COUNTER_lane1_1;
      toplevel_execute_ctrl4_up_GSharePlugin_GSHARE_COUNTER_lane1_2 <= toplevel_execute_ctrl3_down_GSharePlugin_GSHARE_COUNTER_lane1_2;
      toplevel_execute_ctrl4_up_GSharePlugin_GSHARE_COUNTER_lane1_3 <= toplevel_execute_ctrl3_down_GSharePlugin_GSHARE_COUNTER_lane1_3;
      toplevel_execute_ctrl4_up_Prediction_BRANCH_HISTORY_lane1 <= toplevel_execute_ctrl3_down_Prediction_BRANCH_HISTORY_lane1;
      toplevel_execute_ctrl4_up_Decode_INSTRUCTION_SLICE_COUNT_lane1 <= toplevel_execute_ctrl3_down_Decode_INSTRUCTION_SLICE_COUNT_lane1;
      toplevel_execute_ctrl4_up_PC_lane1 <= toplevel_execute_ctrl3_down_PC_lane1;
      toplevel_execute_ctrl4_up_TRAP_lane1 <= toplevel_execute_ctrl3_down_TRAP_lane1;
      toplevel_execute_ctrl4_up_Decode_UOP_ID_lane1 <= toplevel_execute_ctrl3_down_Decode_UOP_ID_lane1;
      toplevel_execute_ctrl4_up_RD_ENABLE_lane1 <= toplevel_execute_ctrl3_down_RD_ENABLE_lane1;
      toplevel_execute_ctrl4_up_RD_PHYS_lane1 <= toplevel_execute_ctrl3_down_RD_PHYS_lane1;
      toplevel_execute_ctrl4_up_LANE_AGE_lane1 <= toplevel_execute_ctrl3_down_LANE_AGE_lane1;
      toplevel_execute_ctrl4_up_COMPLETED_lane1 <= toplevel_execute_ctrl3_down_COMPLETED_lane1;
      toplevel_execute_ctrl4_up_AguPlugin_SIZE_lane0 <= toplevel_execute_ctrl3_down_AguPlugin_SIZE_lane0;
      toplevel_execute_ctrl4_up_integer_RS2_lane0 <= toplevel_execute_ctrl3_down_integer_RS2_lane0;
      toplevel_execute_ctrl4_up_early0_BranchPlugin_SEL_lane0 <= toplevel_execute_ctrl3_down_early0_BranchPlugin_SEL_lane0;
      toplevel_execute_ctrl4_up_early0_MulPlugin_SEL_lane0 <= toplevel_execute_ctrl3_down_early0_MulPlugin_SEL_lane0;
      toplevel_execute_ctrl4_up_late0_IntAluPlugin_SEL_lane0 <= toplevel_execute_ctrl3_down_late0_IntAluPlugin_SEL_lane0;
      toplevel_execute_ctrl4_up_late0_BarrelShifterPlugin_SEL_lane0 <= toplevel_execute_ctrl3_down_late0_BarrelShifterPlugin_SEL_lane0;
      toplevel_execute_ctrl4_up_late0_BranchPlugin_SEL_lane0 <= toplevel_execute_ctrl3_down_late0_BranchPlugin_SEL_lane0;
      toplevel_execute_ctrl4_up_MulPlugin_HIGH_lane0 <= toplevel_execute_ctrl3_down_MulPlugin_HIGH_lane0;
      toplevel_execute_ctrl4_up_AguPlugin_SEL_lane0 <= toplevel_execute_ctrl3_down_AguPlugin_SEL_lane0;
      toplevel_execute_ctrl4_up_LsuPlugin_logic_FENCE_lane0 <= toplevel_execute_ctrl3_down_LsuPlugin_logic_FENCE_lane0;
      toplevel_execute_ctrl4_up_lane0_integer_WriteBackPlugin_SEL_lane0 <= toplevel_execute_ctrl3_down_lane0_integer_WriteBackPlugin_SEL_lane0;
      toplevel_execute_ctrl4_up_COMPLETION_AT_4_lane0 <= toplevel_execute_ctrl3_down_COMPLETION_AT_4_lane0;
      toplevel_execute_ctrl4_up_execute_lane0_logic_completions_onCtrl_2_ENABLE_lane0 <= toplevel_execute_ctrl3_down_execute_lane0_logic_completions_onCtrl_2_ENABLE_lane0;
      toplevel_execute_ctrl4_up_SrcStageables_REVERT_lane0 <= toplevel_execute_ctrl3_down_SrcStageables_REVERT_lane0;
      toplevel_execute_ctrl4_up_SrcStageables_ZERO_lane0 <= toplevel_execute_ctrl3_down_SrcStageables_ZERO_lane0;
      toplevel_execute_ctrl4_up_lane0_IntFormatPlugin_logic_SIGNED_lane0 <= toplevel_execute_ctrl3_down_lane0_IntFormatPlugin_logic_SIGNED_lane0;
      toplevel_execute_ctrl4_up_lane0_IntFormatPlugin_logic_WIDTH_ID_lane0 <= toplevel_execute_ctrl3_down_lane0_IntFormatPlugin_logic_WIDTH_ID_lane0;
      toplevel_execute_ctrl4_up_SrcStageables_UNSIGNED_lane0 <= toplevel_execute_ctrl3_down_SrcStageables_UNSIGNED_lane0;
      toplevel_execute_ctrl4_up_BarrelShifterPlugin_LEFT_lane0 <= toplevel_execute_ctrl3_down_BarrelShifterPlugin_LEFT_lane0;
      toplevel_execute_ctrl4_up_BarrelShifterPlugin_SIGNED_lane0 <= toplevel_execute_ctrl3_down_BarrelShifterPlugin_SIGNED_lane0;
      toplevel_execute_ctrl4_up_BranchPlugin_BRANCH_CTRL_lane0 <= toplevel_execute_ctrl3_down_BranchPlugin_BRANCH_CTRL_lane0;
      toplevel_execute_ctrl4_up_AguPlugin_LOAD_lane0 <= toplevel_execute_ctrl3_down_AguPlugin_LOAD_lane0;
      toplevel_execute_ctrl4_up_AguPlugin_STORE_lane0 <= toplevel_execute_ctrl3_down_AguPlugin_STORE_lane0;
      toplevel_execute_ctrl4_up_AguPlugin_ATOMIC_lane0 <= toplevel_execute_ctrl3_down_AguPlugin_ATOMIC_lane0;
      toplevel_execute_ctrl4_up_AguPlugin_FLOAT_lane0 <= toplevel_execute_ctrl3_down_AguPlugin_FLOAT_lane0;
      toplevel_execute_ctrl4_up_LsuPlugin_logic_LSU_PREFETCH_lane0 <= toplevel_execute_ctrl3_down_LsuPlugin_logic_LSU_PREFETCH_lane0;
      toplevel_execute_ctrl4_up_late0_IntAluPlugin_ALU_ADD_SUB_lane0 <= toplevel_execute_ctrl3_down_late0_IntAluPlugin_ALU_ADD_SUB_lane0;
      toplevel_execute_ctrl4_up_late0_IntAluPlugin_ALU_SLTX_lane0 <= toplevel_execute_ctrl3_down_late0_IntAluPlugin_ALU_SLTX_lane0;
      toplevel_execute_ctrl4_up_late0_IntAluPlugin_ALU_BITWISE_CTRL_lane0 <= toplevel_execute_ctrl3_down_late0_IntAluPlugin_ALU_BITWISE_CTRL_lane0;
      toplevel_execute_ctrl4_up_early1_BranchPlugin_SEL_lane1 <= toplevel_execute_ctrl3_down_early1_BranchPlugin_SEL_lane1;
      toplevel_execute_ctrl4_up_late1_IntAluPlugin_SEL_lane1 <= toplevel_execute_ctrl3_down_late1_IntAluPlugin_SEL_lane1;
      toplevel_execute_ctrl4_up_late1_BarrelShifterPlugin_SEL_lane1 <= toplevel_execute_ctrl3_down_late1_BarrelShifterPlugin_SEL_lane1;
      toplevel_execute_ctrl4_up_late1_BranchPlugin_SEL_lane1 <= toplevel_execute_ctrl3_down_late1_BranchPlugin_SEL_lane1;
      toplevel_execute_ctrl4_up_lane1_integer_WriteBackPlugin_SEL_lane1 <= toplevel_execute_ctrl3_down_lane1_integer_WriteBackPlugin_SEL_lane1;
      toplevel_execute_ctrl4_up_COMPLETION_AT_4_lane1 <= toplevel_execute_ctrl3_down_COMPLETION_AT_4_lane1;
      toplevel_execute_ctrl4_up_execute_lane1_logic_completions_onCtrl_2_ENABLE_lane1 <= toplevel_execute_ctrl3_down_execute_lane1_logic_completions_onCtrl_2_ENABLE_lane1;
      toplevel_execute_ctrl4_up_SrcStageables_REVERT_lane1 <= toplevel_execute_ctrl3_down_SrcStageables_REVERT_lane1;
      toplevel_execute_ctrl4_up_SrcStageables_ZERO_lane1 <= toplevel_execute_ctrl3_down_SrcStageables_ZERO_lane1;
      toplevel_execute_ctrl4_up_SrcStageables_UNSIGNED_lane1 <= toplevel_execute_ctrl3_down_SrcStageables_UNSIGNED_lane1;
      toplevel_execute_ctrl4_up_BarrelShifterPlugin_LEFT_lane1 <= toplevel_execute_ctrl3_down_BarrelShifterPlugin_LEFT_lane1;
      toplevel_execute_ctrl4_up_BarrelShifterPlugin_SIGNED_lane1 <= toplevel_execute_ctrl3_down_BarrelShifterPlugin_SIGNED_lane1;
      toplevel_execute_ctrl4_up_BranchPlugin_BRANCH_CTRL_lane1 <= toplevel_execute_ctrl3_down_BranchPlugin_BRANCH_CTRL_lane1;
      toplevel_execute_ctrl4_up_late1_IntAluPlugin_ALU_ADD_SUB_lane1 <= toplevel_execute_ctrl3_down_late1_IntAluPlugin_ALU_ADD_SUB_lane1;
      toplevel_execute_ctrl4_up_late1_IntAluPlugin_ALU_SLTX_lane1 <= toplevel_execute_ctrl3_down_late1_IntAluPlugin_ALU_SLTX_lane1;
      toplevel_execute_ctrl4_up_late1_IntAluPlugin_ALU_BITWISE_CTRL_lane1 <= toplevel_execute_ctrl3_down_late1_IntAluPlugin_ALU_BITWISE_CTRL_lane1;
      toplevel_execute_ctrl4_up_COMMIT_lane0 <= toplevel_execute_ctrl3_down_COMMIT_lane0;
      toplevel_execute_ctrl4_up_COMMIT_lane1 <= toplevel_execute_ctrl3_down_COMMIT_lane1;
      toplevel_execute_ctrl4_up_early0_BranchPlugin_pcCalc_PC_TRUE_lane0 <= toplevel_execute_ctrl3_down_early0_BranchPlugin_pcCalc_PC_TRUE_lane0;
      toplevel_execute_ctrl4_up_early0_BranchPlugin_pcCalc_PC_FALSE_lane0 <= toplevel_execute_ctrl3_down_early0_BranchPlugin_pcCalc_PC_FALSE_lane0;
      toplevel_execute_ctrl4_up_early0_BranchPlugin_pcCalc_PC_LAST_SLICE_lane0 <= toplevel_execute_ctrl3_down_early0_BranchPlugin_pcCalc_PC_LAST_SLICE_lane0;
      toplevel_execute_ctrl4_up_early1_BranchPlugin_pcCalc_PC_TRUE_lane1 <= toplevel_execute_ctrl3_down_early1_BranchPlugin_pcCalc_PC_TRUE_lane1;
      toplevel_execute_ctrl4_up_early1_BranchPlugin_pcCalc_PC_FALSE_lane1 <= toplevel_execute_ctrl3_down_early1_BranchPlugin_pcCalc_PC_FALSE_lane1;
      toplevel_execute_ctrl4_up_early1_BranchPlugin_pcCalc_PC_LAST_SLICE_lane1 <= toplevel_execute_ctrl3_down_early1_BranchPlugin_pcCalc_PC_LAST_SLICE_lane1;
      toplevel_execute_ctrl4_up_lane0_integer_WriteBackPlugin_logic_DATA_lane0 <= toplevel_execute_ctrl3_down_lane0_integer_WriteBackPlugin_logic_DATA_lane0;
      toplevel_execute_ctrl4_up_lane1_integer_WriteBackPlugin_logic_DATA_lane1 <= toplevel_execute_ctrl3_down_lane1_integer_WriteBackPlugin_logic_DATA_lane1;
      toplevel_execute_ctrl4_up_LsuL1_MIXED_ADDRESS_lane0 <= toplevel_execute_ctrl3_down_LsuL1_MIXED_ADDRESS_lane0;
      toplevel_execute_ctrl4_up_LsuL1Plugin_logic_EVENT_WRITE_DATA_lane0 <= toplevel_execute_ctrl3_down_LsuL1Plugin_logic_EVENT_WRITE_DATA_lane0;
      toplevel_execute_ctrl4_up_LsuL1Plugin_logic_EVENT_WRITE_MASK_lane0 <= toplevel_execute_ctrl3_down_LsuL1Plugin_logic_EVENT_WRITE_MASK_lane0;
      toplevel_execute_ctrl4_up_LsuPlugin_logic_FROM_ACCESS_lane0 <= toplevel_execute_ctrl3_down_LsuPlugin_logic_FROM_ACCESS_lane0;
      toplevel_execute_ctrl4_up_LsuL1_MASK_lane0 <= toplevel_execute_ctrl3_down_LsuL1_MASK_lane0;
      toplevel_execute_ctrl4_up_LsuL1_SIZE_lane0 <= toplevel_execute_ctrl3_down_LsuL1_SIZE_lane0;
      toplevel_execute_ctrl4_up_LsuL1_LOAD_lane0 <= toplevel_execute_ctrl3_down_LsuL1_LOAD_lane0;
      toplevel_execute_ctrl4_up_LsuL1_ATOMIC_lane0 <= toplevel_execute_ctrl3_down_LsuL1_ATOMIC_lane0;
      toplevel_execute_ctrl4_up_LsuL1_STORE_lane0 <= toplevel_execute_ctrl3_down_LsuL1_STORE_lane0;
      toplevel_execute_ctrl4_up_LsuL1_PREFETCH_lane0 <= toplevel_execute_ctrl3_down_LsuL1_PREFETCH_lane0;
      toplevel_execute_ctrl4_up_LsuL1_FLUSH_lane0 <= toplevel_execute_ctrl3_down_LsuL1_FLUSH_lane0;
      toplevel_execute_ctrl4_up_Decode_STORE_ID_lane0 <= toplevel_execute_ctrl3_down_Decode_STORE_ID_lane0;
      toplevel_execute_ctrl4_up_LsuPlugin_logic_FROM_LSU_lane0 <= toplevel_execute_ctrl3_down_LsuPlugin_logic_FROM_LSU_lane0;
      toplevel_execute_ctrl4_up_LsuPlugin_logic_FROM_PREFETCH_lane0 <= toplevel_execute_ctrl3_down_LsuPlugin_logic_FROM_PREFETCH_lane0;
      toplevel_execute_ctrl4_up_LsuL1Plugin_logic_SHARED_lane0_plru_0 <= toplevel_execute_ctrl3_down_LsuL1Plugin_logic_SHARED_lane0_plru_0;
      toplevel_execute_ctrl4_up_LsuL1Plugin_logic_SHARED_lane0_dirty <= toplevel_execute_ctrl3_down_LsuL1Plugin_logic_SHARED_lane0_dirty;
      toplevel_execute_ctrl4_up_early0_MulPlugin_logic_steps_0_adders_0_lane0 <= toplevel_execute_ctrl3_down_early0_MulPlugin_logic_steps_0_adders_0_lane0;
      toplevel_execute_ctrl4_up_early0_MulPlugin_logic_steps_0_adders_1_lane0 <= toplevel_execute_ctrl3_down_early0_MulPlugin_logic_steps_0_adders_1_lane0;
      toplevel_execute_ctrl4_up_late0_SrcPlugin_SRC1_lane0 <= toplevel_execute_ctrl3_down_late0_SrcPlugin_SRC1_lane0;
      toplevel_execute_ctrl4_up_late0_SrcPlugin_SRC2_lane0 <= toplevel_execute_ctrl3_down_late0_SrcPlugin_SRC2_lane0;
      toplevel_execute_ctrl4_up_late1_SrcPlugin_SRC1_lane1 <= toplevel_execute_ctrl3_down_late1_SrcPlugin_SRC1_lane1;
      toplevel_execute_ctrl4_up_late1_SrcPlugin_SRC2_lane1 <= toplevel_execute_ctrl3_down_late1_SrcPlugin_SRC2_lane1;
      toplevel_execute_ctrl4_up_LsuL1Plugin_logic_BANK_BUSY_REMAPPED_lane0 <= toplevel_execute_ctrl3_down_LsuL1Plugin_logic_BANK_BUSY_REMAPPED_lane0;
      toplevel_execute_ctrl4_up_LsuL1Plugin_logic_BANKS_MUXES_lane0_0 <= toplevel_execute_ctrl3_down_LsuL1Plugin_logic_BANKS_MUXES_lane0_0;
      toplevel_execute_ctrl4_up_LsuL1Plugin_logic_BANKS_MUXES_lane0_1 <= toplevel_execute_ctrl3_down_LsuL1Plugin_logic_BANKS_MUXES_lane0_1;
      toplevel_execute_ctrl4_up_LsuL1Plugin_logic_WRITE_TO_READ_HAZARDS_lane0 <= toplevel_execute_ctrl3_down_LsuL1Plugin_logic_WRITE_TO_READ_HAZARDS_lane0;
      toplevel_execute_ctrl4_up_LsuL1_PHYSICAL_ADDRESS_lane0 <= toplevel_execute_ctrl3_down_LsuL1_PHYSICAL_ADDRESS_lane0;
      toplevel_execute_ctrl4_up_LsuL1Plugin_logic_WAYS_TAGS_lane0_0_loaded <= toplevel_execute_ctrl3_down_LsuL1Plugin_logic_WAYS_TAGS_lane0_0_loaded;
      toplevel_execute_ctrl4_up_LsuL1Plugin_logic_WAYS_TAGS_lane0_0_address <= toplevel_execute_ctrl3_down_LsuL1Plugin_logic_WAYS_TAGS_lane0_0_address;
      toplevel_execute_ctrl4_up_LsuL1Plugin_logic_WAYS_TAGS_lane0_0_fault <= toplevel_execute_ctrl3_down_LsuL1Plugin_logic_WAYS_TAGS_lane0_0_fault;
      toplevel_execute_ctrl4_up_LsuL1Plugin_logic_WAYS_TAGS_lane0_1_loaded <= toplevel_execute_ctrl3_down_LsuL1Plugin_logic_WAYS_TAGS_lane0_1_loaded;
      toplevel_execute_ctrl4_up_LsuL1Plugin_logic_WAYS_TAGS_lane0_1_address <= toplevel_execute_ctrl3_down_LsuL1Plugin_logic_WAYS_TAGS_lane0_1_address;
      toplevel_execute_ctrl4_up_LsuL1Plugin_logic_WAYS_TAGS_lane0_1_fault <= toplevel_execute_ctrl3_down_LsuL1Plugin_logic_WAYS_TAGS_lane0_1_fault;
      toplevel_execute_ctrl4_up_LsuL1Plugin_logic_WAYS_HITS_lane0 <= toplevel_execute_ctrl3_down_LsuL1Plugin_logic_WAYS_HITS_lane0;
      toplevel_execute_ctrl4_up_LsuPlugin_logic_onTrigger_HIT_lane0 <= toplevel_execute_ctrl3_down_LsuPlugin_logic_onTrigger_HIT_lane0;
      toplevel_execute_ctrl4_up_MMU_TRANSLATED_lane0 <= toplevel_execute_ctrl3_down_MMU_TRANSLATED_lane0;
      toplevel_execute_ctrl4_up_LsuPlugin_logic_preCtrl_MISS_ALIGNED_lane0 <= toplevel_execute_ctrl3_down_LsuPlugin_logic_preCtrl_MISS_ALIGNED_lane0;
      toplevel_execute_ctrl4_up_LsuPlugin_logic_preCtrl_IS_AMO_lane0 <= toplevel_execute_ctrl3_down_LsuPlugin_logic_preCtrl_IS_AMO_lane0;
      toplevel_execute_ctrl4_up_LsuPlugin_logic_onPma_CACHED_RSP_lane0_fault <= toplevel_execute_ctrl3_down_LsuPlugin_logic_onPma_CACHED_RSP_lane0_fault;
      toplevel_execute_ctrl4_up_LsuPlugin_logic_onPma_CACHED_RSP_lane0_io <= toplevel_execute_ctrl3_down_LsuPlugin_logic_onPma_CACHED_RSP_lane0_io;
      toplevel_execute_ctrl4_up_LsuPlugin_logic_onPma_IO_RSP_lane0_fault <= toplevel_execute_ctrl3_down_LsuPlugin_logic_onPma_IO_RSP_lane0_fault;
      toplevel_execute_ctrl4_up_LsuPlugin_logic_onPma_IO_RSP_lane0_io <= toplevel_execute_ctrl3_down_LsuPlugin_logic_onPma_IO_RSP_lane0_io;
      toplevel_execute_ctrl4_up_LsuPlugin_logic_onPma_IO_lane0 <= toplevel_execute_ctrl3_down_LsuPlugin_logic_onPma_IO_lane0;
      toplevel_execute_ctrl4_up_LsuPlugin_logic_onPma_FROM_LSU_MSB_FAILED_lane0 <= toplevel_execute_ctrl3_down_LsuPlugin_logic_onPma_FROM_LSU_MSB_FAILED_lane0;
      toplevel_execute_ctrl4_up_LsuPlugin_logic_MMU_PAGE_FAULT_lane0 <= toplevel_execute_ctrl3_down_LsuPlugin_logic_MMU_PAGE_FAULT_lane0;
      toplevel_execute_ctrl4_up_LsuPlugin_logic_MMU_FAILURE_lane0 <= toplevel_execute_ctrl3_down_LsuPlugin_logic_MMU_FAILURE_lane0;
      toplevel_execute_ctrl4_up_MMU_ACCESS_FAULT_lane0 <= toplevel_execute_ctrl3_down_MMU_ACCESS_FAULT_lane0;
      toplevel_execute_ctrl4_up_MMU_REFILL_lane0 <= toplevel_execute_ctrl3_down_MMU_REFILL_lane0;
      toplevel_execute_ctrl4_up_MMU_HAZARD_lane0 <= toplevel_execute_ctrl3_down_MMU_HAZARD_lane0;
      toplevel_execute_ctrl4_up_MMU_BYPASS_TRANSLATION_lane0 <= toplevel_execute_ctrl3_down_MMU_BYPASS_TRANSLATION_lane0;
    end
    if(toplevel_execute_ctrl4_down_isReady) begin
      toplevel_execute_ctrl5_up_RD_ENABLE_lane0 <= toplevel_execute_ctrl4_down_RD_ENABLE_lane0;
      toplevel_execute_ctrl5_up_RD_PHYS_lane0 <= toplevel_execute_ctrl4_down_RD_PHYS_lane0;
      toplevel_execute_ctrl5_up_LANE_AGE_lane0 <= toplevel_execute_ctrl4_down_LANE_AGE_lane0;
      toplevel_execute_ctrl5_up_RD_ENABLE_lane1 <= toplevel_execute_ctrl4_down_RD_ENABLE_lane1;
      toplevel_execute_ctrl5_up_RD_PHYS_lane1 <= toplevel_execute_ctrl4_down_RD_PHYS_lane1;
      toplevel_execute_ctrl5_up_LANE_AGE_lane1 <= toplevel_execute_ctrl4_down_LANE_AGE_lane1;
      toplevel_execute_ctrl5_up_COMMIT_lane0 <= toplevel_execute_ctrl4_down_COMMIT_lane0;
      toplevel_execute_ctrl5_up_COMMIT_lane1 <= toplevel_execute_ctrl4_down_COMMIT_lane1;
      toplevel_execute_ctrl5_up_lane0_integer_WriteBackPlugin_logic_DATA_lane0 <= toplevel_execute_ctrl4_down_lane0_integer_WriteBackPlugin_logic_DATA_lane0;
      toplevel_execute_ctrl5_up_lane1_integer_WriteBackPlugin_logic_DATA_lane1 <= toplevel_execute_ctrl4_down_lane1_integer_WriteBackPlugin_logic_DATA_lane1;
    end
    case(LsuPlugin_logic_flusher_stateReg)
      LsuPlugin_logic_flusher_enumDef_CMD : begin
        if(when_LsuPlugin_l297) begin
          LsuPlugin_logic_flusher_waiter <= LsuL1_WRITEBACK_BUSY;
        end
      end
      LsuPlugin_logic_flusher_enumDef_COMPLETION : begin
        LsuPlugin_logic_flusher_waiter <= (LsuPlugin_logic_flusher_waiter & LsuL1_WRITEBACK_BUSY);
      end
      default : begin
        LsuPlugin_logic_flusher_cmdCounter <= 7'h0;
      end
    endcase
    case(TrapPlugin_logic_harts_0_trap_fsm_stateReg)
      TrapPlugin_logic_harts_0_trap_fsm_enumDef_RUNNING : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_enumDef_PROCESS_1 : begin
        TrapPlugin_logic_harts_0_trap_fsm_triggerEbreakReg <= TrapPlugin_logic_harts_0_trap_fsm_triggerEbreak;
      end
      TrapPlugin_logic_harts_0_trap_fsm_enumDef_TRAP_EPC : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_enumDef_TRAP_TVAL : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_enumDef_TRAP_TVEC : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_enumDef_TRAP_APPLY : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_enumDef_XRET_EPC : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_enumDef_XRET_APPLY : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_enumDef_ATS_RSP : begin
        if(TrapPlugin_logic_harts_0_trap_fsm_atsPorts_refill_rsp_valid) begin
          if(when_TrapPlugin_l492) begin
            TrapPlugin_logic_harts_0_trap_pending_state_exception <= 1'b1;
            case(switch_TrapPlugin_l494)
              3'b010 : begin
                TrapPlugin_logic_harts_0_trap_pending_state_code <= 4'b0001;
              end
              3'b000 : begin
                TrapPlugin_logic_harts_0_trap_pending_state_code <= 4'b0101;
              end
              3'b001 : begin
                TrapPlugin_logic_harts_0_trap_pending_state_code <= 4'b0111;
              end
              3'b110 : begin
                TrapPlugin_logic_harts_0_trap_pending_state_code <= 4'b1100;
              end
              3'b100 : begin
                TrapPlugin_logic_harts_0_trap_pending_state_code <= 4'b1101;
              end
              3'b101 : begin
                TrapPlugin_logic_harts_0_trap_pending_state_code <= 4'b1111;
              end
              default : begin
              end
            endcase
          end
        end
      end
      TrapPlugin_logic_harts_0_trap_fsm_enumDef_JUMP : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_enumDef_LSU_FLUSH : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_enumDef_FETCH_FLUSH : begin
      end
      default : begin
      end
    endcase
    case(MmuPlugin_logic_refill_stateReg)
      MmuPlugin_logic_refill_enumDef_IDLE : begin
        if(MmuPlugin_logic_refill_arbiter_io_output_valid) begin
          MmuPlugin_logic_refill_portOhReg <= MmuPlugin_logic_refill_arbiter_io_chosenOH;
          MmuPlugin_logic_refill_storageOhReg <= (2'b01 <<< MmuPlugin_logic_refill_arbiter_io_output_payload_storageId);
          MmuPlugin_logic_refill_virtual <= MmuPlugin_logic_refill_arbiter_io_output_payload_address;
          MmuPlugin_logic_refill_load_address <= {{MmuPlugin_logic_satp_ppn,MmuPlugin_logic_refill_arbiter_io_output_payload_address[31 : 22]},2'b00};
        end
      end
      MmuPlugin_logic_refill_enumDef_CMD_0 : begin
      end
      MmuPlugin_logic_refill_enumDef_CMD_1 : begin
      end
      MmuPlugin_logic_refill_enumDef_RSP_0 : begin
      end
      MmuPlugin_logic_refill_enumDef_RSP_1 : begin
        if(MmuPlugin_logic_refill_load_rsp_valid) begin
          if(!MmuPlugin_logic_refill_load_rsp_payload_redo) begin
            if(!when_MmuPlugin_l471) begin
              MmuPlugin_logic_refill_load_address <= MmuPlugin_logic_refill_load_nextLevelBase;
              MmuPlugin_logic_refill_load_address[11 : 2] <= MmuPlugin_logic_refill_virtual[21 : 12];
            end
          end
        end
      end
      default : begin
      end
    endcase
    case(CsrAccessPlugin_logic_fsm_stateReg)
      CsrAccessPlugin_logic_fsm_enumDef_READ : begin
        CsrAccessPlugin_logic_fsm_regs_aluInput <= CsrAccessPlugin_bus_read_toWriteBits;
        CsrAccessPlugin_logic_fsm_regs_csrValue <= CsrAccessPlugin_logic_fsm_readLogic_csrValue;
      end
      CsrAccessPlugin_logic_fsm_enumDef_WRITE : begin
      end
      CsrAccessPlugin_logic_fsm_enumDef_COMPLETION : begin
      end
      default : begin
        REG_CSR_1952 <= COMB_CSR_1952;
        REG_CSR_1953 <= COMB_CSR_1953;
        REG_CSR_1954 <= COMB_CSR_1954;
        REG_CSR_3857 <= COMB_CSR_3857;
        REG_CSR_3858 <= COMB_CSR_3858;
        REG_CSR_3859 <= COMB_CSR_3859;
        REG_CSR_3860 <= COMB_CSR_3860;
        REG_CSR_769 <= COMB_CSR_769;
        REG_CSR_768 <= COMB_CSR_768;
        REG_CSR_834 <= COMB_CSR_834;
        REG_CSR_836 <= COMB_CSR_836;
        REG_CSR_772 <= COMB_CSR_772;
        REG_CSR_770 <= COMB_CSR_770;
        REG_CSR_771 <= COMB_CSR_771;
        REG_CSR_322 <= COMB_CSR_322;
        REG_CSR_256 <= COMB_CSR_256;
        REG_CSR_260 <= COMB_CSR_260;
        REG_CSR_324 <= COMB_CSR_324;
        REG_CSR_3073 <= COMB_CSR_3073;
        REG_CSR_3201 <= COMB_CSR_3201;
        REG_CSR_PrivilegedPlugin_logic_readAnyWriteLegal_tvecFilter <= COMB_CSR_PrivilegedPlugin_logic_readAnyWriteLegal_tvecFilter;
        REG_CSR_PrivilegedPlugin_logic_readAnyWriteLegal_epcFilter <= COMB_CSR_PrivilegedPlugin_logic_readAnyWriteLegal_epcFilter;
        REG_CSR_384 <= COMB_CSR_384;
        REG_CSR_CsrRamPlugin_csrMapper_selFilter <= COMB_CSR_CsrRamPlugin_csrMapper_selFilter;
        REG_CSR_CsrAccessPlugin_logic_trapNextOnWriteFilter <= COMB_CSR_CsrAccessPlugin_logic_trapNextOnWriteFilter;
      end
    endcase
  end


endmodule

module Apb3Router (
  input  wire [18:0]   io_input_PADDR,
  input  wire [4:0]    io_input_PSEL,
  input  wire          io_input_PENABLE,
  output wire          io_input_PREADY,
  input  wire          io_input_PWRITE,
  input  wire [31:0]   io_input_PWDATA,
  output wire [31:0]   io_input_PRDATA,
  output wire [18:0]   io_outputs_0_PADDR,
  output wire [0:0]    io_outputs_0_PSEL,
  output wire          io_outputs_0_PENABLE,
  input  wire          io_outputs_0_PREADY,
  output wire          io_outputs_0_PWRITE,
  output wire [31:0]   io_outputs_0_PWDATA,
  input  wire [31:0]   io_outputs_0_PRDATA,
  output wire [18:0]   io_outputs_1_PADDR,
  output wire [0:0]    io_outputs_1_PSEL,
  output wire          io_outputs_1_PENABLE,
  input  wire          io_outputs_1_PREADY,
  output wire          io_outputs_1_PWRITE,
  output wire [31:0]   io_outputs_1_PWDATA,
  input  wire [31:0]   io_outputs_1_PRDATA,
  output wire [18:0]   io_outputs_2_PADDR,
  output wire [0:0]    io_outputs_2_PSEL,
  output wire          io_outputs_2_PENABLE,
  input  wire          io_outputs_2_PREADY,
  output wire          io_outputs_2_PWRITE,
  output wire [31:0]   io_outputs_2_PWDATA,
  input  wire [31:0]   io_outputs_2_PRDATA,
  output wire [18:0]   io_outputs_3_PADDR,
  output wire [0:0]    io_outputs_3_PSEL,
  output wire          io_outputs_3_PENABLE,
  input  wire          io_outputs_3_PREADY,
  output wire          io_outputs_3_PWRITE,
  output wire [31:0]   io_outputs_3_PWDATA,
  input  wire [31:0]   io_outputs_3_PRDATA,
  output wire [18:0]   io_outputs_4_PADDR,
  output wire [0:0]    io_outputs_4_PSEL,
  output wire          io_outputs_4_PENABLE,
  input  wire          io_outputs_4_PREADY,
  output wire          io_outputs_4_PWRITE,
  output wire [31:0]   io_outputs_4_PWDATA,
  input  wire [31:0]   io_outputs_4_PRDATA,
  input  wire          clk_peripheral,
  input  wire          reset_peripheral
);

  reg                 _zz_io_input_PREADY;
  reg        [31:0]   _zz_io_input_PRDATA;
  wire                _zz_selIndex;
  wire                _zz_selIndex_1;
  wire                _zz_selIndex_2;
  wire                _zz_selIndex_3;
  reg        [2:0]    selIndex;

  always @(*) begin
    case(selIndex)
      3'b000 : begin
        _zz_io_input_PREADY = io_outputs_0_PREADY;
        _zz_io_input_PRDATA = io_outputs_0_PRDATA;
      end
      3'b001 : begin
        _zz_io_input_PREADY = io_outputs_1_PREADY;
        _zz_io_input_PRDATA = io_outputs_1_PRDATA;
      end
      3'b010 : begin
        _zz_io_input_PREADY = io_outputs_2_PREADY;
        _zz_io_input_PRDATA = io_outputs_2_PRDATA;
      end
      3'b011 : begin
        _zz_io_input_PREADY = io_outputs_3_PREADY;
        _zz_io_input_PRDATA = io_outputs_3_PRDATA;
      end
      default : begin
        _zz_io_input_PREADY = io_outputs_4_PREADY;
        _zz_io_input_PRDATA = io_outputs_4_PRDATA;
      end
    endcase
  end

  assign io_outputs_0_PADDR = io_input_PADDR;
  assign io_outputs_0_PENABLE = io_input_PENABLE;
  assign io_outputs_0_PSEL[0] = io_input_PSEL[0];
  assign io_outputs_0_PWRITE = io_input_PWRITE;
  assign io_outputs_0_PWDATA = io_input_PWDATA;
  assign io_outputs_1_PADDR = io_input_PADDR;
  assign io_outputs_1_PENABLE = io_input_PENABLE;
  assign io_outputs_1_PSEL[0] = io_input_PSEL[1];
  assign io_outputs_1_PWRITE = io_input_PWRITE;
  assign io_outputs_1_PWDATA = io_input_PWDATA;
  assign io_outputs_2_PADDR = io_input_PADDR;
  assign io_outputs_2_PENABLE = io_input_PENABLE;
  assign io_outputs_2_PSEL[0] = io_input_PSEL[2];
  assign io_outputs_2_PWRITE = io_input_PWRITE;
  assign io_outputs_2_PWDATA = io_input_PWDATA;
  assign io_outputs_3_PADDR = io_input_PADDR;
  assign io_outputs_3_PENABLE = io_input_PENABLE;
  assign io_outputs_3_PSEL[0] = io_input_PSEL[3];
  assign io_outputs_3_PWRITE = io_input_PWRITE;
  assign io_outputs_3_PWDATA = io_input_PWDATA;
  assign io_outputs_4_PADDR = io_input_PADDR;
  assign io_outputs_4_PENABLE = io_input_PENABLE;
  assign io_outputs_4_PSEL[0] = io_input_PSEL[4];
  assign io_outputs_4_PWRITE = io_input_PWRITE;
  assign io_outputs_4_PWDATA = io_input_PWDATA;
  assign _zz_selIndex = io_input_PSEL[3];
  assign _zz_selIndex_1 = io_input_PSEL[4];
  assign _zz_selIndex_2 = (io_input_PSEL[1] || _zz_selIndex);
  assign _zz_selIndex_3 = (io_input_PSEL[2] || _zz_selIndex);
  assign io_input_PREADY = _zz_io_input_PREADY;
  assign io_input_PRDATA = _zz_io_input_PRDATA;
  always @(posedge clk_peripheral) begin
    selIndex <= {_zz_selIndex_1,{_zz_selIndex_3,_zz_selIndex_2}};
  end


endmodule

module Apb3Decoder (
  input  wire [18:0]   io_input_PADDR,
  input  wire [0:0]    io_input_PSEL,
  input  wire          io_input_PENABLE,
  output reg           io_input_PREADY,
  input  wire          io_input_PWRITE,
  input  wire [31:0]   io_input_PWDATA,
  output wire [31:0]   io_input_PRDATA,
  output wire [18:0]   io_output_PADDR,
  output reg  [4:0]    io_output_PSEL,
  output wire          io_output_PENABLE,
  input  wire          io_output_PREADY,
  output wire          io_output_PWRITE,
  output wire [31:0]   io_output_PWDATA,
  input  wire [31:0]   io_output_PRDATA
);

  wire                when_Apb3Decoder_l88;

  assign io_output_PADDR = io_input_PADDR;
  assign io_output_PENABLE = io_input_PENABLE;
  assign io_output_PWRITE = io_input_PWRITE;
  assign io_output_PWDATA = io_input_PWDATA;
  always @(*) begin
    io_output_PSEL[0] = (((io_input_PADDR & (~ 19'h0000f)) == 19'h10000) && io_input_PSEL[0]);
    io_output_PSEL[1] = (((io_input_PADDR & (~ 19'h00007)) == 19'h20000) && io_input_PSEL[0]);
    io_output_PSEL[2] = (((io_input_PADDR & (~ 19'h0001f)) == 19'h30000) && io_input_PSEL[0]);
    io_output_PSEL[3] = (((io_input_PADDR & (~ 19'h00fff)) == 19'h40000) && io_input_PSEL[0]);
    io_output_PSEL[4] = (((io_input_PADDR & (~ 19'h00fff)) == 19'h41000) && io_input_PSEL[0]);
  end

  always @(*) begin
    io_input_PREADY = io_output_PREADY;
    if(when_Apb3Decoder_l88) begin
      io_input_PREADY = 1'b1;
    end
  end

  assign io_input_PRDATA = io_output_PRDATA;
  assign when_Apb3Decoder_l88 = (io_input_PSEL[0] && (io_output_PSEL == 5'h0));

endmodule

module EndeavourUSB (
  inout  wire          io_usb1_dp,
  inout  wire          io_usb1_dn,
  inout  wire          io_usb2_dp,
  inout  wire          io_usb2_dn,
  input  wire [11:0]   io_apb_ctrl_PADDR,
  input  wire [0:0]    io_apb_ctrl_PSEL,
  input  wire          io_apb_ctrl_PENABLE,
  output wire          io_apb_ctrl_PREADY,
  input  wire          io_apb_ctrl_PWRITE,
  input  wire [31:0]   io_apb_ctrl_PWDATA,
  output wire [31:0]   io_apb_ctrl_PRDATA,
  input  wire [11:0]   io_apb_dma_PADDR,
  input  wire [0:0]    io_apb_dma_PSEL,
  input  wire          io_apb_dma_PENABLE,
  output wire          io_apb_dma_PREADY,
  input  wire          io_apb_dma_PWRITE,
  input  wire [31:0]   io_apb_dma_PWDATA,
  output wire [31:0]   io_apb_dma_PRDATA,
  output wire          io_interrupt,
  output wire          _zz_io_interrupt,
  input  wire          clk_peripheral,
  input  wire          reset_peripheral
);

  wire                ohci_io_ctrl_cmd_valid;
  wire       [0:0]    ohci_io_ctrl_cmd_payload_fragment_opcode;
  wire       [11:0]   ram_1_io_buses_0_cmd_payload_fragment_address;
  wire                ram_1_io_buses_1_cmd_valid;
  wire       [0:0]    ram_1_io_buses_1_cmd_payload_fragment_opcode;
  wire                ohci_io_ctrl_cmd_ready;
  wire                ohci_io_ctrl_rsp_valid;
  wire                ohci_io_ctrl_rsp_payload_last;
  wire       [0:0]    ohci_io_ctrl_rsp_payload_fragment_opcode;
  wire       [31:0]   ohci_io_ctrl_rsp_payload_fragment_data;
  wire                ohci_io_phy_lowSpeed;
  wire                ohci_io_phy_usbReset;
  wire                ohci_io_phy_usbResume;
  wire                ohci_io_phy_tx_valid;
  wire                ohci_io_phy_tx_payload_last;
  wire       [7:0]    ohci_io_phy_tx_payload_fragment;
  wire                ohci_io_phy_ports_0_removable;
  wire                ohci_io_phy_ports_0_power;
  wire                ohci_io_phy_ports_0_reset_valid;
  wire                ohci_io_phy_ports_0_suspend_valid;
  wire                ohci_io_phy_ports_0_resume_valid;
  wire                ohci_io_phy_ports_0_disable_valid;
  wire                ohci_io_phy_ports_1_removable;
  wire                ohci_io_phy_ports_1_power;
  wire                ohci_io_phy_ports_1_reset_valid;
  wire                ohci_io_phy_ports_1_suspend_valid;
  wire                ohci_io_phy_ports_1_resume_valid;
  wire                ohci_io_phy_ports_1_disable_valid;
  wire                ohci_io_dma_cmd_valid;
  wire                ohci_io_dma_cmd_payload_last;
  wire       [0:0]    ohci_io_dma_cmd_payload_fragment_opcode;
  wire       [31:0]   ohci_io_dma_cmd_payload_fragment_address;
  wire       [5:0]    ohci_io_dma_cmd_payload_fragment_length;
  wire       [31:0]   ohci_io_dma_cmd_payload_fragment_data;
  wire       [3:0]    ohci_io_dma_cmd_payload_fragment_mask;
  wire                ohci_io_dma_rsp_ready;
  wire                ohci_io_interrupt;
  wire                ohci_io_interruptBios;
  wire                phy_io_ctrl_overcurrent;
  wire                phy_io_ctrl_tick;
  wire                phy_io_ctrl_tx_ready;
  wire                phy_io_ctrl_txEop;
  wire                phy_io_ctrl_rx_flow_valid;
  wire                phy_io_ctrl_rx_flow_payload_stuffingError;
  wire       [7:0]    phy_io_ctrl_rx_flow_payload_data;
  wire                phy_io_ctrl_rx_active;
  wire                phy_io_ctrl_ports_0_reset_ready;
  wire                phy_io_ctrl_ports_0_suspend_ready;
  wire                phy_io_ctrl_ports_0_resume_ready;
  wire                phy_io_ctrl_ports_0_disable_ready;
  wire                phy_io_ctrl_ports_0_connect;
  wire                phy_io_ctrl_ports_0_disconnect;
  wire                phy_io_ctrl_ports_0_overcurrent;
  wire                phy_io_ctrl_ports_0_lowSpeed;
  wire                phy_io_ctrl_ports_0_remoteResume;
  wire                phy_io_ctrl_ports_1_reset_ready;
  wire                phy_io_ctrl_ports_1_suspend_ready;
  wire                phy_io_ctrl_ports_1_resume_ready;
  wire                phy_io_ctrl_ports_1_disable_ready;
  wire                phy_io_ctrl_ports_1_connect;
  wire                phy_io_ctrl_ports_1_disconnect;
  wire                phy_io_ctrl_ports_1_overcurrent;
  wire                phy_io_ctrl_ports_1_lowSpeed;
  wire                phy_io_ctrl_ports_1_remoteResume;
  wire                phy_io_usb_0_tx_enable;
  wire                phy_io_usb_0_tx_data;
  wire                phy_io_usb_0_tx_se0;
  wire                phy_io_usb_1_tx_enable;
  wire                phy_io_usb_1_tx_data;
  wire                phy_io_usb_1_tx_se0;
  wire                phy_io_management_0_power;
  wire                phy_io_management_1_power;
  wire                ram_1_io_buses_0_cmd_ready;
  wire                ram_1_io_buses_0_rsp_valid;
  wire                ram_1_io_buses_0_rsp_payload_last;
  wire       [0:0]    ram_1_io_buses_0_rsp_payload_fragment_opcode;
  wire       [31:0]   ram_1_io_buses_0_rsp_payload_fragment_data;
  wire                ram_1_io_buses_1_cmd_ready;
  wire                ram_1_io_buses_1_rsp_valid;
  wire                ram_1_io_buses_1_rsp_payload_last;
  wire       [0:0]    ram_1_io_buses_1_rsp_payload_fragment_opcode;
  wire       [31:0]   ram_1_io_buses_1_rsp_payload_fragment_data;
  reg                 _zz_io_usb2_dn;
  reg                 _zz_io_usb2_dp;
  reg                 _zz_io_usb1_dn;
  reg                 _zz_io_usb1_dp;
  wire                usb1_tri_dp_read;
  wire                usb1_tri_dp_write;
  wire                usb1_tri_dp_writeEnable;
  wire                usb1_tri_dm_read;
  wire                usb1_tri_dm_write;
  wire                usb1_tri_dm_writeEnable;
  wire                usb2_tri_dp_read;
  wire                usb2_tri_dp_write;
  wire                usb2_tri_dp_writeEnable;
  wire                usb2_tri_dm_read;
  wire                usb2_tri_dm_write;
  wire                usb2_tri_dm_writeEnable;
  wire                _zz_when_usb_l96;
  reg                 _zz_when_usb_l96_1;
  wire                when_usb_l96;
  wire                when_usb_l96_1;
  wire                _zz_when_usb_l96_2;
  reg                 _zz_when_usb_l96_3;
  wire                when_usb_l96_2;
  wire                when_usb_l96_3;

  UsbOhci ohci (
    .io_ctrl_cmd_valid                    (ohci_io_ctrl_cmd_valid                          ), //i
    .io_ctrl_cmd_ready                    (ohci_io_ctrl_cmd_ready                          ), //o
    .io_ctrl_cmd_payload_last             (1'b1                                            ), //i
    .io_ctrl_cmd_payload_fragment_opcode  (ohci_io_ctrl_cmd_payload_fragment_opcode        ), //i
    .io_ctrl_cmd_payload_fragment_address (io_apb_ctrl_PADDR[11:0]                         ), //i
    .io_ctrl_cmd_payload_fragment_length  (2'b11                                           ), //i
    .io_ctrl_cmd_payload_fragment_data    (io_apb_ctrl_PWDATA[31:0]                        ), //i
    .io_ctrl_cmd_payload_fragment_mask    (4'b1111                                         ), //i
    .io_ctrl_rsp_valid                    (ohci_io_ctrl_rsp_valid                          ), //o
    .io_ctrl_rsp_ready                    (1'b1                                            ), //i
    .io_ctrl_rsp_payload_last             (ohci_io_ctrl_rsp_payload_last                   ), //o
    .io_ctrl_rsp_payload_fragment_opcode  (ohci_io_ctrl_rsp_payload_fragment_opcode        ), //o
    .io_ctrl_rsp_payload_fragment_data    (ohci_io_ctrl_rsp_payload_fragment_data[31:0]    ), //o
    .io_phy_lowSpeed                      (ohci_io_phy_lowSpeed                            ), //o
    .io_phy_tx_valid                      (ohci_io_phy_tx_valid                            ), //o
    .io_phy_tx_ready                      (phy_io_ctrl_tx_ready                            ), //i
    .io_phy_tx_payload_last               (ohci_io_phy_tx_payload_last                     ), //o
    .io_phy_tx_payload_fragment           (ohci_io_phy_tx_payload_fragment[7:0]            ), //o
    .io_phy_txEop                         (phy_io_ctrl_txEop                               ), //i
    .io_phy_rx_flow_valid                 (phy_io_ctrl_rx_flow_valid                       ), //i
    .io_phy_rx_flow_payload_stuffingError (phy_io_ctrl_rx_flow_payload_stuffingError       ), //i
    .io_phy_rx_flow_payload_data          (phy_io_ctrl_rx_flow_payload_data[7:0]           ), //i
    .io_phy_rx_active                     (phy_io_ctrl_rx_active                           ), //i
    .io_phy_usbReset                      (ohci_io_phy_usbReset                            ), //o
    .io_phy_usbResume                     (ohci_io_phy_usbResume                           ), //o
    .io_phy_overcurrent                   (phy_io_ctrl_overcurrent                         ), //i
    .io_phy_tick                          (phy_io_ctrl_tick                                ), //i
    .io_phy_ports_0_disable_valid         (ohci_io_phy_ports_0_disable_valid               ), //o
    .io_phy_ports_0_disable_ready         (phy_io_ctrl_ports_0_disable_ready               ), //i
    .io_phy_ports_0_removable             (ohci_io_phy_ports_0_removable                   ), //o
    .io_phy_ports_0_power                 (ohci_io_phy_ports_0_power                       ), //o
    .io_phy_ports_0_reset_valid           (ohci_io_phy_ports_0_reset_valid                 ), //o
    .io_phy_ports_0_reset_ready           (phy_io_ctrl_ports_0_reset_ready                 ), //i
    .io_phy_ports_0_suspend_valid         (ohci_io_phy_ports_0_suspend_valid               ), //o
    .io_phy_ports_0_suspend_ready         (phy_io_ctrl_ports_0_suspend_ready               ), //i
    .io_phy_ports_0_resume_valid          (ohci_io_phy_ports_0_resume_valid                ), //o
    .io_phy_ports_0_resume_ready          (phy_io_ctrl_ports_0_resume_ready                ), //i
    .io_phy_ports_0_connect               (phy_io_ctrl_ports_0_connect                     ), //i
    .io_phy_ports_0_disconnect            (phy_io_ctrl_ports_0_disconnect                  ), //i
    .io_phy_ports_0_overcurrent           (phy_io_ctrl_ports_0_overcurrent                 ), //i
    .io_phy_ports_0_remoteResume          (phy_io_ctrl_ports_0_remoteResume                ), //i
    .io_phy_ports_0_lowSpeed              (phy_io_ctrl_ports_0_lowSpeed                    ), //i
    .io_phy_ports_1_disable_valid         (ohci_io_phy_ports_1_disable_valid               ), //o
    .io_phy_ports_1_disable_ready         (phy_io_ctrl_ports_1_disable_ready               ), //i
    .io_phy_ports_1_removable             (ohci_io_phy_ports_1_removable                   ), //o
    .io_phy_ports_1_power                 (ohci_io_phy_ports_1_power                       ), //o
    .io_phy_ports_1_reset_valid           (ohci_io_phy_ports_1_reset_valid                 ), //o
    .io_phy_ports_1_reset_ready           (phy_io_ctrl_ports_1_reset_ready                 ), //i
    .io_phy_ports_1_suspend_valid         (ohci_io_phy_ports_1_suspend_valid               ), //o
    .io_phy_ports_1_suspend_ready         (phy_io_ctrl_ports_1_suspend_ready               ), //i
    .io_phy_ports_1_resume_valid          (ohci_io_phy_ports_1_resume_valid                ), //o
    .io_phy_ports_1_resume_ready          (phy_io_ctrl_ports_1_resume_ready                ), //i
    .io_phy_ports_1_connect               (phy_io_ctrl_ports_1_connect                     ), //i
    .io_phy_ports_1_disconnect            (phy_io_ctrl_ports_1_disconnect                  ), //i
    .io_phy_ports_1_overcurrent           (phy_io_ctrl_ports_1_overcurrent                 ), //i
    .io_phy_ports_1_remoteResume          (phy_io_ctrl_ports_1_remoteResume                ), //i
    .io_phy_ports_1_lowSpeed              (phy_io_ctrl_ports_1_lowSpeed                    ), //i
    .io_dma_cmd_valid                     (ohci_io_dma_cmd_valid                           ), //o
    .io_dma_cmd_ready                     (ram_1_io_buses_0_cmd_ready                      ), //i
    .io_dma_cmd_payload_last              (ohci_io_dma_cmd_payload_last                    ), //o
    .io_dma_cmd_payload_fragment_opcode   (ohci_io_dma_cmd_payload_fragment_opcode         ), //o
    .io_dma_cmd_payload_fragment_address  (ohci_io_dma_cmd_payload_fragment_address[31:0]  ), //o
    .io_dma_cmd_payload_fragment_length   (ohci_io_dma_cmd_payload_fragment_length[5:0]    ), //o
    .io_dma_cmd_payload_fragment_data     (ohci_io_dma_cmd_payload_fragment_data[31:0]     ), //o
    .io_dma_cmd_payload_fragment_mask     (ohci_io_dma_cmd_payload_fragment_mask[3:0]      ), //o
    .io_dma_rsp_valid                     (ram_1_io_buses_0_rsp_valid                      ), //i
    .io_dma_rsp_ready                     (ohci_io_dma_rsp_ready                           ), //o
    .io_dma_rsp_payload_last              (ram_1_io_buses_0_rsp_payload_last               ), //i
    .io_dma_rsp_payload_fragment_opcode   (ram_1_io_buses_0_rsp_payload_fragment_opcode    ), //i
    .io_dma_rsp_payload_fragment_data     (ram_1_io_buses_0_rsp_payload_fragment_data[31:0]), //i
    .io_interrupt                         (ohci_io_interrupt                               ), //o
    .io_interruptBios                     (ohci_io_interruptBios                           ), //o
    .clk_peripheral                       (clk_peripheral                                  ), //i
    .reset_peripheral                     (reset_peripheral                                )  //i
  );
  UsbLsFsPhyModified phy (
    .io_ctrl_lowSpeed                      (ohci_io_phy_lowSpeed                     ), //i
    .io_ctrl_tx_valid                      (ohci_io_phy_tx_valid                     ), //i
    .io_ctrl_tx_ready                      (phy_io_ctrl_tx_ready                     ), //o
    .io_ctrl_tx_payload_last               (ohci_io_phy_tx_payload_last              ), //i
    .io_ctrl_tx_payload_fragment           (ohci_io_phy_tx_payload_fragment[7:0]     ), //i
    .io_ctrl_txEop                         (phy_io_ctrl_txEop                        ), //o
    .io_ctrl_rx_flow_valid                 (phy_io_ctrl_rx_flow_valid                ), //o
    .io_ctrl_rx_flow_payload_stuffingError (phy_io_ctrl_rx_flow_payload_stuffingError), //o
    .io_ctrl_rx_flow_payload_data          (phy_io_ctrl_rx_flow_payload_data[7:0]    ), //o
    .io_ctrl_rx_active                     (phy_io_ctrl_rx_active                    ), //o
    .io_ctrl_usbReset                      (ohci_io_phy_usbReset                     ), //i
    .io_ctrl_usbResume                     (ohci_io_phy_usbResume                    ), //i
    .io_ctrl_overcurrent                   (phy_io_ctrl_overcurrent                  ), //o
    .io_ctrl_tick                          (phy_io_ctrl_tick                         ), //o
    .io_ctrl_ports_0_disable_valid         (ohci_io_phy_ports_0_disable_valid        ), //i
    .io_ctrl_ports_0_disable_ready         (phy_io_ctrl_ports_0_disable_ready        ), //o
    .io_ctrl_ports_0_removable             (ohci_io_phy_ports_0_removable            ), //i
    .io_ctrl_ports_0_power                 (ohci_io_phy_ports_0_power                ), //i
    .io_ctrl_ports_0_reset_valid           (ohci_io_phy_ports_0_reset_valid          ), //i
    .io_ctrl_ports_0_reset_ready           (phy_io_ctrl_ports_0_reset_ready          ), //o
    .io_ctrl_ports_0_suspend_valid         (ohci_io_phy_ports_0_suspend_valid        ), //i
    .io_ctrl_ports_0_suspend_ready         (phy_io_ctrl_ports_0_suspend_ready        ), //o
    .io_ctrl_ports_0_resume_valid          (ohci_io_phy_ports_0_resume_valid         ), //i
    .io_ctrl_ports_0_resume_ready          (phy_io_ctrl_ports_0_resume_ready         ), //o
    .io_ctrl_ports_0_connect               (phy_io_ctrl_ports_0_connect              ), //o
    .io_ctrl_ports_0_disconnect            (phy_io_ctrl_ports_0_disconnect           ), //o
    .io_ctrl_ports_0_overcurrent           (phy_io_ctrl_ports_0_overcurrent          ), //o
    .io_ctrl_ports_0_remoteResume          (phy_io_ctrl_ports_0_remoteResume         ), //o
    .io_ctrl_ports_0_lowSpeed              (phy_io_ctrl_ports_0_lowSpeed             ), //o
    .io_ctrl_ports_1_disable_valid         (ohci_io_phy_ports_1_disable_valid        ), //i
    .io_ctrl_ports_1_disable_ready         (phy_io_ctrl_ports_1_disable_ready        ), //o
    .io_ctrl_ports_1_removable             (ohci_io_phy_ports_1_removable            ), //i
    .io_ctrl_ports_1_power                 (ohci_io_phy_ports_1_power                ), //i
    .io_ctrl_ports_1_reset_valid           (ohci_io_phy_ports_1_reset_valid          ), //i
    .io_ctrl_ports_1_reset_ready           (phy_io_ctrl_ports_1_reset_ready          ), //o
    .io_ctrl_ports_1_suspend_valid         (ohci_io_phy_ports_1_suspend_valid        ), //i
    .io_ctrl_ports_1_suspend_ready         (phy_io_ctrl_ports_1_suspend_ready        ), //o
    .io_ctrl_ports_1_resume_valid          (ohci_io_phy_ports_1_resume_valid         ), //i
    .io_ctrl_ports_1_resume_ready          (phy_io_ctrl_ports_1_resume_ready         ), //o
    .io_ctrl_ports_1_connect               (phy_io_ctrl_ports_1_connect              ), //o
    .io_ctrl_ports_1_disconnect            (phy_io_ctrl_ports_1_disconnect           ), //o
    .io_ctrl_ports_1_overcurrent           (phy_io_ctrl_ports_1_overcurrent          ), //o
    .io_ctrl_ports_1_remoteResume          (phy_io_ctrl_ports_1_remoteResume         ), //o
    .io_ctrl_ports_1_lowSpeed              (phy_io_ctrl_ports_1_lowSpeed             ), //o
    .io_usb_0_tx_enable                    (phy_io_usb_0_tx_enable                   ), //o
    .io_usb_0_tx_data                      (phy_io_usb_0_tx_data                     ), //o
    .io_usb_0_tx_se0                       (phy_io_usb_0_tx_se0                      ), //o
    .io_usb_0_rx_dp                        (usb1_tri_dp_read                         ), //i
    .io_usb_0_rx_dm                        (usb1_tri_dm_read                         ), //i
    .io_usb_1_tx_enable                    (phy_io_usb_1_tx_enable                   ), //o
    .io_usb_1_tx_data                      (phy_io_usb_1_tx_data                     ), //o
    .io_usb_1_tx_se0                       (phy_io_usb_1_tx_se0                      ), //o
    .io_usb_1_rx_dp                        (usb2_tri_dp_read                         ), //i
    .io_usb_1_rx_dm                        (usb2_tri_dm_read                         ), //i
    .io_management_0_overcurrent           (1'b0                                     ), //i
    .io_management_0_power                 (phy_io_management_0_power                ), //o
    .io_management_1_overcurrent           (1'b0                                     ), //i
    .io_management_1_power                 (phy_io_management_1_power                ), //o
    .clk_peripheral                        (clk_peripheral                           ), //i
    .reset_peripheral                      (reset_peripheral                         )  //i
  );
  BmbOnChipRamMultiPort ram_1 (
    .io_buses_0_cmd_valid                    (ohci_io_dma_cmd_valid                              ), //i
    .io_buses_0_cmd_ready                    (ram_1_io_buses_0_cmd_ready                         ), //o
    .io_buses_0_cmd_payload_last             (ohci_io_dma_cmd_payload_last                       ), //i
    .io_buses_0_cmd_payload_fragment_opcode  (ohci_io_dma_cmd_payload_fragment_opcode            ), //i
    .io_buses_0_cmd_payload_fragment_address (ram_1_io_buses_0_cmd_payload_fragment_address[11:0]), //i
    .io_buses_0_cmd_payload_fragment_length  (ohci_io_dma_cmd_payload_fragment_length[5:0]       ), //i
    .io_buses_0_cmd_payload_fragment_data    (ohci_io_dma_cmd_payload_fragment_data[31:0]        ), //i
    .io_buses_0_cmd_payload_fragment_mask    (ohci_io_dma_cmd_payload_fragment_mask[3:0]         ), //i
    .io_buses_0_rsp_valid                    (ram_1_io_buses_0_rsp_valid                         ), //o
    .io_buses_0_rsp_ready                    (ohci_io_dma_rsp_ready                              ), //i
    .io_buses_0_rsp_payload_last             (ram_1_io_buses_0_rsp_payload_last                  ), //o
    .io_buses_0_rsp_payload_fragment_opcode  (ram_1_io_buses_0_rsp_payload_fragment_opcode       ), //o
    .io_buses_0_rsp_payload_fragment_data    (ram_1_io_buses_0_rsp_payload_fragment_data[31:0]   ), //o
    .io_buses_1_cmd_valid                    (ram_1_io_buses_1_cmd_valid                         ), //i
    .io_buses_1_cmd_ready                    (ram_1_io_buses_1_cmd_ready                         ), //o
    .io_buses_1_cmd_payload_last             (1'b1                                               ), //i
    .io_buses_1_cmd_payload_fragment_opcode  (ram_1_io_buses_1_cmd_payload_fragment_opcode       ), //i
    .io_buses_1_cmd_payload_fragment_address (io_apb_dma_PADDR[11:0]                             ), //i
    .io_buses_1_cmd_payload_fragment_length  (2'b11                                              ), //i
    .io_buses_1_cmd_payload_fragment_data    (io_apb_dma_PWDATA[31:0]                            ), //i
    .io_buses_1_cmd_payload_fragment_mask    (4'b1111                                            ), //i
    .io_buses_1_rsp_valid                    (ram_1_io_buses_1_rsp_valid                         ), //o
    .io_buses_1_rsp_ready                    (1'b1                                               ), //i
    .io_buses_1_rsp_payload_last             (ram_1_io_buses_1_rsp_payload_last                  ), //o
    .io_buses_1_rsp_payload_fragment_opcode  (ram_1_io_buses_1_rsp_payload_fragment_opcode       ), //o
    .io_buses_1_rsp_payload_fragment_data    (ram_1_io_buses_1_rsp_payload_fragment_data[31:0]   ), //o
    .clk_peripheral                          (clk_peripheral                                     ), //i
    .reset_peripheral                        (reset_peripheral                                   )  //i
  );
  assign io_usb1_dp = _zz_io_usb1_dp ? usb1_tri_dp_write : 1'bz;
  assign io_usb1_dn = _zz_io_usb1_dn ? usb1_tri_dm_write : 1'bz;
  assign io_usb2_dp = _zz_io_usb2_dp ? usb2_tri_dp_write : 1'bz;
  assign io_usb2_dn = _zz_io_usb2_dn ? usb2_tri_dm_write : 1'bz;
  always @(*) begin
    _zz_io_usb2_dn = 1'b0;
    if(usb2_tri_dm_writeEnable) begin
      _zz_io_usb2_dn = 1'b1;
    end
  end

  always @(*) begin
    _zz_io_usb2_dp = 1'b0;
    if(usb2_tri_dp_writeEnable) begin
      _zz_io_usb2_dp = 1'b1;
    end
  end

  always @(*) begin
    _zz_io_usb1_dn = 1'b0;
    if(usb1_tri_dm_writeEnable) begin
      _zz_io_usb1_dn = 1'b1;
    end
  end

  always @(*) begin
    _zz_io_usb1_dp = 1'b0;
    if(usb1_tri_dp_writeEnable) begin
      _zz_io_usb1_dp = 1'b1;
    end
  end

  assign _zz_io_interrupt = ohci_io_interrupt;
  assign io_interrupt = _zz_io_interrupt;
  assign usb1_tri_dp_writeEnable = phy_io_usb_0_tx_enable;
  assign usb1_tri_dm_writeEnable = phy_io_usb_0_tx_enable;
  assign usb1_tri_dp_write = ((! phy_io_usb_0_tx_se0) && phy_io_usb_0_tx_data);
  assign usb1_tri_dm_write = ((! phy_io_usb_0_tx_se0) && (! phy_io_usb_0_tx_data));
  assign usb1_tri_dp_read = io_usb1_dp;
  assign usb1_tri_dm_read = io_usb1_dn;
  assign usb2_tri_dp_writeEnable = phy_io_usb_1_tx_enable;
  assign usb2_tri_dm_writeEnable = phy_io_usb_1_tx_enable;
  assign usb2_tri_dp_write = ((! phy_io_usb_1_tx_se0) && phy_io_usb_1_tx_data);
  assign usb2_tri_dm_write = ((! phy_io_usb_1_tx_se0) && (! phy_io_usb_1_tx_data));
  assign usb2_tri_dp_read = io_usb2_dp;
  assign usb2_tri_dm_read = io_usb2_dn;
  assign ram_1_io_buses_0_cmd_payload_fragment_address = ohci_io_dma_cmd_payload_fragment_address[11 : 0];
  assign ohci_io_ctrl_cmd_payload_fragment_opcode = io_apb_ctrl_PWRITE;
  assign io_apb_ctrl_PRDATA = ohci_io_ctrl_rsp_payload_fragment_data;
  assign io_apb_ctrl_PREADY = ohci_io_ctrl_rsp_valid;
  assign _zz_when_usb_l96 = (io_apb_ctrl_PSEL[0] && io_apb_ctrl_PENABLE);
  assign when_usb_l96 = (ohci_io_ctrl_cmd_valid && ohci_io_ctrl_cmd_ready);
  assign when_usb_l96_1 = (_zz_when_usb_l96_1 && (! _zz_when_usb_l96));
  assign ohci_io_ctrl_cmd_valid = (_zz_when_usb_l96 && (! _zz_when_usb_l96_1));
  assign ram_1_io_buses_1_cmd_payload_fragment_opcode = io_apb_dma_PWRITE;
  assign io_apb_dma_PRDATA = ram_1_io_buses_1_rsp_payload_fragment_data;
  assign io_apb_dma_PREADY = ram_1_io_buses_1_rsp_valid;
  assign _zz_when_usb_l96_2 = (io_apb_dma_PSEL[0] && io_apb_dma_PENABLE);
  assign when_usb_l96_2 = (ram_1_io_buses_1_cmd_valid && ram_1_io_buses_1_cmd_ready);
  assign when_usb_l96_3 = (_zz_when_usb_l96_3 && (! _zz_when_usb_l96_2));
  assign ram_1_io_buses_1_cmd_valid = (_zz_when_usb_l96_2 && (! _zz_when_usb_l96_3));
  always @(posedge clk_peripheral or posedge reset_peripheral) begin
    if(reset_peripheral) begin
      _zz_when_usb_l96_1 <= 1'b0;
      _zz_when_usb_l96_3 <= 1'b0;
    end else begin
      if(when_usb_l96) begin
        _zz_when_usb_l96_1 <= 1'b1;
      end
      if(when_usb_l96_1) begin
        _zz_when_usb_l96_1 <= 1'b0;
      end
      if(when_usb_l96_2) begin
        _zz_when_usb_l96_3 <= 1'b1;
      end
      if(when_usb_l96_3) begin
        _zz_when_usb_l96_3 <= 1'b0;
      end
    end
  end


endmodule

module StreamArbiter_8 (
  input  wire          io_inputs_0_valid,
  output wire          io_inputs_0_ready,
  input  wire [2:0]    io_inputs_0_payload_opcode,
  input  wire [2:0]    io_inputs_0_payload_param,
  input  wire [2:0]    io_inputs_0_payload_source,
  input  wire [2:0]    io_inputs_0_payload_size,
  input  wire          io_inputs_0_payload_denied,
  input  wire [31:0]   io_inputs_0_payload_data,
  input  wire          io_inputs_0_payload_corrupt,
  input  wire          io_inputs_1_valid,
  output wire          io_inputs_1_ready,
  input  wire [2:0]    io_inputs_1_payload_opcode,
  input  wire [2:0]    io_inputs_1_payload_param,
  input  wire [2:0]    io_inputs_1_payload_source,
  input  wire [2:0]    io_inputs_1_payload_size,
  input  wire          io_inputs_1_payload_denied,
  input  wire [31:0]   io_inputs_1_payload_data,
  input  wire          io_inputs_1_payload_corrupt,
  output wire          io_output_valid,
  input  wire          io_output_ready,
  output wire [2:0]    io_output_payload_opcode,
  output wire [2:0]    io_output_payload_param,
  output wire [2:0]    io_output_payload_source,
  output wire [2:0]    io_output_payload_size,
  output wire          io_output_payload_denied,
  output wire [31:0]   io_output_payload_data,
  output wire          io_output_payload_corrupt,
  output wire [0:0]    io_chosen,
  output wire [1:0]    io_chosenOH,
  input  wire          clk_cpu,
  input  wire          reset_cpu
);
  localparam D_ACCESS_ACK = 3'd0;
  localparam D_ACCESS_ACK_DATA = 3'd1;
  localparam D_GRANT = 3'd4;
  localparam D_GRANT_DATA = 3'd5;
  localparam D_RELEASE_ACK = 3'd6;

  wire       [3:0]    _zz__zz_maskProposal_0_2;
  wire       [3:0]    _zz__zz_maskProposal_0_2_1;
  wire       [1:0]    _zz__zz_maskProposal_0_2_2;
  reg        [3:0]    _zz_io_output_tracker_last;
  reg                 locked;
  wire                maskProposal_0;
  wire                maskProposal_1;
  reg                 maskLocked_0;
  reg                 maskLocked_1;
  wire                maskRouted_0;
  wire                maskRouted_1;
  wire       [1:0]    _zz_maskProposal_0;
  wire       [3:0]    _zz_maskProposal_0_1;
  wire       [3:0]    _zz_maskProposal_0_2;
  wire       [1:0]    _zz_maskProposal_0_3;
  wire                io_output_fire;
  reg        [3:0]    io_output_tracker_beat;
  wire                io_output_tracker_last;
  wire                when_Stream_l794;
  wire       [2:0]    _zz_io_output_payload_opcode;
  wire                _zz_io_chosen;
  `ifndef SYNTHESIS
  reg [119:0] io_inputs_0_payload_opcode_string;
  reg [119:0] io_inputs_1_payload_opcode_string;
  reg [119:0] io_output_payload_opcode_string;
  reg [119:0] _zz_io_output_payload_opcode_string;
  `endif


  assign _zz__zz_maskProposal_0_2 = (_zz_maskProposal_0_1 - _zz__zz_maskProposal_0_2_1);
  assign _zz__zz_maskProposal_0_2_2 = {maskLocked_0,maskLocked_1};
  assign _zz__zz_maskProposal_0_2_1 = {2'd0, _zz__zz_maskProposal_0_2_2};
  always @(*) begin
    case(io_output_payload_size)
      3'b000 : _zz_io_output_tracker_last = 4'b0000;
      3'b001 : _zz_io_output_tracker_last = 4'b0000;
      3'b010 : _zz_io_output_tracker_last = 4'b0000;
      3'b011 : _zz_io_output_tracker_last = 4'b0001;
      3'b100 : _zz_io_output_tracker_last = 4'b0011;
      3'b101 : _zz_io_output_tracker_last = 4'b0111;
      default : _zz_io_output_tracker_last = 4'b1111;
    endcase
  end

  `ifndef SYNTHESIS
  always @(*) begin
    case(io_inputs_0_payload_opcode)
      D_ACCESS_ACK : io_inputs_0_payload_opcode_string = "ACCESS_ACK     ";
      D_ACCESS_ACK_DATA : io_inputs_0_payload_opcode_string = "ACCESS_ACK_DATA";
      D_GRANT : io_inputs_0_payload_opcode_string = "GRANT          ";
      D_GRANT_DATA : io_inputs_0_payload_opcode_string = "GRANT_DATA     ";
      D_RELEASE_ACK : io_inputs_0_payload_opcode_string = "RELEASE_ACK    ";
      default : io_inputs_0_payload_opcode_string = "???????????????";
    endcase
  end
  always @(*) begin
    case(io_inputs_1_payload_opcode)
      D_ACCESS_ACK : io_inputs_1_payload_opcode_string = "ACCESS_ACK     ";
      D_ACCESS_ACK_DATA : io_inputs_1_payload_opcode_string = "ACCESS_ACK_DATA";
      D_GRANT : io_inputs_1_payload_opcode_string = "GRANT          ";
      D_GRANT_DATA : io_inputs_1_payload_opcode_string = "GRANT_DATA     ";
      D_RELEASE_ACK : io_inputs_1_payload_opcode_string = "RELEASE_ACK    ";
      default : io_inputs_1_payload_opcode_string = "???????????????";
    endcase
  end
  always @(*) begin
    case(io_output_payload_opcode)
      D_ACCESS_ACK : io_output_payload_opcode_string = "ACCESS_ACK     ";
      D_ACCESS_ACK_DATA : io_output_payload_opcode_string = "ACCESS_ACK_DATA";
      D_GRANT : io_output_payload_opcode_string = "GRANT          ";
      D_GRANT_DATA : io_output_payload_opcode_string = "GRANT_DATA     ";
      D_RELEASE_ACK : io_output_payload_opcode_string = "RELEASE_ACK    ";
      default : io_output_payload_opcode_string = "???????????????";
    endcase
  end
  always @(*) begin
    case(_zz_io_output_payload_opcode)
      D_ACCESS_ACK : _zz_io_output_payload_opcode_string = "ACCESS_ACK     ";
      D_ACCESS_ACK_DATA : _zz_io_output_payload_opcode_string = "ACCESS_ACK_DATA";
      D_GRANT : _zz_io_output_payload_opcode_string = "GRANT          ";
      D_GRANT_DATA : _zz_io_output_payload_opcode_string = "GRANT_DATA     ";
      D_RELEASE_ACK : _zz_io_output_payload_opcode_string = "RELEASE_ACK    ";
      default : _zz_io_output_payload_opcode_string = "???????????????";
    endcase
  end
  `endif

  assign maskRouted_0 = (locked ? maskLocked_0 : maskProposal_0);
  assign maskRouted_1 = (locked ? maskLocked_1 : maskProposal_1);
  assign _zz_maskProposal_0 = {io_inputs_1_valid,io_inputs_0_valid};
  assign _zz_maskProposal_0_1 = {_zz_maskProposal_0,_zz_maskProposal_0};
  assign _zz_maskProposal_0_2 = (_zz_maskProposal_0_1 & (~ _zz__zz_maskProposal_0_2));
  assign _zz_maskProposal_0_3 = (_zz_maskProposal_0_2[3 : 2] | _zz_maskProposal_0_2[1 : 0]);
  assign maskProposal_0 = _zz_maskProposal_0_3[0];
  assign maskProposal_1 = _zz_maskProposal_0_3[1];
  assign io_output_fire = (io_output_valid && io_output_ready);
  assign io_output_tracker_last = ((! ((1'b0 || (D_ACCESS_ACK_DATA == io_output_payload_opcode)) || (D_GRANT_DATA == io_output_payload_opcode))) || (io_output_tracker_beat == _zz_io_output_tracker_last));
  assign when_Stream_l794 = (io_output_fire && io_output_tracker_last);
  assign io_output_valid = ((io_inputs_0_valid && maskRouted_0) || (io_inputs_1_valid && maskRouted_1));
  assign _zz_io_output_payload_opcode = (maskRouted_0 ? io_inputs_0_payload_opcode : io_inputs_1_payload_opcode);
  assign io_output_payload_opcode = _zz_io_output_payload_opcode;
  assign io_output_payload_param = (maskRouted_0 ? io_inputs_0_payload_param : io_inputs_1_payload_param);
  assign io_output_payload_source = (maskRouted_0 ? io_inputs_0_payload_source : io_inputs_1_payload_source);
  assign io_output_payload_size = (maskRouted_0 ? io_inputs_0_payload_size : io_inputs_1_payload_size);
  assign io_output_payload_denied = (maskRouted_0 ? io_inputs_0_payload_denied : io_inputs_1_payload_denied);
  assign io_output_payload_data = (maskRouted_0 ? io_inputs_0_payload_data : io_inputs_1_payload_data);
  assign io_output_payload_corrupt = (maskRouted_0 ? io_inputs_0_payload_corrupt : io_inputs_1_payload_corrupt);
  assign io_inputs_0_ready = (maskRouted_0 && io_output_ready);
  assign io_inputs_1_ready = (maskRouted_1 && io_output_ready);
  assign io_chosenOH = {maskRouted_1,maskRouted_0};
  assign _zz_io_chosen = io_chosenOH[1];
  assign io_chosen = _zz_io_chosen;
  always @(posedge clk_cpu or posedge reset_cpu) begin
    if(reset_cpu) begin
      locked <= 1'b0;
      maskLocked_0 <= 1'b0;
      maskLocked_1 <= 1'b1;
      io_output_tracker_beat <= 4'b0000;
    end else begin
      if(io_output_valid) begin
        maskLocked_0 <= maskRouted_0;
        maskLocked_1 <= maskRouted_1;
      end
      if(io_output_valid) begin
        locked <= 1'b1;
      end
      if(io_output_fire) begin
        io_output_tracker_beat <= (io_output_tracker_beat + 4'b0001);
        if(io_output_tracker_last) begin
          io_output_tracker_beat <= 4'b0000;
        end
      end
      if(when_Stream_l794) begin
        locked <= 1'b0;
      end
    end
  end


endmodule

module StreamArbiter_7 (
  input  wire          io_inputs_0_valid,
  output wire          io_inputs_0_ready,
  input  wire [2:0]    io_inputs_0_payload_opcode,
  input  wire [2:0]    io_inputs_0_payload_param,
  input  wire [2:0]    io_inputs_0_payload_source,
  input  wire [2:0]    io_inputs_0_payload_size,
  input  wire          io_inputs_0_payload_denied,
  input  wire [63:0]   io_inputs_0_payload_data,
  input  wire          io_inputs_0_payload_corrupt,
  input  wire          io_inputs_1_valid,
  output wire          io_inputs_1_ready,
  input  wire [2:0]    io_inputs_1_payload_opcode,
  input  wire [2:0]    io_inputs_1_payload_param,
  input  wire [2:0]    io_inputs_1_payload_source,
  input  wire [2:0]    io_inputs_1_payload_size,
  input  wire          io_inputs_1_payload_denied,
  input  wire [63:0]   io_inputs_1_payload_data,
  input  wire          io_inputs_1_payload_corrupt,
  output wire          io_output_valid,
  input  wire          io_output_ready,
  output wire [2:0]    io_output_payload_opcode,
  output wire [2:0]    io_output_payload_param,
  output wire [2:0]    io_output_payload_source,
  output wire [2:0]    io_output_payload_size,
  output wire          io_output_payload_denied,
  output wire [63:0]   io_output_payload_data,
  output wire          io_output_payload_corrupt,
  output wire [0:0]    io_chosen,
  output wire [1:0]    io_chosenOH,
  input  wire          clk_cpu,
  input  wire          reset_cpu
);
  localparam D_ACCESS_ACK = 3'd0;
  localparam D_ACCESS_ACK_DATA = 3'd1;
  localparam D_GRANT = 3'd4;
  localparam D_GRANT_DATA = 3'd5;
  localparam D_RELEASE_ACK = 3'd6;

  wire       [3:0]    _zz__zz_maskProposal_0_2;
  wire       [3:0]    _zz__zz_maskProposal_0_2_1;
  wire       [1:0]    _zz__zz_maskProposal_0_2_2;
  reg        [2:0]    _zz_io_output_tracker_last;
  reg                 locked;
  wire                maskProposal_0;
  wire                maskProposal_1;
  reg                 maskLocked_0;
  reg                 maskLocked_1;
  wire                maskRouted_0;
  wire                maskRouted_1;
  wire       [1:0]    _zz_maskProposal_0;
  wire       [3:0]    _zz_maskProposal_0_1;
  wire       [3:0]    _zz_maskProposal_0_2;
  wire       [1:0]    _zz_maskProposal_0_3;
  wire                io_output_fire;
  reg        [2:0]    io_output_tracker_beat;
  wire                io_output_tracker_last;
  wire                when_Stream_l794;
  wire       [2:0]    _zz_io_output_payload_opcode;
  wire                _zz_io_chosen;
  `ifndef SYNTHESIS
  reg [119:0] io_inputs_0_payload_opcode_string;
  reg [119:0] io_inputs_1_payload_opcode_string;
  reg [119:0] io_output_payload_opcode_string;
  reg [119:0] _zz_io_output_payload_opcode_string;
  `endif


  assign _zz__zz_maskProposal_0_2 = (_zz_maskProposal_0_1 - _zz__zz_maskProposal_0_2_1);
  assign _zz__zz_maskProposal_0_2_2 = {maskLocked_0,maskLocked_1};
  assign _zz__zz_maskProposal_0_2_1 = {2'd0, _zz__zz_maskProposal_0_2_2};
  always @(*) begin
    case(io_output_payload_size)
      3'b000 : _zz_io_output_tracker_last = 3'b000;
      3'b001 : _zz_io_output_tracker_last = 3'b000;
      3'b010 : _zz_io_output_tracker_last = 3'b000;
      3'b011 : _zz_io_output_tracker_last = 3'b000;
      3'b100 : _zz_io_output_tracker_last = 3'b001;
      3'b101 : _zz_io_output_tracker_last = 3'b011;
      default : _zz_io_output_tracker_last = 3'b111;
    endcase
  end

  `ifndef SYNTHESIS
  always @(*) begin
    case(io_inputs_0_payload_opcode)
      D_ACCESS_ACK : io_inputs_0_payload_opcode_string = "ACCESS_ACK     ";
      D_ACCESS_ACK_DATA : io_inputs_0_payload_opcode_string = "ACCESS_ACK_DATA";
      D_GRANT : io_inputs_0_payload_opcode_string = "GRANT          ";
      D_GRANT_DATA : io_inputs_0_payload_opcode_string = "GRANT_DATA     ";
      D_RELEASE_ACK : io_inputs_0_payload_opcode_string = "RELEASE_ACK    ";
      default : io_inputs_0_payload_opcode_string = "???????????????";
    endcase
  end
  always @(*) begin
    case(io_inputs_1_payload_opcode)
      D_ACCESS_ACK : io_inputs_1_payload_opcode_string = "ACCESS_ACK     ";
      D_ACCESS_ACK_DATA : io_inputs_1_payload_opcode_string = "ACCESS_ACK_DATA";
      D_GRANT : io_inputs_1_payload_opcode_string = "GRANT          ";
      D_GRANT_DATA : io_inputs_1_payload_opcode_string = "GRANT_DATA     ";
      D_RELEASE_ACK : io_inputs_1_payload_opcode_string = "RELEASE_ACK    ";
      default : io_inputs_1_payload_opcode_string = "???????????????";
    endcase
  end
  always @(*) begin
    case(io_output_payload_opcode)
      D_ACCESS_ACK : io_output_payload_opcode_string = "ACCESS_ACK     ";
      D_ACCESS_ACK_DATA : io_output_payload_opcode_string = "ACCESS_ACK_DATA";
      D_GRANT : io_output_payload_opcode_string = "GRANT          ";
      D_GRANT_DATA : io_output_payload_opcode_string = "GRANT_DATA     ";
      D_RELEASE_ACK : io_output_payload_opcode_string = "RELEASE_ACK    ";
      default : io_output_payload_opcode_string = "???????????????";
    endcase
  end
  always @(*) begin
    case(_zz_io_output_payload_opcode)
      D_ACCESS_ACK : _zz_io_output_payload_opcode_string = "ACCESS_ACK     ";
      D_ACCESS_ACK_DATA : _zz_io_output_payload_opcode_string = "ACCESS_ACK_DATA";
      D_GRANT : _zz_io_output_payload_opcode_string = "GRANT          ";
      D_GRANT_DATA : _zz_io_output_payload_opcode_string = "GRANT_DATA     ";
      D_RELEASE_ACK : _zz_io_output_payload_opcode_string = "RELEASE_ACK    ";
      default : _zz_io_output_payload_opcode_string = "???????????????";
    endcase
  end
  `endif

  assign maskRouted_0 = (locked ? maskLocked_0 : maskProposal_0);
  assign maskRouted_1 = (locked ? maskLocked_1 : maskProposal_1);
  assign _zz_maskProposal_0 = {io_inputs_1_valid,io_inputs_0_valid};
  assign _zz_maskProposal_0_1 = {_zz_maskProposal_0,_zz_maskProposal_0};
  assign _zz_maskProposal_0_2 = (_zz_maskProposal_0_1 & (~ _zz__zz_maskProposal_0_2));
  assign _zz_maskProposal_0_3 = (_zz_maskProposal_0_2[3 : 2] | _zz_maskProposal_0_2[1 : 0]);
  assign maskProposal_0 = _zz_maskProposal_0_3[0];
  assign maskProposal_1 = _zz_maskProposal_0_3[1];
  assign io_output_fire = (io_output_valid && io_output_ready);
  assign io_output_tracker_last = ((! ((1'b0 || (D_ACCESS_ACK_DATA == io_output_payload_opcode)) || (D_GRANT_DATA == io_output_payload_opcode))) || (io_output_tracker_beat == _zz_io_output_tracker_last));
  assign when_Stream_l794 = (io_output_fire && io_output_tracker_last);
  assign io_output_valid = ((io_inputs_0_valid && maskRouted_0) || (io_inputs_1_valid && maskRouted_1));
  assign _zz_io_output_payload_opcode = (maskRouted_0 ? io_inputs_0_payload_opcode : io_inputs_1_payload_opcode);
  assign io_output_payload_opcode = _zz_io_output_payload_opcode;
  assign io_output_payload_param = (maskRouted_0 ? io_inputs_0_payload_param : io_inputs_1_payload_param);
  assign io_output_payload_source = (maskRouted_0 ? io_inputs_0_payload_source : io_inputs_1_payload_source);
  assign io_output_payload_size = (maskRouted_0 ? io_inputs_0_payload_size : io_inputs_1_payload_size);
  assign io_output_payload_denied = (maskRouted_0 ? io_inputs_0_payload_denied : io_inputs_1_payload_denied);
  assign io_output_payload_data = (maskRouted_0 ? io_inputs_0_payload_data : io_inputs_1_payload_data);
  assign io_output_payload_corrupt = (maskRouted_0 ? io_inputs_0_payload_corrupt : io_inputs_1_payload_corrupt);
  assign io_inputs_0_ready = (maskRouted_0 && io_output_ready);
  assign io_inputs_1_ready = (maskRouted_1 && io_output_ready);
  assign io_chosenOH = {maskRouted_1,maskRouted_0};
  assign _zz_io_chosen = io_chosenOH[1];
  assign io_chosen = _zz_io_chosen;
  always @(posedge clk_cpu or posedge reset_cpu) begin
    if(reset_cpu) begin
      locked <= 1'b0;
      maskLocked_0 <= 1'b0;
      maskLocked_1 <= 1'b1;
      io_output_tracker_beat <= 3'b000;
    end else begin
      if(io_output_valid) begin
        maskLocked_0 <= maskRouted_0;
        maskLocked_1 <= maskRouted_1;
      end
      if(io_output_valid) begin
        locked <= 1'b1;
      end
      if(io_output_fire) begin
        io_output_tracker_beat <= (io_output_tracker_beat + 3'b001);
        if(io_output_tracker_last) begin
          io_output_tracker_beat <= 3'b000;
        end
      end
      if(when_Stream_l794) begin
        locked <= 1'b0;
      end
    end
  end


endmodule

module StreamFifoCC_3 (
  input  wire          io_push_valid,
  output wire          io_push_ready,
  input  wire [2:0]    io_push_payload_id,
  input  wire [1:0]    io_push_payload_resp,
  output wire          io_pop_valid,
  input  wire          io_pop_ready,
  output wire [2:0]    io_pop_payload_id,
  output wire [1:0]    io_pop_payload_resp,
  output wire [1:0]    io_pushOccupancy,
  output wire [1:0]    io_popOccupancy,
  input  wire          clk_ram_bus,
  input  wire          reset_ram,
  input  wire          clk_cpu,
  input  wire          ram_axi_cc_toplevel_board_ctrl_reset_ram_synchronized_1
);

  reg        [4:0]    ram_1_spinal_port1;
  wire       [1:0]    popToPushGray_buffercc_io_dataOut;
  wire       [1:0]    pushToPopGray_buffercc_io_dataOut;
  wire       [1:0]    _zz_pushCC_pushPtrGray;
  wire       [0:0]    _zz_ram_1_port;
  wire       [4:0]    _zz_ram_1_port_1;
  wire       [1:0]    _zz_popCC_popPtrGray;
  reg                 _zz_1;
  wire       [1:0]    popToPushGray;
  wire       [1:0]    pushToPopGray;
  reg        [1:0]    pushCC_pushPtr;
  wire       [1:0]    pushCC_pushPtrPlus;
  wire                io_push_fire;
  reg        [1:0]    pushCC_pushPtrGray;
  wire       [1:0]    pushCC_popPtrGray;
  wire                pushCC_full;
  wire                _zz_io_pushOccupancy;
  reg        [1:0]    popCC_popPtr;
  (* keep , syn_keep *) wire       [1:0]    popCC_popPtrPlus /* synthesis syn_keep = 1 */ ;
  wire       [1:0]    popCC_popPtrGray;
  wire       [1:0]    popCC_pushPtrGray;
  wire                popCC_addressGen_valid;
  reg                 popCC_addressGen_ready;
  wire       [0:0]    popCC_addressGen_payload;
  wire                popCC_empty;
  wire                popCC_addressGen_fire;
  wire                popCC_readArbitation_valid;
  wire                popCC_readArbitation_ready;
  wire       [0:0]    popCC_readArbitation_payload;
  reg                 popCC_addressGen_rValid;
  reg        [0:0]    popCC_addressGen_rData;
  wire                when_Stream_l393;
  wire                popCC_readPort_cmd_valid;
  wire       [0:0]    popCC_readPort_cmd_payload;
  wire       [2:0]    popCC_readPort_rsp_id;
  wire       [1:0]    popCC_readPort_rsp_resp;
  wire       [4:0]    _zz_popCC_readPort_rsp_id;
  wire                popCC_readArbitation_translated_valid;
  wire                popCC_readArbitation_translated_ready;
  wire       [2:0]    popCC_readArbitation_translated_payload_id;
  wire       [1:0]    popCC_readArbitation_translated_payload_resp;
  wire                popCC_readArbitation_fire;
  reg        [1:0]    popCC_ptrToPush;
  reg        [1:0]    popCC_ptrToOccupancy;
  wire                _zz_io_popOccupancy;
  reg [4:0] ram_1 [0:1];

  assign _zz_pushCC_pushPtrGray = (pushCC_pushPtrPlus >>> 1'b1);
  assign _zz_ram_1_port = pushCC_pushPtr[0:0];
  assign _zz_popCC_popPtrGray = (popCC_popPtr >>> 1'b1);
  assign _zz_ram_1_port_1 = {io_push_payload_resp,io_push_payload_id};
  always @(posedge clk_ram_bus) begin
    if(_zz_1) begin
      ram_1[_zz_ram_1_port] <= _zz_ram_1_port_1;
    end
  end

  always @(posedge clk_cpu) begin
    if(popCC_readPort_cmd_valid) begin
      ram_1_spinal_port1 <= ram_1[popCC_readPort_cmd_payload];
    end
  end

  (* keep_hierarchy = "TRUE" *) BufferCC_8 popToPushGray_buffercc (
    .io_dataIn   (popToPushGray[1:0]                    ), //i
    .io_dataOut  (popToPushGray_buffercc_io_dataOut[1:0]), //o
    .clk_ram_bus (clk_ram_bus                           ), //i
    .reset_ram   (reset_ram                             )  //i
  );
  (* keep_hierarchy = "TRUE" *) BufferCC_9 pushToPopGray_buffercc (
    .io_dataIn                                               (pushToPopGray[1:0]                                     ), //i
    .io_dataOut                                              (pushToPopGray_buffercc_io_dataOut[1:0]                 ), //o
    .clk_cpu                                                 (clk_cpu                                                ), //i
    .ram_axi_cc_toplevel_board_ctrl_reset_ram_synchronized_1 (ram_axi_cc_toplevel_board_ctrl_reset_ram_synchronized_1)  //i
  );
  always @(*) begin
    _zz_1 = 1'b0;
    if(io_push_fire) begin
      _zz_1 = 1'b1;
    end
  end

  assign pushCC_pushPtrPlus = (pushCC_pushPtr + 2'b01);
  assign io_push_fire = (io_push_valid && io_push_ready);
  assign pushCC_popPtrGray = popToPushGray_buffercc_io_dataOut;
  assign pushCC_full = ((pushCC_pushPtrGray[1 : 0] == (~ pushCC_popPtrGray[1 : 0])) && 1'b1);
  assign io_push_ready = (! pushCC_full);
  assign _zz_io_pushOccupancy = pushCC_popPtrGray[1];
  assign io_pushOccupancy = (pushCC_pushPtr - {_zz_io_pushOccupancy,(pushCC_popPtrGray[0] ^ _zz_io_pushOccupancy)});
  assign popCC_popPtrPlus = (popCC_popPtr + 2'b01);
  assign popCC_popPtrGray = (_zz_popCC_popPtrGray ^ popCC_popPtr);
  assign popCC_pushPtrGray = pushToPopGray_buffercc_io_dataOut;
  assign popCC_empty = (popCC_popPtrGray == popCC_pushPtrGray);
  assign popCC_addressGen_valid = (! popCC_empty);
  assign popCC_addressGen_payload = popCC_popPtr[0:0];
  assign popCC_addressGen_fire = (popCC_addressGen_valid && popCC_addressGen_ready);
  always @(*) begin
    popCC_addressGen_ready = popCC_readArbitation_ready;
    if(when_Stream_l393) begin
      popCC_addressGen_ready = 1'b1;
    end
  end

  assign when_Stream_l393 = (! popCC_readArbitation_valid);
  assign popCC_readArbitation_valid = popCC_addressGen_rValid;
  assign popCC_readArbitation_payload = popCC_addressGen_rData;
  assign _zz_popCC_readPort_rsp_id = ram_1_spinal_port1;
  assign popCC_readPort_rsp_id = _zz_popCC_readPort_rsp_id[2 : 0];
  assign popCC_readPort_rsp_resp = _zz_popCC_readPort_rsp_id[4 : 3];
  assign popCC_readPort_cmd_valid = popCC_addressGen_fire;
  assign popCC_readPort_cmd_payload = popCC_addressGen_payload;
  assign popCC_readArbitation_translated_valid = popCC_readArbitation_valid;
  assign popCC_readArbitation_ready = popCC_readArbitation_translated_ready;
  assign popCC_readArbitation_translated_payload_id = popCC_readPort_rsp_id;
  assign popCC_readArbitation_translated_payload_resp = popCC_readPort_rsp_resp;
  assign io_pop_valid = popCC_readArbitation_translated_valid;
  assign popCC_readArbitation_translated_ready = io_pop_ready;
  assign io_pop_payload_id = popCC_readArbitation_translated_payload_id;
  assign io_pop_payload_resp = popCC_readArbitation_translated_payload_resp;
  assign popCC_readArbitation_fire = (popCC_readArbitation_valid && popCC_readArbitation_ready);
  assign _zz_io_popOccupancy = popCC_pushPtrGray[1];
  assign io_popOccupancy = ({_zz_io_popOccupancy,(popCC_pushPtrGray[0] ^ _zz_io_popOccupancy)} - popCC_ptrToOccupancy);
  assign pushToPopGray = pushCC_pushPtrGray;
  assign popToPushGray = popCC_ptrToPush;
  always @(posedge clk_ram_bus or posedge reset_ram) begin
    if(reset_ram) begin
      pushCC_pushPtr <= 2'b00;
      pushCC_pushPtrGray <= 2'b00;
    end else begin
      if(io_push_fire) begin
        pushCC_pushPtrGray <= (_zz_pushCC_pushPtrGray ^ pushCC_pushPtrPlus);
      end
      if(io_push_fire) begin
        pushCC_pushPtr <= pushCC_pushPtrPlus;
      end
    end
  end

  always @(posedge clk_cpu or posedge ram_axi_cc_toplevel_board_ctrl_reset_ram_synchronized_1) begin
    if(ram_axi_cc_toplevel_board_ctrl_reset_ram_synchronized_1) begin
      popCC_popPtr <= 2'b00;
      popCC_addressGen_rValid <= 1'b0;
      popCC_ptrToPush <= 2'b00;
      popCC_ptrToOccupancy <= 2'b00;
    end else begin
      if(popCC_addressGen_fire) begin
        popCC_popPtr <= popCC_popPtrPlus;
      end
      if(popCC_addressGen_ready) begin
        popCC_addressGen_rValid <= popCC_addressGen_valid;
      end
      if(popCC_readArbitation_fire) begin
        popCC_ptrToPush <= popCC_popPtrGray;
      end
      if(popCC_readArbitation_fire) begin
        popCC_ptrToOccupancy <= popCC_popPtr;
      end
    end
  end

  always @(posedge clk_cpu) begin
    if(popCC_addressGen_ready) begin
      popCC_addressGen_rData <= popCC_addressGen_payload;
    end
  end


endmodule

module StreamFifoCC_2 (
  input  wire          io_push_valid,
  output wire          io_push_ready,
  input  wire [63:0]   io_push_payload_data,
  input  wire [7:0]    io_push_payload_strb,
  input  wire          io_push_payload_last,
  output wire          io_pop_valid,
  input  wire          io_pop_ready,
  output wire [63:0]   io_pop_payload_data,
  output wire [7:0]    io_pop_payload_strb,
  output wire          io_pop_payload_last,
  output wire [4:0]    io_pushOccupancy,
  output wire [4:0]    io_popOccupancy,
  input  wire          clk_cpu,
  input  wire          reset_cpu,
  input  wire          clk_ram_bus,
  input  wire          ram_axi_cc_toplevel_board_ctrl_reset_cpu_synchronized_1
);

  reg        [72:0]   ram_1_spinal_port1;
  wire       [4:0]    popToPushGray_buffercc_io_dataOut;
  wire       [4:0]    pushToPopGray_buffercc_io_dataOut;
  wire       [4:0]    _zz_pushCC_pushPtrGray;
  wire       [3:0]    _zz_ram_1_port;
  wire       [72:0]   _zz_ram_1_port_1;
  wire       [4:0]    _zz_popCC_popPtrGray;
  reg                 _zz_1;
  wire       [4:0]    popToPushGray;
  wire       [4:0]    pushToPopGray;
  reg        [4:0]    pushCC_pushPtr;
  wire       [4:0]    pushCC_pushPtrPlus;
  wire                io_push_fire;
  reg        [4:0]    pushCC_pushPtrGray;
  wire       [4:0]    pushCC_popPtrGray;
  wire                pushCC_full;
  wire                _zz_io_pushOccupancy;
  wire                _zz_io_pushOccupancy_1;
  wire                _zz_io_pushOccupancy_2;
  wire                _zz_io_pushOccupancy_3;
  reg        [4:0]    popCC_popPtr;
  (* keep , syn_keep *) wire       [4:0]    popCC_popPtrPlus /* synthesis syn_keep = 1 */ ;
  wire       [4:0]    popCC_popPtrGray;
  wire       [4:0]    popCC_pushPtrGray;
  wire                popCC_addressGen_valid;
  reg                 popCC_addressGen_ready;
  wire       [3:0]    popCC_addressGen_payload;
  wire                popCC_empty;
  wire                popCC_addressGen_fire;
  wire                popCC_readArbitation_valid;
  wire                popCC_readArbitation_ready;
  wire       [3:0]    popCC_readArbitation_payload;
  reg                 popCC_addressGen_rValid;
  reg        [3:0]    popCC_addressGen_rData;
  wire                when_Stream_l393;
  wire                popCC_readPort_cmd_valid;
  wire       [3:0]    popCC_readPort_cmd_payload;
  wire       [63:0]   popCC_readPort_rsp_data;
  wire       [7:0]    popCC_readPort_rsp_strb;
  wire                popCC_readPort_rsp_last;
  wire       [72:0]   _zz_popCC_readPort_rsp_data;
  wire                popCC_readArbitation_translated_valid;
  wire                popCC_readArbitation_translated_ready;
  wire       [63:0]   popCC_readArbitation_translated_payload_data;
  wire       [7:0]    popCC_readArbitation_translated_payload_strb;
  wire                popCC_readArbitation_translated_payload_last;
  wire                popCC_readArbitation_fire;
  reg        [4:0]    popCC_ptrToPush;
  reg        [4:0]    popCC_ptrToOccupancy;
  wire                _zz_io_popOccupancy;
  wire                _zz_io_popOccupancy_1;
  wire                _zz_io_popOccupancy_2;
  wire                _zz_io_popOccupancy_3;
  reg [72:0] ram_1 [0:15];

  assign _zz_pushCC_pushPtrGray = (pushCC_pushPtrPlus >>> 1'b1);
  assign _zz_ram_1_port = pushCC_pushPtr[3:0];
  assign _zz_popCC_popPtrGray = (popCC_popPtr >>> 1'b1);
  assign _zz_ram_1_port_1 = {io_push_payload_last,{io_push_payload_strb,io_push_payload_data}};
  always @(posedge clk_cpu) begin
    if(_zz_1) begin
      ram_1[_zz_ram_1_port] <= _zz_ram_1_port_1;
    end
  end

  always @(posedge clk_ram_bus) begin
    if(popCC_readPort_cmd_valid) begin
      ram_1_spinal_port1 <= ram_1[popCC_readPort_cmd_payload];
    end
  end

  (* keep_hierarchy = "TRUE" *) BufferCC_6 popToPushGray_buffercc (
    .io_dataIn  (popToPushGray[4:0]                    ), //i
    .io_dataOut (popToPushGray_buffercc_io_dataOut[4:0]), //o
    .clk_cpu    (clk_cpu                               ), //i
    .reset_cpu  (reset_cpu                             )  //i
  );
  (* keep_hierarchy = "TRUE" *) BufferCC_7 pushToPopGray_buffercc (
    .io_dataIn                                               (pushToPopGray[4:0]                                     ), //i
    .io_dataOut                                              (pushToPopGray_buffercc_io_dataOut[4:0]                 ), //o
    .clk_ram_bus                                             (clk_ram_bus                                            ), //i
    .ram_axi_cc_toplevel_board_ctrl_reset_cpu_synchronized_1 (ram_axi_cc_toplevel_board_ctrl_reset_cpu_synchronized_1)  //i
  );
  always @(*) begin
    _zz_1 = 1'b0;
    if(io_push_fire) begin
      _zz_1 = 1'b1;
    end
  end

  assign pushCC_pushPtrPlus = (pushCC_pushPtr + 5'h01);
  assign io_push_fire = (io_push_valid && io_push_ready);
  assign pushCC_popPtrGray = popToPushGray_buffercc_io_dataOut;
  assign pushCC_full = ((pushCC_pushPtrGray[4 : 3] == (~ pushCC_popPtrGray[4 : 3])) && (pushCC_pushPtrGray[2 : 0] == pushCC_popPtrGray[2 : 0]));
  assign io_push_ready = (! pushCC_full);
  assign _zz_io_pushOccupancy = (pushCC_popPtrGray[1] ^ _zz_io_pushOccupancy_1);
  assign _zz_io_pushOccupancy_1 = (pushCC_popPtrGray[2] ^ _zz_io_pushOccupancy_2);
  assign _zz_io_pushOccupancy_2 = (pushCC_popPtrGray[3] ^ _zz_io_pushOccupancy_3);
  assign _zz_io_pushOccupancy_3 = pushCC_popPtrGray[4];
  assign io_pushOccupancy = (pushCC_pushPtr - {_zz_io_pushOccupancy_3,{_zz_io_pushOccupancy_2,{_zz_io_pushOccupancy_1,{_zz_io_pushOccupancy,(pushCC_popPtrGray[0] ^ _zz_io_pushOccupancy)}}}});
  assign popCC_popPtrPlus = (popCC_popPtr + 5'h01);
  assign popCC_popPtrGray = (_zz_popCC_popPtrGray ^ popCC_popPtr);
  assign popCC_pushPtrGray = pushToPopGray_buffercc_io_dataOut;
  assign popCC_empty = (popCC_popPtrGray == popCC_pushPtrGray);
  assign popCC_addressGen_valid = (! popCC_empty);
  assign popCC_addressGen_payload = popCC_popPtr[3:0];
  assign popCC_addressGen_fire = (popCC_addressGen_valid && popCC_addressGen_ready);
  always @(*) begin
    popCC_addressGen_ready = popCC_readArbitation_ready;
    if(when_Stream_l393) begin
      popCC_addressGen_ready = 1'b1;
    end
  end

  assign when_Stream_l393 = (! popCC_readArbitation_valid);
  assign popCC_readArbitation_valid = popCC_addressGen_rValid;
  assign popCC_readArbitation_payload = popCC_addressGen_rData;
  assign _zz_popCC_readPort_rsp_data = ram_1_spinal_port1;
  assign popCC_readPort_rsp_data = _zz_popCC_readPort_rsp_data[63 : 0];
  assign popCC_readPort_rsp_strb = _zz_popCC_readPort_rsp_data[71 : 64];
  assign popCC_readPort_rsp_last = _zz_popCC_readPort_rsp_data[72];
  assign popCC_readPort_cmd_valid = popCC_addressGen_fire;
  assign popCC_readPort_cmd_payload = popCC_addressGen_payload;
  assign popCC_readArbitation_translated_valid = popCC_readArbitation_valid;
  assign popCC_readArbitation_ready = popCC_readArbitation_translated_ready;
  assign popCC_readArbitation_translated_payload_data = popCC_readPort_rsp_data;
  assign popCC_readArbitation_translated_payload_strb = popCC_readPort_rsp_strb;
  assign popCC_readArbitation_translated_payload_last = popCC_readPort_rsp_last;
  assign io_pop_valid = popCC_readArbitation_translated_valid;
  assign popCC_readArbitation_translated_ready = io_pop_ready;
  assign io_pop_payload_data = popCC_readArbitation_translated_payload_data;
  assign io_pop_payload_strb = popCC_readArbitation_translated_payload_strb;
  assign io_pop_payload_last = popCC_readArbitation_translated_payload_last;
  assign popCC_readArbitation_fire = (popCC_readArbitation_valid && popCC_readArbitation_ready);
  assign _zz_io_popOccupancy = (popCC_pushPtrGray[1] ^ _zz_io_popOccupancy_1);
  assign _zz_io_popOccupancy_1 = (popCC_pushPtrGray[2] ^ _zz_io_popOccupancy_2);
  assign _zz_io_popOccupancy_2 = (popCC_pushPtrGray[3] ^ _zz_io_popOccupancy_3);
  assign _zz_io_popOccupancy_3 = popCC_pushPtrGray[4];
  assign io_popOccupancy = ({_zz_io_popOccupancy_3,{_zz_io_popOccupancy_2,{_zz_io_popOccupancy_1,{_zz_io_popOccupancy,(popCC_pushPtrGray[0] ^ _zz_io_popOccupancy)}}}} - popCC_ptrToOccupancy);
  assign pushToPopGray = pushCC_pushPtrGray;
  assign popToPushGray = popCC_ptrToPush;
  always @(posedge clk_cpu or posedge reset_cpu) begin
    if(reset_cpu) begin
      pushCC_pushPtr <= 5'h0;
      pushCC_pushPtrGray <= 5'h0;
    end else begin
      if(io_push_fire) begin
        pushCC_pushPtrGray <= (_zz_pushCC_pushPtrGray ^ pushCC_pushPtrPlus);
      end
      if(io_push_fire) begin
        pushCC_pushPtr <= pushCC_pushPtrPlus;
      end
    end
  end

  always @(posedge clk_ram_bus or posedge ram_axi_cc_toplevel_board_ctrl_reset_cpu_synchronized_1) begin
    if(ram_axi_cc_toplevel_board_ctrl_reset_cpu_synchronized_1) begin
      popCC_popPtr <= 5'h0;
      popCC_addressGen_rValid <= 1'b0;
      popCC_ptrToPush <= 5'h0;
      popCC_ptrToOccupancy <= 5'h0;
    end else begin
      if(popCC_addressGen_fire) begin
        popCC_popPtr <= popCC_popPtrPlus;
      end
      if(popCC_addressGen_ready) begin
        popCC_addressGen_rValid <= popCC_addressGen_valid;
      end
      if(popCC_readArbitation_fire) begin
        popCC_ptrToPush <= popCC_popPtrGray;
      end
      if(popCC_readArbitation_fire) begin
        popCC_ptrToOccupancy <= popCC_popPtr;
      end
    end
  end

  always @(posedge clk_ram_bus) begin
    if(popCC_addressGen_ready) begin
      popCC_addressGen_rData <= popCC_addressGen_payload;
    end
  end


endmodule

module StreamFifoCC_1 (
  input  wire          io_push_valid,
  output wire          io_push_ready,
  input  wire [63:0]   io_push_payload_data,
  input  wire [2:0]    io_push_payload_id,
  input  wire [1:0]    io_push_payload_resp,
  input  wire          io_push_payload_last,
  output wire          io_pop_valid,
  input  wire          io_pop_ready,
  output wire [63:0]   io_pop_payload_data,
  output wire [2:0]    io_pop_payload_id,
  output wire [1:0]    io_pop_payload_resp,
  output wire          io_pop_payload_last,
  output wire [7:0]    io_pushOccupancy,
  output wire [7:0]    io_popOccupancy,
  input  wire          clk_ram_bus,
  input  wire          reset_ram,
  input  wire          clk_cpu,
  output wire          ram_axi_cc_toplevel_board_ctrl_reset_ram_synchronized_1
);

  reg        [69:0]   ram_1_spinal_port1;
  wire       [7:0]    popToPushGray_buffercc_io_dataOut;
  wire                ram_axi_cc_toplevel_board_ctrl_reset_ram_asyncAssertSyncDeassert_buffercc_io_dataOut;
  wire       [7:0]    pushToPopGray_buffercc_io_dataOut;
  wire       [7:0]    _zz_pushCC_pushPtrGray;
  wire       [6:0]    _zz_ram_1_port;
  wire       [69:0]   _zz_ram_1_port_1;
  wire       [7:0]    _zz_popCC_popPtrGray;
  reg                 _zz_1;
  wire       [7:0]    popToPushGray;
  wire       [7:0]    pushToPopGray;
  reg        [7:0]    pushCC_pushPtr;
  wire       [7:0]    pushCC_pushPtrPlus;
  wire                io_push_fire;
  reg        [7:0]    pushCC_pushPtrGray;
  wire       [7:0]    pushCC_popPtrGray;
  wire                pushCC_full;
  wire                _zz_io_pushOccupancy;
  wire                _zz_io_pushOccupancy_1;
  wire                _zz_io_pushOccupancy_2;
  wire                _zz_io_pushOccupancy_3;
  wire                _zz_io_pushOccupancy_4;
  wire                _zz_io_pushOccupancy_5;
  wire                _zz_io_pushOccupancy_6;
  wire                ram_axi_cc_toplevel_board_ctrl_reset_ram_asyncAssertSyncDeassert;
  wire                ram_axi_cc_toplevel_board_ctrl_reset_ram_synchronized;
  reg        [7:0]    popCC_popPtr;
  (* keep , syn_keep *) wire       [7:0]    popCC_popPtrPlus /* synthesis syn_keep = 1 */ ;
  wire       [7:0]    popCC_popPtrGray;
  wire       [7:0]    popCC_pushPtrGray;
  wire                popCC_addressGen_valid;
  reg                 popCC_addressGen_ready;
  wire       [6:0]    popCC_addressGen_payload;
  wire                popCC_empty;
  wire                popCC_addressGen_fire;
  wire                popCC_readArbitation_valid;
  wire                popCC_readArbitation_ready;
  wire       [6:0]    popCC_readArbitation_payload;
  reg                 popCC_addressGen_rValid;
  reg        [6:0]    popCC_addressGen_rData;
  wire                when_Stream_l393;
  wire                popCC_readPort_cmd_valid;
  wire       [6:0]    popCC_readPort_cmd_payload;
  wire       [63:0]   popCC_readPort_rsp_data;
  wire       [2:0]    popCC_readPort_rsp_id;
  wire       [1:0]    popCC_readPort_rsp_resp;
  wire                popCC_readPort_rsp_last;
  wire       [69:0]   _zz_popCC_readPort_rsp_data;
  wire                popCC_readArbitation_translated_valid;
  wire                popCC_readArbitation_translated_ready;
  wire       [63:0]   popCC_readArbitation_translated_payload_data;
  wire       [2:0]    popCC_readArbitation_translated_payload_id;
  wire       [1:0]    popCC_readArbitation_translated_payload_resp;
  wire                popCC_readArbitation_translated_payload_last;
  wire                popCC_readArbitation_fire;
  reg        [7:0]    popCC_ptrToPush;
  reg        [7:0]    popCC_ptrToOccupancy;
  wire                _zz_io_popOccupancy;
  wire                _zz_io_popOccupancy_1;
  wire                _zz_io_popOccupancy_2;
  wire                _zz_io_popOccupancy_3;
  wire                _zz_io_popOccupancy_4;
  wire                _zz_io_popOccupancy_5;
  wire                _zz_io_popOccupancy_6;
  reg [69:0] ram_1 [0:127];

  assign _zz_pushCC_pushPtrGray = (pushCC_pushPtrPlus >>> 1'b1);
  assign _zz_ram_1_port = pushCC_pushPtr[6:0];
  assign _zz_popCC_popPtrGray = (popCC_popPtr >>> 1'b1);
  assign _zz_ram_1_port_1 = {io_push_payload_last,{io_push_payload_resp,{io_push_payload_id,io_push_payload_data}}};
  always @(posedge clk_ram_bus) begin
    if(_zz_1) begin
      ram_1[_zz_ram_1_port] <= _zz_ram_1_port_1;
    end
  end

  always @(posedge clk_cpu) begin
    if(popCC_readPort_cmd_valid) begin
      ram_1_spinal_port1 <= ram_1[popCC_readPort_cmd_payload];
    end
  end

  (* keep_hierarchy = "TRUE" *) BufferCC_3 popToPushGray_buffercc (
    .io_dataIn   (popToPushGray[7:0]                    ), //i
    .io_dataOut  (popToPushGray_buffercc_io_dataOut[7:0]), //o
    .clk_ram_bus (clk_ram_bus                           ), //i
    .reset_ram   (reset_ram                             )  //i
  );
  (* keep_hierarchy = "TRUE" *) BufferCC_4 ram_axi_cc_toplevel_board_ctrl_reset_ram_asyncAssertSyncDeassert_buffercc (
    .io_dataIn  (ram_axi_cc_toplevel_board_ctrl_reset_ram_asyncAssertSyncDeassert                    ), //i
    .io_dataOut (ram_axi_cc_toplevel_board_ctrl_reset_ram_asyncAssertSyncDeassert_buffercc_io_dataOut), //o
    .clk_cpu    (clk_cpu                                                                             ), //i
    .reset_ram  (reset_ram                                                                           )  //i
  );
  (* keep_hierarchy = "TRUE" *) BufferCC_5 pushToPopGray_buffercc (
    .io_dataIn                                             (pushToPopGray[7:0]                                   ), //i
    .io_dataOut                                            (pushToPopGray_buffercc_io_dataOut[7:0]               ), //o
    .clk_cpu                                               (clk_cpu                                              ), //i
    .ram_axi_cc_toplevel_board_ctrl_reset_ram_synchronized (ram_axi_cc_toplevel_board_ctrl_reset_ram_synchronized)  //i
  );
  always @(*) begin
    _zz_1 = 1'b0;
    if(io_push_fire) begin
      _zz_1 = 1'b1;
    end
  end

  assign pushCC_pushPtrPlus = (pushCC_pushPtr + 8'h01);
  assign io_push_fire = (io_push_valid && io_push_ready);
  assign pushCC_popPtrGray = popToPushGray_buffercc_io_dataOut;
  assign pushCC_full = ((pushCC_pushPtrGray[7 : 6] == (~ pushCC_popPtrGray[7 : 6])) && (pushCC_pushPtrGray[5 : 0] == pushCC_popPtrGray[5 : 0]));
  assign io_push_ready = (! pushCC_full);
  assign _zz_io_pushOccupancy = (pushCC_popPtrGray[1] ^ _zz_io_pushOccupancy_1);
  assign _zz_io_pushOccupancy_1 = (pushCC_popPtrGray[2] ^ _zz_io_pushOccupancy_2);
  assign _zz_io_pushOccupancy_2 = (pushCC_popPtrGray[3] ^ _zz_io_pushOccupancy_3);
  assign _zz_io_pushOccupancy_3 = (pushCC_popPtrGray[4] ^ _zz_io_pushOccupancy_4);
  assign _zz_io_pushOccupancy_4 = (pushCC_popPtrGray[5] ^ _zz_io_pushOccupancy_5);
  assign _zz_io_pushOccupancy_5 = (pushCC_popPtrGray[6] ^ _zz_io_pushOccupancy_6);
  assign _zz_io_pushOccupancy_6 = pushCC_popPtrGray[7];
  assign io_pushOccupancy = (pushCC_pushPtr - {_zz_io_pushOccupancy_6,{_zz_io_pushOccupancy_5,{_zz_io_pushOccupancy_4,{_zz_io_pushOccupancy_3,{_zz_io_pushOccupancy_2,{_zz_io_pushOccupancy_1,{_zz_io_pushOccupancy,(pushCC_popPtrGray[0] ^ _zz_io_pushOccupancy)}}}}}}});
  assign ram_axi_cc_toplevel_board_ctrl_reset_ram_asyncAssertSyncDeassert = (1'b0 ^ 1'b0);
  assign ram_axi_cc_toplevel_board_ctrl_reset_ram_synchronized = ram_axi_cc_toplevel_board_ctrl_reset_ram_asyncAssertSyncDeassert_buffercc_io_dataOut;
  assign popCC_popPtrPlus = (popCC_popPtr + 8'h01);
  assign popCC_popPtrGray = (_zz_popCC_popPtrGray ^ popCC_popPtr);
  assign popCC_pushPtrGray = pushToPopGray_buffercc_io_dataOut;
  assign popCC_empty = (popCC_popPtrGray == popCC_pushPtrGray);
  assign popCC_addressGen_valid = (! popCC_empty);
  assign popCC_addressGen_payload = popCC_popPtr[6:0];
  assign popCC_addressGen_fire = (popCC_addressGen_valid && popCC_addressGen_ready);
  always @(*) begin
    popCC_addressGen_ready = popCC_readArbitation_ready;
    if(when_Stream_l393) begin
      popCC_addressGen_ready = 1'b1;
    end
  end

  assign when_Stream_l393 = (! popCC_readArbitation_valid);
  assign popCC_readArbitation_valid = popCC_addressGen_rValid;
  assign popCC_readArbitation_payload = popCC_addressGen_rData;
  assign _zz_popCC_readPort_rsp_data = ram_1_spinal_port1;
  assign popCC_readPort_rsp_data = _zz_popCC_readPort_rsp_data[63 : 0];
  assign popCC_readPort_rsp_id = _zz_popCC_readPort_rsp_data[66 : 64];
  assign popCC_readPort_rsp_resp = _zz_popCC_readPort_rsp_data[68 : 67];
  assign popCC_readPort_rsp_last = _zz_popCC_readPort_rsp_data[69];
  assign popCC_readPort_cmd_valid = popCC_addressGen_fire;
  assign popCC_readPort_cmd_payload = popCC_addressGen_payload;
  assign popCC_readArbitation_translated_valid = popCC_readArbitation_valid;
  assign popCC_readArbitation_ready = popCC_readArbitation_translated_ready;
  assign popCC_readArbitation_translated_payload_data = popCC_readPort_rsp_data;
  assign popCC_readArbitation_translated_payload_id = popCC_readPort_rsp_id;
  assign popCC_readArbitation_translated_payload_resp = popCC_readPort_rsp_resp;
  assign popCC_readArbitation_translated_payload_last = popCC_readPort_rsp_last;
  assign io_pop_valid = popCC_readArbitation_translated_valid;
  assign popCC_readArbitation_translated_ready = io_pop_ready;
  assign io_pop_payload_data = popCC_readArbitation_translated_payload_data;
  assign io_pop_payload_id = popCC_readArbitation_translated_payload_id;
  assign io_pop_payload_resp = popCC_readArbitation_translated_payload_resp;
  assign io_pop_payload_last = popCC_readArbitation_translated_payload_last;
  assign popCC_readArbitation_fire = (popCC_readArbitation_valid && popCC_readArbitation_ready);
  assign _zz_io_popOccupancy = (popCC_pushPtrGray[1] ^ _zz_io_popOccupancy_1);
  assign _zz_io_popOccupancy_1 = (popCC_pushPtrGray[2] ^ _zz_io_popOccupancy_2);
  assign _zz_io_popOccupancy_2 = (popCC_pushPtrGray[3] ^ _zz_io_popOccupancy_3);
  assign _zz_io_popOccupancy_3 = (popCC_pushPtrGray[4] ^ _zz_io_popOccupancy_4);
  assign _zz_io_popOccupancy_4 = (popCC_pushPtrGray[5] ^ _zz_io_popOccupancy_5);
  assign _zz_io_popOccupancy_5 = (popCC_pushPtrGray[6] ^ _zz_io_popOccupancy_6);
  assign _zz_io_popOccupancy_6 = popCC_pushPtrGray[7];
  assign io_popOccupancy = ({_zz_io_popOccupancy_6,{_zz_io_popOccupancy_5,{_zz_io_popOccupancy_4,{_zz_io_popOccupancy_3,{_zz_io_popOccupancy_2,{_zz_io_popOccupancy_1,{_zz_io_popOccupancy,(popCC_pushPtrGray[0] ^ _zz_io_popOccupancy)}}}}}}} - popCC_ptrToOccupancy);
  assign pushToPopGray = pushCC_pushPtrGray;
  assign popToPushGray = popCC_ptrToPush;
  assign ram_axi_cc_toplevel_board_ctrl_reset_ram_synchronized_1 = ram_axi_cc_toplevel_board_ctrl_reset_ram_synchronized;
  always @(posedge clk_ram_bus or posedge reset_ram) begin
    if(reset_ram) begin
      pushCC_pushPtr <= 8'h0;
      pushCC_pushPtrGray <= 8'h0;
    end else begin
      if(io_push_fire) begin
        pushCC_pushPtrGray <= (_zz_pushCC_pushPtrGray ^ pushCC_pushPtrPlus);
      end
      if(io_push_fire) begin
        pushCC_pushPtr <= pushCC_pushPtrPlus;
      end
    end
  end

  always @(posedge clk_cpu or posedge ram_axi_cc_toplevel_board_ctrl_reset_ram_synchronized) begin
    if(ram_axi_cc_toplevel_board_ctrl_reset_ram_synchronized) begin
      popCC_popPtr <= 8'h0;
      popCC_addressGen_rValid <= 1'b0;
      popCC_ptrToPush <= 8'h0;
      popCC_ptrToOccupancy <= 8'h0;
    end else begin
      if(popCC_addressGen_fire) begin
        popCC_popPtr <= popCC_popPtrPlus;
      end
      if(popCC_addressGen_ready) begin
        popCC_addressGen_rValid <= popCC_addressGen_valid;
      end
      if(popCC_readArbitation_fire) begin
        popCC_ptrToPush <= popCC_popPtrGray;
      end
      if(popCC_readArbitation_fire) begin
        popCC_ptrToOccupancy <= popCC_popPtr;
      end
    end
  end

  always @(posedge clk_cpu) begin
    if(popCC_addressGen_ready) begin
      popCC_addressGen_rData <= popCC_addressGen_payload;
    end
  end


endmodule

module StreamFifoCC (
  input  wire          io_push_valid,
  output wire          io_push_ready,
  input  wire [26:0]   io_push_payload_addr,
  input  wire [2:0]    io_push_payload_id,
  input  wire [7:0]    io_push_payload_len,
  input  wire [2:0]    io_push_payload_size,
  input  wire [1:0]    io_push_payload_burst,
  input  wire          io_push_payload_allStrb,
  input  wire          io_push_payload_write,
  output wire          io_pop_valid,
  input  wire          io_pop_ready,
  output wire [26:0]   io_pop_payload_addr,
  output wire [2:0]    io_pop_payload_id,
  output wire [7:0]    io_pop_payload_len,
  output wire [2:0]    io_pop_payload_size,
  output wire [1:0]    io_pop_payload_burst,
  output wire          io_pop_payload_allStrb,
  output wire          io_pop_payload_write,
  output wire [1:0]    io_pushOccupancy,
  output wire [1:0]    io_popOccupancy,
  input  wire          clk_cpu,
  input  wire          reset_cpu,
  input  wire          clk_ram_bus,
  output wire          ram_axi_cc_toplevel_board_ctrl_reset_cpu_synchronized_1
);

  reg        [44:0]   ram_1_spinal_port1;
  wire       [1:0]    popToPushGray_buffercc_io_dataOut;
  wire                ram_axi_cc_toplevel_board_ctrl_reset_cpu_asyncAssertSyncDeassert_buffercc_io_dataOut;
  wire       [1:0]    pushToPopGray_buffercc_io_dataOut;
  wire       [1:0]    _zz_pushCC_pushPtrGray;
  wire       [0:0]    _zz_ram_1_port;
  wire       [44:0]   _zz_ram_1_port_1;
  wire       [1:0]    _zz_popCC_popPtrGray;
  reg                 _zz_1;
  wire       [1:0]    popToPushGray;
  wire       [1:0]    pushToPopGray;
  reg        [1:0]    pushCC_pushPtr;
  wire       [1:0]    pushCC_pushPtrPlus;
  wire                io_push_fire;
  reg        [1:0]    pushCC_pushPtrGray;
  wire       [1:0]    pushCC_popPtrGray;
  wire                pushCC_full;
  wire                _zz_io_pushOccupancy;
  wire                ram_axi_cc_toplevel_board_ctrl_reset_cpu_asyncAssertSyncDeassert;
  wire                ram_axi_cc_toplevel_board_ctrl_reset_cpu_synchronized;
  reg        [1:0]    popCC_popPtr;
  (* keep , syn_keep *) wire       [1:0]    popCC_popPtrPlus /* synthesis syn_keep = 1 */ ;
  wire       [1:0]    popCC_popPtrGray;
  wire       [1:0]    popCC_pushPtrGray;
  wire                popCC_addressGen_valid;
  reg                 popCC_addressGen_ready;
  wire       [0:0]    popCC_addressGen_payload;
  wire                popCC_empty;
  wire                popCC_addressGen_fire;
  wire                popCC_readArbitation_valid;
  wire                popCC_readArbitation_ready;
  wire       [0:0]    popCC_readArbitation_payload;
  reg                 popCC_addressGen_rValid;
  reg        [0:0]    popCC_addressGen_rData;
  wire                when_Stream_l393;
  wire                popCC_readPort_cmd_valid;
  wire       [0:0]    popCC_readPort_cmd_payload;
  wire       [26:0]   popCC_readPort_rsp_addr;
  wire       [2:0]    popCC_readPort_rsp_id;
  wire       [7:0]    popCC_readPort_rsp_len;
  wire       [2:0]    popCC_readPort_rsp_size;
  wire       [1:0]    popCC_readPort_rsp_burst;
  wire                popCC_readPort_rsp_allStrb;
  wire                popCC_readPort_rsp_write;
  wire       [44:0]   _zz_popCC_readPort_rsp_addr;
  wire                popCC_readArbitation_translated_valid;
  wire                popCC_readArbitation_translated_ready;
  wire       [26:0]   popCC_readArbitation_translated_payload_addr;
  wire       [2:0]    popCC_readArbitation_translated_payload_id;
  wire       [7:0]    popCC_readArbitation_translated_payload_len;
  wire       [2:0]    popCC_readArbitation_translated_payload_size;
  wire       [1:0]    popCC_readArbitation_translated_payload_burst;
  wire                popCC_readArbitation_translated_payload_allStrb;
  wire                popCC_readArbitation_translated_payload_write;
  wire                popCC_readArbitation_fire;
  reg        [1:0]    popCC_ptrToPush;
  reg        [1:0]    popCC_ptrToOccupancy;
  wire                _zz_io_popOccupancy;
  reg [44:0] ram_1 [0:1];

  assign _zz_pushCC_pushPtrGray = (pushCC_pushPtrPlus >>> 1'b1);
  assign _zz_ram_1_port = pushCC_pushPtr[0:0];
  assign _zz_popCC_popPtrGray = (popCC_popPtr >>> 1'b1);
  assign _zz_ram_1_port_1 = {io_push_payload_write,{io_push_payload_allStrb,{io_push_payload_burst,{io_push_payload_size,{io_push_payload_len,{io_push_payload_id,io_push_payload_addr}}}}}};
  always @(posedge clk_cpu) begin
    if(_zz_1) begin
      ram_1[_zz_ram_1_port] <= _zz_ram_1_port_1;
    end
  end

  always @(posedge clk_ram_bus) begin
    if(popCC_readPort_cmd_valid) begin
      ram_1_spinal_port1 <= ram_1[popCC_readPort_cmd_payload];
    end
  end

  (* keep_hierarchy = "TRUE" *) BufferCC popToPushGray_buffercc (
    .io_dataIn  (popToPushGray[1:0]                    ), //i
    .io_dataOut (popToPushGray_buffercc_io_dataOut[1:0]), //o
    .clk_cpu    (clk_cpu                               ), //i
    .reset_cpu  (reset_cpu                             )  //i
  );
  (* keep_hierarchy = "TRUE" *) BufferCC_1 ram_axi_cc_toplevel_board_ctrl_reset_cpu_asyncAssertSyncDeassert_buffercc (
    .io_dataIn   (ram_axi_cc_toplevel_board_ctrl_reset_cpu_asyncAssertSyncDeassert                    ), //i
    .io_dataOut  (ram_axi_cc_toplevel_board_ctrl_reset_cpu_asyncAssertSyncDeassert_buffercc_io_dataOut), //o
    .clk_ram_bus (clk_ram_bus                                                                         ), //i
    .reset_cpu   (reset_cpu                                                                           )  //i
  );
  (* keep_hierarchy = "TRUE" *) BufferCC_2 pushToPopGray_buffercc (
    .io_dataIn                                             (pushToPopGray[1:0]                                   ), //i
    .io_dataOut                                            (pushToPopGray_buffercc_io_dataOut[1:0]               ), //o
    .clk_ram_bus                                           (clk_ram_bus                                          ), //i
    .ram_axi_cc_toplevel_board_ctrl_reset_cpu_synchronized (ram_axi_cc_toplevel_board_ctrl_reset_cpu_synchronized)  //i
  );
  always @(*) begin
    _zz_1 = 1'b0;
    if(io_push_fire) begin
      _zz_1 = 1'b1;
    end
  end

  assign pushCC_pushPtrPlus = (pushCC_pushPtr + 2'b01);
  assign io_push_fire = (io_push_valid && io_push_ready);
  assign pushCC_popPtrGray = popToPushGray_buffercc_io_dataOut;
  assign pushCC_full = ((pushCC_pushPtrGray[1 : 0] == (~ pushCC_popPtrGray[1 : 0])) && 1'b1);
  assign io_push_ready = (! pushCC_full);
  assign _zz_io_pushOccupancy = pushCC_popPtrGray[1];
  assign io_pushOccupancy = (pushCC_pushPtr - {_zz_io_pushOccupancy,(pushCC_popPtrGray[0] ^ _zz_io_pushOccupancy)});
  assign ram_axi_cc_toplevel_board_ctrl_reset_cpu_asyncAssertSyncDeassert = (1'b0 ^ 1'b0);
  assign ram_axi_cc_toplevel_board_ctrl_reset_cpu_synchronized = ram_axi_cc_toplevel_board_ctrl_reset_cpu_asyncAssertSyncDeassert_buffercc_io_dataOut;
  assign popCC_popPtrPlus = (popCC_popPtr + 2'b01);
  assign popCC_popPtrGray = (_zz_popCC_popPtrGray ^ popCC_popPtr);
  assign popCC_pushPtrGray = pushToPopGray_buffercc_io_dataOut;
  assign popCC_empty = (popCC_popPtrGray == popCC_pushPtrGray);
  assign popCC_addressGen_valid = (! popCC_empty);
  assign popCC_addressGen_payload = popCC_popPtr[0:0];
  assign popCC_addressGen_fire = (popCC_addressGen_valid && popCC_addressGen_ready);
  always @(*) begin
    popCC_addressGen_ready = popCC_readArbitation_ready;
    if(when_Stream_l393) begin
      popCC_addressGen_ready = 1'b1;
    end
  end

  assign when_Stream_l393 = (! popCC_readArbitation_valid);
  assign popCC_readArbitation_valid = popCC_addressGen_rValid;
  assign popCC_readArbitation_payload = popCC_addressGen_rData;
  assign _zz_popCC_readPort_rsp_addr = ram_1_spinal_port1;
  assign popCC_readPort_rsp_addr = _zz_popCC_readPort_rsp_addr[26 : 0];
  assign popCC_readPort_rsp_id = _zz_popCC_readPort_rsp_addr[29 : 27];
  assign popCC_readPort_rsp_len = _zz_popCC_readPort_rsp_addr[37 : 30];
  assign popCC_readPort_rsp_size = _zz_popCC_readPort_rsp_addr[40 : 38];
  assign popCC_readPort_rsp_burst = _zz_popCC_readPort_rsp_addr[42 : 41];
  assign popCC_readPort_rsp_allStrb = _zz_popCC_readPort_rsp_addr[43];
  assign popCC_readPort_rsp_write = _zz_popCC_readPort_rsp_addr[44];
  assign popCC_readPort_cmd_valid = popCC_addressGen_fire;
  assign popCC_readPort_cmd_payload = popCC_addressGen_payload;
  assign popCC_readArbitation_translated_valid = popCC_readArbitation_valid;
  assign popCC_readArbitation_ready = popCC_readArbitation_translated_ready;
  assign popCC_readArbitation_translated_payload_addr = popCC_readPort_rsp_addr;
  assign popCC_readArbitation_translated_payload_id = popCC_readPort_rsp_id;
  assign popCC_readArbitation_translated_payload_len = popCC_readPort_rsp_len;
  assign popCC_readArbitation_translated_payload_size = popCC_readPort_rsp_size;
  assign popCC_readArbitation_translated_payload_burst = popCC_readPort_rsp_burst;
  assign popCC_readArbitation_translated_payload_allStrb = popCC_readPort_rsp_allStrb;
  assign popCC_readArbitation_translated_payload_write = popCC_readPort_rsp_write;
  assign io_pop_valid = popCC_readArbitation_translated_valid;
  assign popCC_readArbitation_translated_ready = io_pop_ready;
  assign io_pop_payload_addr = popCC_readArbitation_translated_payload_addr;
  assign io_pop_payload_id = popCC_readArbitation_translated_payload_id;
  assign io_pop_payload_len = popCC_readArbitation_translated_payload_len;
  assign io_pop_payload_size = popCC_readArbitation_translated_payload_size;
  assign io_pop_payload_burst = popCC_readArbitation_translated_payload_burst;
  assign io_pop_payload_allStrb = popCC_readArbitation_translated_payload_allStrb;
  assign io_pop_payload_write = popCC_readArbitation_translated_payload_write;
  assign popCC_readArbitation_fire = (popCC_readArbitation_valid && popCC_readArbitation_ready);
  assign _zz_io_popOccupancy = popCC_pushPtrGray[1];
  assign io_popOccupancy = ({_zz_io_popOccupancy,(popCC_pushPtrGray[0] ^ _zz_io_popOccupancy)} - popCC_ptrToOccupancy);
  assign pushToPopGray = pushCC_pushPtrGray;
  assign popToPushGray = popCC_ptrToPush;
  assign ram_axi_cc_toplevel_board_ctrl_reset_cpu_synchronized_1 = ram_axi_cc_toplevel_board_ctrl_reset_cpu_synchronized;
  always @(posedge clk_cpu or posedge reset_cpu) begin
    if(reset_cpu) begin
      pushCC_pushPtr <= 2'b00;
      pushCC_pushPtrGray <= 2'b00;
    end else begin
      if(io_push_fire) begin
        pushCC_pushPtrGray <= (_zz_pushCC_pushPtrGray ^ pushCC_pushPtrPlus);
      end
      if(io_push_fire) begin
        pushCC_pushPtr <= pushCC_pushPtrPlus;
      end
    end
  end

  always @(posedge clk_ram_bus or posedge ram_axi_cc_toplevel_board_ctrl_reset_cpu_synchronized) begin
    if(ram_axi_cc_toplevel_board_ctrl_reset_cpu_synchronized) begin
      popCC_popPtr <= 2'b00;
      popCC_addressGen_rValid <= 1'b0;
      popCC_ptrToPush <= 2'b00;
      popCC_ptrToOccupancy <= 2'b00;
    end else begin
      if(popCC_addressGen_fire) begin
        popCC_popPtr <= popCC_popPtrPlus;
      end
      if(popCC_addressGen_ready) begin
        popCC_addressGen_rValid <= popCC_addressGen_valid;
      end
      if(popCC_readArbitation_fire) begin
        popCC_ptrToPush <= popCC_popPtrGray;
      end
      if(popCC_readArbitation_fire) begin
        popCC_ptrToOccupancy <= popCC_popPtr;
      end
    end
  end

  always @(posedge clk_ram_bus) begin
    if(popCC_addressGen_ready) begin
      popCC_addressGen_rData <= popCC_addressGen_payload;
    end
  end


endmodule

module ContextAsyncBufferFull_1 (
  input  wire          io_add_valid,
  output wire          io_add_ready,
  input  wire [0:0]    io_add_payload_context,
  input  wire          io_remove_valid,
  output wire [0:0]    io_query_context,
  input  wire          clk_cpu,
  input  wire          reset_cpu
);

  reg                 when_Phase_l773;
  wire                write_valid;
  wire       [0:0]    write_payload_data;
  wire       [0:0]    read_data;
  wire       [0:0]    _zz_read_data;
  reg        [0:0]    _zz_read_data_1;

  always @(*) begin
    when_Phase_l773 = 1'b0;
    if(write_valid) begin
      when_Phase_l773 = 1'b1;
    end
  end

  assign write_valid = io_add_valid;
  assign write_payload_data = io_add_payload_context;
  assign io_add_ready = 1'b1;
  assign read_data = _zz_read_data;
  assign io_query_context = read_data;
  assign _zz_read_data = _zz_read_data_1;
  always @(posedge clk_cpu) begin
    if(when_Phase_l773) begin
      _zz_read_data_1 <= write_payload_data;
    end
  end


endmodule

module StreamArbiter_6 (
  input  wire          io_inputs_0_valid,
  output wire          io_inputs_0_ready,
  input  wire [2:0]    io_inputs_0_payload_source,
  input  wire          io_inputs_0_payload_denied,
  input  wire          io_inputs_0_payload_last,
  input  wire          io_inputs_1_valid,
  output wire          io_inputs_1_ready,
  input  wire [2:0]    io_inputs_1_payload_source,
  input  wire          io_inputs_1_payload_denied,
  input  wire          io_inputs_1_payload_last,
  output wire          io_output_valid,
  input  wire          io_output_ready,
  output wire [2:0]    io_output_payload_source,
  output wire          io_output_payload_denied,
  output wire          io_output_payload_last,
  output wire [0:0]    io_chosen,
  output wire [1:0]    io_chosenOH,
  input  wire          clk_cpu,
  input  wire          reset_cpu
);

  wire       [3:0]    _zz__zz_maskProposal_0_2;
  wire       [3:0]    _zz__zz_maskProposal_0_2_1;
  wire       [1:0]    _zz__zz_maskProposal_0_2_2;
  reg                 locked;
  wire                maskProposal_0;
  wire                maskProposal_1;
  reg                 maskLocked_0;
  reg                 maskLocked_1;
  wire                maskRouted_0;
  wire                maskRouted_1;
  wire       [1:0]    _zz_maskProposal_0;
  wire       [3:0]    _zz_maskProposal_0_1;
  wire       [3:0]    _zz_maskProposal_0_2;
  wire       [1:0]    _zz_maskProposal_0_3;
  wire                io_output_fire;
  wire                when_Stream_l794;
  wire                _zz_io_chosen;

  assign _zz__zz_maskProposal_0_2 = (_zz_maskProposal_0_1 - _zz__zz_maskProposal_0_2_1);
  assign _zz__zz_maskProposal_0_2_2 = {maskLocked_0,maskLocked_1};
  assign _zz__zz_maskProposal_0_2_1 = {2'd0, _zz__zz_maskProposal_0_2_2};
  assign maskRouted_0 = (locked ? maskLocked_0 : maskProposal_0);
  assign maskRouted_1 = (locked ? maskLocked_1 : maskProposal_1);
  assign _zz_maskProposal_0 = {io_inputs_1_valid,io_inputs_0_valid};
  assign _zz_maskProposal_0_1 = {_zz_maskProposal_0,_zz_maskProposal_0};
  assign _zz_maskProposal_0_2 = (_zz_maskProposal_0_1 & (~ _zz__zz_maskProposal_0_2));
  assign _zz_maskProposal_0_3 = (_zz_maskProposal_0_2[3 : 2] | _zz_maskProposal_0_2[1 : 0]);
  assign maskProposal_0 = _zz_maskProposal_0_3[0];
  assign maskProposal_1 = _zz_maskProposal_0_3[1];
  assign io_output_fire = (io_output_valid && io_output_ready);
  assign when_Stream_l794 = (io_output_fire && io_output_payload_last);
  assign io_output_valid = ((io_inputs_0_valid && maskRouted_0) || (io_inputs_1_valid && maskRouted_1));
  assign io_output_payload_source = (maskRouted_0 ? io_inputs_0_payload_source : io_inputs_1_payload_source);
  assign io_output_payload_denied = (maskRouted_0 ? io_inputs_0_payload_denied : io_inputs_1_payload_denied);
  assign io_output_payload_last = (maskRouted_0 ? io_inputs_0_payload_last : io_inputs_1_payload_last);
  assign io_inputs_0_ready = (maskRouted_0 && io_output_ready);
  assign io_inputs_1_ready = (maskRouted_1 && io_output_ready);
  assign io_chosenOH = {maskRouted_1,maskRouted_0};
  assign _zz_io_chosen = io_chosenOH[1];
  assign io_chosen = _zz_io_chosen;
  always @(posedge clk_cpu or posedge reset_cpu) begin
    if(reset_cpu) begin
      locked <= 1'b0;
      maskLocked_0 <= 1'b0;
      maskLocked_1 <= 1'b1;
    end else begin
      if(io_output_valid) begin
        maskLocked_0 <= maskRouted_0;
        maskLocked_1 <= maskRouted_1;
      end
      if(io_output_valid) begin
        locked <= 1'b1;
      end
      if(when_Stream_l794) begin
        locked <= 1'b0;
      end
    end
  end


endmodule

module ContextAsyncBufferFull (
  input  wire          io_add_valid,
  output wire          io_add_ready,
  input  wire [2:0]    io_add_payload_id,
  input  wire [2:0]    io_add_payload_context,
  input  wire          io_remove_valid,
  input  wire [2:0]    io_remove_payload_id,
  input  wire [2:0]    io_query_id,
  output wire [2:0]    io_query_context,
  input  wire          clk_cpu,
  input  wire          reset_cpu
);

  wire       [2:0]    contexts_spinal_port1;
  wire       [2:0]    _zz_contexts_port;
  reg                 _zz_1;
  wire                write_valid;
  wire       [2:0]    write_payload_address;
  wire       [2:0]    write_payload_data;
  wire       [2:0]    read_address;
  wire       [2:0]    read_data;
  (* ram_style = "distributed" *) reg [2:0] contexts [0:7];

  assign _zz_contexts_port = write_payload_data;
  always @(posedge clk_cpu) begin
    if(_zz_1) begin
      contexts[write_payload_address] <= _zz_contexts_port;
    end
  end

  assign contexts_spinal_port1 = contexts[read_address];
  always @(*) begin
    _zz_1 = 1'b0;
    if(write_valid) begin
      _zz_1 = 1'b1;
    end
  end

  assign write_valid = io_add_valid;
  assign write_payload_address = io_add_payload_id;
  assign write_payload_data = io_add_payload_context;
  assign io_add_ready = 1'b1;
  assign read_data = contexts_spinal_port1;
  assign read_address = io_query_id;
  assign io_query_context = read_data;

endmodule

module StreamArbiter_5 (
  input  wire          io_inputs_0_valid,
  output wire          io_inputs_0_ready,
  input  wire [2:0]    io_inputs_0_payload_opcode,
  input  wire [2:0]    io_inputs_0_payload_param,
  input  wire [2:0]    io_inputs_0_payload_source,
  input  wire [31:0]   io_inputs_0_payload_address,
  input  wire [2:0]    io_inputs_0_payload_size,
  input  wire [7:0]    io_inputs_0_payload_mask,
  input  wire [63:0]   io_inputs_0_payload_data,
  input  wire          io_inputs_0_payload_corrupt,
  input  wire          io_inputs_1_valid,
  output wire          io_inputs_1_ready,
  input  wire [2:0]    io_inputs_1_payload_opcode,
  input  wire [2:0]    io_inputs_1_payload_param,
  input  wire [2:0]    io_inputs_1_payload_source,
  input  wire [31:0]   io_inputs_1_payload_address,
  input  wire [2:0]    io_inputs_1_payload_size,
  input  wire [7:0]    io_inputs_1_payload_mask,
  input  wire [63:0]   io_inputs_1_payload_data,
  input  wire          io_inputs_1_payload_corrupt,
  input  wire          io_inputs_2_valid,
  output wire          io_inputs_2_ready,
  input  wire [2:0]    io_inputs_2_payload_opcode,
  input  wire [2:0]    io_inputs_2_payload_param,
  input  wire [2:0]    io_inputs_2_payload_source,
  input  wire [31:0]   io_inputs_2_payload_address,
  input  wire [2:0]    io_inputs_2_payload_size,
  input  wire [7:0]    io_inputs_2_payload_mask,
  input  wire [63:0]   io_inputs_2_payload_data,
  input  wire          io_inputs_2_payload_corrupt,
  output wire          io_output_valid,
  input  wire          io_output_ready,
  output wire [2:0]    io_output_payload_opcode,
  output wire [2:0]    io_output_payload_param,
  output wire [2:0]    io_output_payload_source,
  output wire [31:0]   io_output_payload_address,
  output wire [2:0]    io_output_payload_size,
  output wire [7:0]    io_output_payload_mask,
  output wire [63:0]   io_output_payload_data,
  output wire          io_output_payload_corrupt,
  output wire [1:0]    io_chosen,
  output wire [2:0]    io_chosenOH,
  input  wire          clk_cpu,
  input  wire          reset_cpu
);
  localparam A_PUT_FULL_DATA = 3'd0;
  localparam A_PUT_PARTIAL_DATA = 3'd1;
  localparam A_GET = 3'd4;
  localparam A_ACQUIRE_BLOCK = 3'd6;
  localparam A_ACQUIRE_PERM = 3'd7;

  wire       [5:0]    _zz__zz_maskProposal_0_2;
  wire       [5:0]    _zz__zz_maskProposal_0_2_1;
  wire       [2:0]    _zz__zz_maskProposal_0_2_2;
  reg        [2:0]    _zz_io_output_tracker_last;
  reg        [2:0]    _zz__zz_io_output_payload_opcode;
  reg        [2:0]    _zz_io_output_payload_param_1;
  reg        [2:0]    _zz_io_output_payload_source;
  reg        [31:0]   _zz_io_output_payload_address;
  reg        [2:0]    _zz_io_output_payload_size;
  reg        [7:0]    _zz_io_output_payload_mask;
  reg        [63:0]   _zz_io_output_payload_data;
  reg                 _zz_io_output_payload_corrupt;
  reg                 locked;
  wire                maskProposal_0;
  wire                maskProposal_1;
  wire                maskProposal_2;
  reg                 maskLocked_0;
  reg                 maskLocked_1;
  reg                 maskLocked_2;
  wire                maskRouted_0;
  wire                maskRouted_1;
  wire                maskRouted_2;
  wire       [2:0]    _zz_maskProposal_0;
  wire       [5:0]    _zz_maskProposal_0_1;
  wire       [5:0]    _zz_maskProposal_0_2;
  wire       [2:0]    _zz_maskProposal_0_3;
  wire                io_output_fire;
  reg        [2:0]    io_output_tracker_beat;
  wire                io_output_tracker_last;
  wire                when_Stream_l794;
  wire       [1:0]    _zz_io_output_payload_param;
  wire       [2:0]    _zz_io_output_payload_opcode;
  wire                _zz_io_chosen;
  wire                _zz_io_chosen_1;
  `ifndef SYNTHESIS
  reg [127:0] io_inputs_0_payload_opcode_string;
  reg [127:0] io_inputs_1_payload_opcode_string;
  reg [127:0] io_inputs_2_payload_opcode_string;
  reg [127:0] io_output_payload_opcode_string;
  reg [127:0] _zz_io_output_payload_opcode_string;
  `endif


  assign _zz__zz_maskProposal_0_2 = (_zz_maskProposal_0_1 - _zz__zz_maskProposal_0_2_1);
  assign _zz__zz_maskProposal_0_2_2 = {maskLocked_1,{maskLocked_0,maskLocked_2}};
  assign _zz__zz_maskProposal_0_2_1 = {3'd0, _zz__zz_maskProposal_0_2_2};
  always @(*) begin
    case(io_output_payload_size)
      3'b000 : _zz_io_output_tracker_last = 3'b000;
      3'b001 : _zz_io_output_tracker_last = 3'b000;
      3'b010 : _zz_io_output_tracker_last = 3'b000;
      3'b011 : _zz_io_output_tracker_last = 3'b000;
      3'b100 : _zz_io_output_tracker_last = 3'b001;
      3'b101 : _zz_io_output_tracker_last = 3'b011;
      default : _zz_io_output_tracker_last = 3'b111;
    endcase
  end

  always @(*) begin
    case(_zz_io_output_payload_param)
      2'b00 : begin
        _zz__zz_io_output_payload_opcode = io_inputs_0_payload_opcode;
        _zz_io_output_payload_param_1 = io_inputs_0_payload_param;
        _zz_io_output_payload_source = io_inputs_0_payload_source;
        _zz_io_output_payload_address = io_inputs_0_payload_address;
        _zz_io_output_payload_size = io_inputs_0_payload_size;
        _zz_io_output_payload_mask = io_inputs_0_payload_mask;
        _zz_io_output_payload_data = io_inputs_0_payload_data;
        _zz_io_output_payload_corrupt = io_inputs_0_payload_corrupt;
      end
      2'b01 : begin
        _zz__zz_io_output_payload_opcode = io_inputs_1_payload_opcode;
        _zz_io_output_payload_param_1 = io_inputs_1_payload_param;
        _zz_io_output_payload_source = io_inputs_1_payload_source;
        _zz_io_output_payload_address = io_inputs_1_payload_address;
        _zz_io_output_payload_size = io_inputs_1_payload_size;
        _zz_io_output_payload_mask = io_inputs_1_payload_mask;
        _zz_io_output_payload_data = io_inputs_1_payload_data;
        _zz_io_output_payload_corrupt = io_inputs_1_payload_corrupt;
      end
      default : begin
        _zz__zz_io_output_payload_opcode = io_inputs_2_payload_opcode;
        _zz_io_output_payload_param_1 = io_inputs_2_payload_param;
        _zz_io_output_payload_source = io_inputs_2_payload_source;
        _zz_io_output_payload_address = io_inputs_2_payload_address;
        _zz_io_output_payload_size = io_inputs_2_payload_size;
        _zz_io_output_payload_mask = io_inputs_2_payload_mask;
        _zz_io_output_payload_data = io_inputs_2_payload_data;
        _zz_io_output_payload_corrupt = io_inputs_2_payload_corrupt;
      end
    endcase
  end

  `ifndef SYNTHESIS
  always @(*) begin
    case(io_inputs_0_payload_opcode)
      A_PUT_FULL_DATA : io_inputs_0_payload_opcode_string = "PUT_FULL_DATA   ";
      A_PUT_PARTIAL_DATA : io_inputs_0_payload_opcode_string = "PUT_PARTIAL_DATA";
      A_GET : io_inputs_0_payload_opcode_string = "GET             ";
      A_ACQUIRE_BLOCK : io_inputs_0_payload_opcode_string = "ACQUIRE_BLOCK   ";
      A_ACQUIRE_PERM : io_inputs_0_payload_opcode_string = "ACQUIRE_PERM    ";
      default : io_inputs_0_payload_opcode_string = "????????????????";
    endcase
  end
  always @(*) begin
    case(io_inputs_1_payload_opcode)
      A_PUT_FULL_DATA : io_inputs_1_payload_opcode_string = "PUT_FULL_DATA   ";
      A_PUT_PARTIAL_DATA : io_inputs_1_payload_opcode_string = "PUT_PARTIAL_DATA";
      A_GET : io_inputs_1_payload_opcode_string = "GET             ";
      A_ACQUIRE_BLOCK : io_inputs_1_payload_opcode_string = "ACQUIRE_BLOCK   ";
      A_ACQUIRE_PERM : io_inputs_1_payload_opcode_string = "ACQUIRE_PERM    ";
      default : io_inputs_1_payload_opcode_string = "????????????????";
    endcase
  end
  always @(*) begin
    case(io_inputs_2_payload_opcode)
      A_PUT_FULL_DATA : io_inputs_2_payload_opcode_string = "PUT_FULL_DATA   ";
      A_PUT_PARTIAL_DATA : io_inputs_2_payload_opcode_string = "PUT_PARTIAL_DATA";
      A_GET : io_inputs_2_payload_opcode_string = "GET             ";
      A_ACQUIRE_BLOCK : io_inputs_2_payload_opcode_string = "ACQUIRE_BLOCK   ";
      A_ACQUIRE_PERM : io_inputs_2_payload_opcode_string = "ACQUIRE_PERM    ";
      default : io_inputs_2_payload_opcode_string = "????????????????";
    endcase
  end
  always @(*) begin
    case(io_output_payload_opcode)
      A_PUT_FULL_DATA : io_output_payload_opcode_string = "PUT_FULL_DATA   ";
      A_PUT_PARTIAL_DATA : io_output_payload_opcode_string = "PUT_PARTIAL_DATA";
      A_GET : io_output_payload_opcode_string = "GET             ";
      A_ACQUIRE_BLOCK : io_output_payload_opcode_string = "ACQUIRE_BLOCK   ";
      A_ACQUIRE_PERM : io_output_payload_opcode_string = "ACQUIRE_PERM    ";
      default : io_output_payload_opcode_string = "????????????????";
    endcase
  end
  always @(*) begin
    case(_zz_io_output_payload_opcode)
      A_PUT_FULL_DATA : _zz_io_output_payload_opcode_string = "PUT_FULL_DATA   ";
      A_PUT_PARTIAL_DATA : _zz_io_output_payload_opcode_string = "PUT_PARTIAL_DATA";
      A_GET : _zz_io_output_payload_opcode_string = "GET             ";
      A_ACQUIRE_BLOCK : _zz_io_output_payload_opcode_string = "ACQUIRE_BLOCK   ";
      A_ACQUIRE_PERM : _zz_io_output_payload_opcode_string = "ACQUIRE_PERM    ";
      default : _zz_io_output_payload_opcode_string = "????????????????";
    endcase
  end
  `endif

  assign maskRouted_0 = (locked ? maskLocked_0 : maskProposal_0);
  assign maskRouted_1 = (locked ? maskLocked_1 : maskProposal_1);
  assign maskRouted_2 = (locked ? maskLocked_2 : maskProposal_2);
  assign _zz_maskProposal_0 = {io_inputs_2_valid,{io_inputs_1_valid,io_inputs_0_valid}};
  assign _zz_maskProposal_0_1 = {_zz_maskProposal_0,_zz_maskProposal_0};
  assign _zz_maskProposal_0_2 = (_zz_maskProposal_0_1 & (~ _zz__zz_maskProposal_0_2));
  assign _zz_maskProposal_0_3 = (_zz_maskProposal_0_2[5 : 3] | _zz_maskProposal_0_2[2 : 0]);
  assign maskProposal_0 = _zz_maskProposal_0_3[0];
  assign maskProposal_1 = _zz_maskProposal_0_3[1];
  assign maskProposal_2 = _zz_maskProposal_0_3[2];
  assign io_output_fire = (io_output_valid && io_output_ready);
  assign io_output_tracker_last = ((! ((1'b0 || (A_PUT_FULL_DATA == io_output_payload_opcode)) || (A_PUT_PARTIAL_DATA == io_output_payload_opcode))) || (io_output_tracker_beat == _zz_io_output_tracker_last));
  assign when_Stream_l794 = (io_output_fire && io_output_tracker_last);
  assign io_output_valid = (((io_inputs_0_valid && maskRouted_0) || (io_inputs_1_valid && maskRouted_1)) || (io_inputs_2_valid && maskRouted_2));
  assign _zz_io_output_payload_param = {maskRouted_2,maskRouted_1};
  assign _zz_io_output_payload_opcode = _zz__zz_io_output_payload_opcode;
  assign io_output_payload_opcode = _zz_io_output_payload_opcode;
  assign io_output_payload_param = _zz_io_output_payload_param_1;
  assign io_output_payload_source = _zz_io_output_payload_source;
  assign io_output_payload_address = _zz_io_output_payload_address;
  assign io_output_payload_size = _zz_io_output_payload_size;
  assign io_output_payload_mask = _zz_io_output_payload_mask;
  assign io_output_payload_data = _zz_io_output_payload_data;
  assign io_output_payload_corrupt = _zz_io_output_payload_corrupt;
  assign io_inputs_0_ready = (maskRouted_0 && io_output_ready);
  assign io_inputs_1_ready = (maskRouted_1 && io_output_ready);
  assign io_inputs_2_ready = (maskRouted_2 && io_output_ready);
  assign io_chosenOH = {maskRouted_2,{maskRouted_1,maskRouted_0}};
  assign _zz_io_chosen = io_chosenOH[1];
  assign _zz_io_chosen_1 = io_chosenOH[2];
  assign io_chosen = {_zz_io_chosen_1,_zz_io_chosen};
  always @(posedge clk_cpu or posedge reset_cpu) begin
    if(reset_cpu) begin
      locked <= 1'b0;
      maskLocked_0 <= 1'b0;
      maskLocked_1 <= 1'b0;
      maskLocked_2 <= 1'b1;
      io_output_tracker_beat <= 3'b000;
    end else begin
      if(io_output_valid) begin
        maskLocked_0 <= maskRouted_0;
        maskLocked_1 <= maskRouted_1;
        maskLocked_2 <= maskRouted_2;
      end
      if(io_output_valid) begin
        locked <= 1'b1;
      end
      if(io_output_fire) begin
        io_output_tracker_beat <= (io_output_tracker_beat + 3'b001);
        if(io_output_tracker_last) begin
          io_output_tracker_beat <= 3'b000;
        end
      end
      if(when_Stream_l794) begin
        locked <= 1'b0;
      end
    end
  end


endmodule

module RegFileMem (
  input  wire          io_writes_0_valid,
  input  wire [4:0]    io_writes_0_address,
  input  wire [31:0]   io_writes_0_data,
  input  wire [15:0]   io_writes_0_uopId,
  input  wire          io_writes_1_valid,
  input  wire [4:0]    io_writes_1_address,
  input  wire [31:0]   io_writes_1_data,
  input  wire [15:0]   io_writes_1_uopId,
  input  wire          io_reads_0_valid,
  input  wire [4:0]    io_reads_0_address,
  output wire [31:0]   io_reads_0_data,
  input  wire          io_reads_1_valid,
  input  wire [4:0]    io_reads_1_address,
  output wire [31:0]   io_reads_1_data,
  input  wire          io_reads_2_valid,
  input  wire [4:0]    io_reads_2_address,
  output wire [31:0]   io_reads_2_data,
  input  wire          io_reads_3_valid,
  input  wire [4:0]    io_reads_3_address,
  output wire [31:0]   io_reads_3_data,
  input  wire          clk_cpu,
  input  wire          reset_cpu
);

  wire       [31:0]   ramSyncMwMux_1_io_read_0_rsp;
  wire       [31:0]   ramSyncMwMux_1_io_read_1_rsp;
  wire       [31:0]   ramSyncMwMux_1_io_read_2_rsp;
  wire       [31:0]   ramSyncMwMux_1_io_read_3_rsp;
  wire                conv_writes_0_valid;
  wire       [4:0]    conv_writes_0_payload_address;
  wire       [31:0]   conv_writes_0_payload_data;
  wire                conv_writes_1_valid;
  wire       [4:0]    conv_writes_1_payload_address;
  wire       [31:0]   conv_writes_1_payload_data;
  wire                conv_read_0_cmd_valid;
  wire       [4:0]    conv_read_0_cmd_payload;
  wire       [31:0]   conv_read_0_rsp;
  wire                conv_read_1_cmd_valid;
  wire       [4:0]    conv_read_1_cmd_payload;
  wire       [31:0]   conv_read_1_rsp;
  wire                conv_read_2_cmd_valid;
  wire       [4:0]    conv_read_2_cmd_payload;
  wire       [31:0]   conv_read_2_rsp;
  wire                conv_read_3_cmd_valid;
  wire       [4:0]    conv_read_3_cmd_payload;
  wire       [31:0]   conv_read_3_rsp;

  RamSyncMwMux ramSyncMwMux_1 (
    .io_writes_0_valid           (conv_writes_0_valid               ), //i
    .io_writes_0_payload_address (conv_writes_0_payload_address[4:0]), //i
    .io_writes_0_payload_data    (conv_writes_0_payload_data[31:0]  ), //i
    .io_writes_1_valid           (conv_writes_1_valid               ), //i
    .io_writes_1_payload_address (conv_writes_1_payload_address[4:0]), //i
    .io_writes_1_payload_data    (conv_writes_1_payload_data[31:0]  ), //i
    .io_read_0_cmd_valid         (conv_read_0_cmd_valid             ), //i
    .io_read_0_cmd_payload       (conv_read_0_cmd_payload[4:0]      ), //i
    .io_read_0_rsp               (ramSyncMwMux_1_io_read_0_rsp[31:0]), //o
    .io_read_1_cmd_valid         (conv_read_1_cmd_valid             ), //i
    .io_read_1_cmd_payload       (conv_read_1_cmd_payload[4:0]      ), //i
    .io_read_1_rsp               (ramSyncMwMux_1_io_read_1_rsp[31:0]), //o
    .io_read_2_cmd_valid         (conv_read_2_cmd_valid             ), //i
    .io_read_2_cmd_payload       (conv_read_2_cmd_payload[4:0]      ), //i
    .io_read_2_rsp               (ramSyncMwMux_1_io_read_2_rsp[31:0]), //o
    .io_read_3_cmd_valid         (conv_read_3_cmd_valid             ), //i
    .io_read_3_cmd_payload       (conv_read_3_cmd_payload[4:0]      ), //i
    .io_read_3_rsp               (ramSyncMwMux_1_io_read_3_rsp[31:0]), //o
    .clk_cpu                     (clk_cpu                           ), //i
    .reset_cpu                   (reset_cpu                         )  //i
  );
  assign conv_writes_0_valid = io_writes_0_valid;
  assign conv_writes_0_payload_address = io_writes_0_address;
  assign conv_writes_0_payload_data = io_writes_0_data;
  assign conv_writes_1_valid = io_writes_1_valid;
  assign conv_writes_1_payload_address = io_writes_1_address;
  assign conv_writes_1_payload_data = io_writes_1_data;
  assign conv_read_0_cmd_valid = io_reads_0_valid;
  assign conv_read_0_cmd_payload = io_reads_0_address;
  assign io_reads_0_data = conv_read_0_rsp;
  assign conv_read_1_cmd_valid = io_reads_1_valid;
  assign conv_read_1_cmd_payload = io_reads_1_address;
  assign io_reads_1_data = conv_read_1_rsp;
  assign conv_read_2_cmd_valid = io_reads_2_valid;
  assign conv_read_2_cmd_payload = io_reads_2_address;
  assign io_reads_2_data = conv_read_2_rsp;
  assign conv_read_3_cmd_valid = io_reads_3_valid;
  assign conv_read_3_cmd_payload = io_reads_3_address;
  assign io_reads_3_data = conv_read_3_rsp;
  assign conv_read_0_rsp = ramSyncMwMux_1_io_read_0_rsp;
  assign conv_read_1_rsp = ramSyncMwMux_1_io_read_1_rsp;
  assign conv_read_2_rsp = ramSyncMwMux_1_io_read_2_rsp;
  assign conv_read_3_rsp = ramSyncMwMux_1_io_read_3_rsp;

endmodule

module StreamArbiter_4 (
  input  wire          io_inputs_0_valid,
  output wire          io_inputs_0_ready,
  output wire          io_output_valid,
  input  wire          io_output_ready,
  output wire [0:0]    io_chosenOH,
  input  wire          clk_cpu,
  input  wire          reset_cpu
);

  wire       [1:0]    _zz__zz_maskProposal_0_2;
  wire       [1:0]    _zz__zz_maskProposal_0_2_1;
  wire       [0:0]    _zz__zz_maskProposal_0_2_2;
  wire       [0:0]    _zz_maskProposal_0_3;
  reg                 locked;
  wire                maskProposal_0;
  reg                 maskLocked_0;
  wire                maskRouted_0;
  wire       [0:0]    _zz_maskProposal_0;
  wire       [1:0]    _zz_maskProposal_0_1;
  wire       [1:0]    _zz_maskProposal_0_2;
  wire                io_output_fire;

  assign _zz__zz_maskProposal_0_2 = (_zz_maskProposal_0_1 - _zz__zz_maskProposal_0_2_1);
  assign _zz__zz_maskProposal_0_2_2 = maskLocked_0;
  assign _zz__zz_maskProposal_0_2_1 = {1'd0, _zz__zz_maskProposal_0_2_2};
  assign _zz_maskProposal_0_3 = (_zz_maskProposal_0_2[1 : 1] | _zz_maskProposal_0_2[0 : 0]);
  assign maskRouted_0 = (locked ? maskLocked_0 : maskProposal_0);
  assign _zz_maskProposal_0 = io_inputs_0_valid;
  assign _zz_maskProposal_0_1 = {_zz_maskProposal_0,_zz_maskProposal_0};
  assign _zz_maskProposal_0_2 = (_zz_maskProposal_0_1 & (~ _zz__zz_maskProposal_0_2));
  assign maskProposal_0 = _zz_maskProposal_0_3[0];
  assign io_output_fire = (io_output_valid && io_output_ready);
  assign io_output_valid = (io_inputs_0_valid && maskRouted_0);
  assign io_inputs_0_ready = (maskRouted_0 && io_output_ready);
  assign io_chosenOH = maskRouted_0;
  always @(posedge clk_cpu or posedge reset_cpu) begin
    if(reset_cpu) begin
      locked <= 1'b0;
      maskLocked_0 <= 1'b1;
    end else begin
      if(io_output_valid) begin
        maskLocked_0 <= maskRouted_0;
      end
      if(io_output_valid) begin
        locked <= 1'b1;
      end
      if(io_output_fire) begin
        locked <= 1'b0;
      end
    end
  end


endmodule

module StreamArbiter_3 (
  input  wire          io_inputs_0_valid,
  output wire          io_inputs_0_ready,
  input  wire [31:0]   io_inputs_0_payload_address,
  input  wire [0:0]    io_inputs_0_payload_storageId,
  output wire          io_output_valid,
  input  wire          io_output_ready,
  output wire [31:0]   io_output_payload_address,
  output wire [0:0]    io_output_payload_storageId,
  output wire [0:0]    io_chosenOH,
  input  wire          clk_cpu,
  input  wire          reset_cpu
);

  wire       [1:0]    _zz__zz_maskProposal_0_2;
  wire       [1:0]    _zz__zz_maskProposal_0_2_1;
  wire       [0:0]    _zz__zz_maskProposal_0_2_2;
  wire       [0:0]    _zz_maskProposal_0_3;
  reg                 locked;
  wire                maskProposal_0;
  reg                 maskLocked_0;
  wire                maskRouted_0;
  wire       [0:0]    _zz_maskProposal_0;
  wire       [1:0]    _zz_maskProposal_0_1;
  wire       [1:0]    _zz_maskProposal_0_2;
  wire                io_output_fire;

  assign _zz__zz_maskProposal_0_2 = (_zz_maskProposal_0_1 - _zz__zz_maskProposal_0_2_1);
  assign _zz__zz_maskProposal_0_2_2 = maskLocked_0;
  assign _zz__zz_maskProposal_0_2_1 = {1'd0, _zz__zz_maskProposal_0_2_2};
  assign _zz_maskProposal_0_3 = (_zz_maskProposal_0_2[1 : 1] | _zz_maskProposal_0_2[0 : 0]);
  assign maskRouted_0 = (locked ? maskLocked_0 : maskProposal_0);
  assign _zz_maskProposal_0 = io_inputs_0_valid;
  assign _zz_maskProposal_0_1 = {_zz_maskProposal_0,_zz_maskProposal_0};
  assign _zz_maskProposal_0_2 = (_zz_maskProposal_0_1 & (~ _zz__zz_maskProposal_0_2));
  assign maskProposal_0 = _zz_maskProposal_0_3[0];
  assign io_output_fire = (io_output_valid && io_output_ready);
  assign io_output_valid = (io_inputs_0_valid && maskRouted_0);
  assign io_output_payload_address = io_inputs_0_payload_address;
  assign io_output_payload_storageId = io_inputs_0_payload_storageId;
  assign io_inputs_0_ready = (maskRouted_0 && io_output_ready);
  assign io_chosenOH = maskRouted_0;
  always @(posedge clk_cpu or posedge reset_cpu) begin
    if(reset_cpu) begin
      locked <= 1'b0;
      maskLocked_0 <= 1'b1;
    end else begin
      if(io_output_valid) begin
        maskLocked_0 <= maskRouted_0;
      end
      if(io_output_valid) begin
        locked <= 1'b1;
      end
      if(io_output_fire) begin
        locked <= 1'b0;
      end
    end
  end


endmodule

module StreamArbiter_2 (
  input  wire          io_inputs_0_valid,
  output wire          io_inputs_0_ready,
  input  wire [2:0]    io_inputs_0_payload_op,
  input  wire [31:0]   io_inputs_0_payload_address,
  input  wire [1:0]    io_inputs_0_payload_size,
  input  wire          io_inputs_0_payload_load,
  input  wire          io_inputs_0_payload_store,
  input  wire          io_inputs_0_payload_atomic,
  input  wire [11:0]   io_inputs_0_payload_storeId,
  input  wire          io_inputs_1_valid,
  output wire          io_inputs_1_ready,
  input  wire [2:0]    io_inputs_1_payload_op,
  input  wire [31:0]   io_inputs_1_payload_address,
  input  wire [1:0]    io_inputs_1_payload_size,
  input  wire          io_inputs_1_payload_load,
  input  wire          io_inputs_1_payload_store,
  input  wire          io_inputs_1_payload_atomic,
  input  wire [11:0]   io_inputs_1_payload_storeId,
  input  wire          io_inputs_2_valid,
  output wire          io_inputs_2_ready,
  input  wire [2:0]    io_inputs_2_payload_op,
  input  wire [31:0]   io_inputs_2_payload_address,
  input  wire [1:0]    io_inputs_2_payload_size,
  input  wire          io_inputs_2_payload_load,
  input  wire          io_inputs_2_payload_store,
  input  wire          io_inputs_2_payload_atomic,
  input  wire [11:0]   io_inputs_2_payload_storeId,
  output wire          io_output_valid,
  input  wire          io_output_ready,
  output wire [2:0]    io_output_payload_op,
  output wire [31:0]   io_output_payload_address,
  output wire [1:0]    io_output_payload_size,
  output wire          io_output_payload_load,
  output wire          io_output_payload_store,
  output wire          io_output_payload_atomic,
  output wire [11:0]   io_output_payload_storeId,
  output wire [1:0]    io_chosen,
  output wire [2:0]    io_chosenOH,
  input  wire          clk_cpu,
  input  wire          reset_cpu
);
  localparam LsuL1CmdOpcode_LSU = 3'd0;
  localparam LsuL1CmdOpcode_ACCESS_1 = 3'd1;
  localparam LsuL1CmdOpcode_STORE_BUFFER = 3'd2;
  localparam LsuL1CmdOpcode_FLUSH = 3'd3;
  localparam LsuL1CmdOpcode_PREFETCH = 3'd4;

  wire       [2:0]    _zz__zz_maskProposal_1_1;
  reg        [2:0]    _zz__zz_io_output_payload_op;
  reg        [31:0]   _zz_io_output_payload_address_1;
  reg        [1:0]    _zz_io_output_payload_size;
  reg                 _zz_io_output_payload_load;
  reg                 _zz_io_output_payload_store;
  reg                 _zz_io_output_payload_atomic;
  reg        [11:0]   _zz_io_output_payload_storeId;
  wire                locked;
  wire                maskProposal_0;
  wire                maskProposal_1;
  wire                maskProposal_2;
  reg                 maskLocked_0;
  reg                 maskLocked_1;
  reg                 maskLocked_2;
  wire                maskRouted_0;
  wire                maskRouted_1;
  wire                maskRouted_2;
  wire       [2:0]    _zz_maskProposal_1;
  wire       [2:0]    _zz_maskProposal_1_1;
  wire       [1:0]    _zz_io_output_payload_address;
  wire       [2:0]    _zz_io_output_payload_op;
  wire                _zz_io_chosen;
  wire                _zz_io_chosen_1;
  `ifndef SYNTHESIS
  reg [95:0] io_inputs_0_payload_op_string;
  reg [95:0] io_inputs_1_payload_op_string;
  reg [95:0] io_inputs_2_payload_op_string;
  reg [95:0] io_output_payload_op_string;
  reg [95:0] _zz_io_output_payload_op_string;
  `endif


  assign _zz__zz_maskProposal_1_1 = (_zz_maskProposal_1 - 3'b001);
  always @(*) begin
    case(_zz_io_output_payload_address)
      2'b00 : begin
        _zz__zz_io_output_payload_op = io_inputs_0_payload_op;
        _zz_io_output_payload_address_1 = io_inputs_0_payload_address;
        _zz_io_output_payload_size = io_inputs_0_payload_size;
        _zz_io_output_payload_load = io_inputs_0_payload_load;
        _zz_io_output_payload_store = io_inputs_0_payload_store;
        _zz_io_output_payload_atomic = io_inputs_0_payload_atomic;
        _zz_io_output_payload_storeId = io_inputs_0_payload_storeId;
      end
      2'b01 : begin
        _zz__zz_io_output_payload_op = io_inputs_1_payload_op;
        _zz_io_output_payload_address_1 = io_inputs_1_payload_address;
        _zz_io_output_payload_size = io_inputs_1_payload_size;
        _zz_io_output_payload_load = io_inputs_1_payload_load;
        _zz_io_output_payload_store = io_inputs_1_payload_store;
        _zz_io_output_payload_atomic = io_inputs_1_payload_atomic;
        _zz_io_output_payload_storeId = io_inputs_1_payload_storeId;
      end
      default : begin
        _zz__zz_io_output_payload_op = io_inputs_2_payload_op;
        _zz_io_output_payload_address_1 = io_inputs_2_payload_address;
        _zz_io_output_payload_size = io_inputs_2_payload_size;
        _zz_io_output_payload_load = io_inputs_2_payload_load;
        _zz_io_output_payload_store = io_inputs_2_payload_store;
        _zz_io_output_payload_atomic = io_inputs_2_payload_atomic;
        _zz_io_output_payload_storeId = io_inputs_2_payload_storeId;
      end
    endcase
  end

  `ifndef SYNTHESIS
  always @(*) begin
    case(io_inputs_0_payload_op)
      LsuL1CmdOpcode_LSU : io_inputs_0_payload_op_string = "LSU         ";
      LsuL1CmdOpcode_ACCESS_1 : io_inputs_0_payload_op_string = "ACCESS_1    ";
      LsuL1CmdOpcode_STORE_BUFFER : io_inputs_0_payload_op_string = "STORE_BUFFER";
      LsuL1CmdOpcode_FLUSH : io_inputs_0_payload_op_string = "FLUSH       ";
      LsuL1CmdOpcode_PREFETCH : io_inputs_0_payload_op_string = "PREFETCH    ";
      default : io_inputs_0_payload_op_string = "????????????";
    endcase
  end
  always @(*) begin
    case(io_inputs_1_payload_op)
      LsuL1CmdOpcode_LSU : io_inputs_1_payload_op_string = "LSU         ";
      LsuL1CmdOpcode_ACCESS_1 : io_inputs_1_payload_op_string = "ACCESS_1    ";
      LsuL1CmdOpcode_STORE_BUFFER : io_inputs_1_payload_op_string = "STORE_BUFFER";
      LsuL1CmdOpcode_FLUSH : io_inputs_1_payload_op_string = "FLUSH       ";
      LsuL1CmdOpcode_PREFETCH : io_inputs_1_payload_op_string = "PREFETCH    ";
      default : io_inputs_1_payload_op_string = "????????????";
    endcase
  end
  always @(*) begin
    case(io_inputs_2_payload_op)
      LsuL1CmdOpcode_LSU : io_inputs_2_payload_op_string = "LSU         ";
      LsuL1CmdOpcode_ACCESS_1 : io_inputs_2_payload_op_string = "ACCESS_1    ";
      LsuL1CmdOpcode_STORE_BUFFER : io_inputs_2_payload_op_string = "STORE_BUFFER";
      LsuL1CmdOpcode_FLUSH : io_inputs_2_payload_op_string = "FLUSH       ";
      LsuL1CmdOpcode_PREFETCH : io_inputs_2_payload_op_string = "PREFETCH    ";
      default : io_inputs_2_payload_op_string = "????????????";
    endcase
  end
  always @(*) begin
    case(io_output_payload_op)
      LsuL1CmdOpcode_LSU : io_output_payload_op_string = "LSU         ";
      LsuL1CmdOpcode_ACCESS_1 : io_output_payload_op_string = "ACCESS_1    ";
      LsuL1CmdOpcode_STORE_BUFFER : io_output_payload_op_string = "STORE_BUFFER";
      LsuL1CmdOpcode_FLUSH : io_output_payload_op_string = "FLUSH       ";
      LsuL1CmdOpcode_PREFETCH : io_output_payload_op_string = "PREFETCH    ";
      default : io_output_payload_op_string = "????????????";
    endcase
  end
  always @(*) begin
    case(_zz_io_output_payload_op)
      LsuL1CmdOpcode_LSU : _zz_io_output_payload_op_string = "LSU         ";
      LsuL1CmdOpcode_ACCESS_1 : _zz_io_output_payload_op_string = "ACCESS_1    ";
      LsuL1CmdOpcode_STORE_BUFFER : _zz_io_output_payload_op_string = "STORE_BUFFER";
      LsuL1CmdOpcode_FLUSH : _zz_io_output_payload_op_string = "FLUSH       ";
      LsuL1CmdOpcode_PREFETCH : _zz_io_output_payload_op_string = "PREFETCH    ";
      default : _zz_io_output_payload_op_string = "????????????";
    endcase
  end
  `endif

  assign locked = 1'b0;
  assign maskRouted_0 = (locked ? maskLocked_0 : maskProposal_0);
  assign maskRouted_1 = (locked ? maskLocked_1 : maskProposal_1);
  assign maskRouted_2 = (locked ? maskLocked_2 : maskProposal_2);
  assign _zz_maskProposal_1 = {io_inputs_2_valid,{io_inputs_1_valid,io_inputs_0_valid}};
  assign _zz_maskProposal_1_1 = (_zz_maskProposal_1 & (~ _zz__zz_maskProposal_1_1));
  assign maskProposal_0 = io_inputs_0_valid;
  assign maskProposal_1 = _zz_maskProposal_1_1[1];
  assign maskProposal_2 = _zz_maskProposal_1_1[2];
  assign io_output_valid = (((io_inputs_0_valid && maskRouted_0) || (io_inputs_1_valid && maskRouted_1)) || (io_inputs_2_valid && maskRouted_2));
  assign _zz_io_output_payload_address = {maskRouted_2,maskRouted_1};
  assign _zz_io_output_payload_op = _zz__zz_io_output_payload_op;
  assign io_output_payload_op = _zz_io_output_payload_op;
  assign io_output_payload_address = _zz_io_output_payload_address_1;
  assign io_output_payload_size = _zz_io_output_payload_size;
  assign io_output_payload_load = _zz_io_output_payload_load;
  assign io_output_payload_store = _zz_io_output_payload_store;
  assign io_output_payload_atomic = _zz_io_output_payload_atomic;
  assign io_output_payload_storeId = _zz_io_output_payload_storeId;
  assign io_inputs_0_ready = (maskRouted_0 && io_output_ready);
  assign io_inputs_1_ready = (maskRouted_1 && io_output_ready);
  assign io_inputs_2_ready = (maskRouted_2 && io_output_ready);
  assign io_chosenOH = {maskRouted_2,{maskRouted_1,maskRouted_0}};
  assign _zz_io_chosen = io_chosenOH[1];
  assign _zz_io_chosen_1 = io_chosenOH[2];
  assign io_chosen = {_zz_io_chosen_1,_zz_io_chosen};
  always @(posedge clk_cpu) begin
    if(io_output_valid) begin
      maskLocked_0 <= maskRouted_0;
      maskLocked_1 <= maskRouted_1;
      maskLocked_2 <= maskRouted_2;
    end
  end


endmodule

module StreamArbiter_1 (
  input  wire          io_inputs_0_valid,
  output wire          io_inputs_0_ready,
  input  wire [31:0]   io_inputs_0_payload_pcOnLastSlice,
  input  wire [31:0]   io_inputs_0_payload_pcTarget,
  input  wire          io_inputs_0_payload_taken,
  input  wire          io_inputs_0_payload_isBranch,
  input  wire          io_inputs_0_payload_isPush,
  input  wire          io_inputs_0_payload_isPop,
  input  wire          io_inputs_0_payload_wasWrong,
  input  wire          io_inputs_0_payload_badPredictedTarget,
  input  wire [11:0]   io_inputs_0_payload_history,
  input  wire [15:0]   io_inputs_0_payload_uopId,
  input  wire [1:0]    io_inputs_0_payload_ctx_GSharePlugin_GSHARE_COUNTER_0,
  input  wire [1:0]    io_inputs_0_payload_ctx_GSharePlugin_GSHARE_COUNTER_1,
  input  wire [1:0]    io_inputs_0_payload_ctx_GSharePlugin_GSHARE_COUNTER_2,
  input  wire [1:0]    io_inputs_0_payload_ctx_GSharePlugin_GSHARE_COUNTER_3,
  input  wire          io_inputs_1_valid,
  output wire          io_inputs_1_ready,
  input  wire [31:0]   io_inputs_1_payload_pcOnLastSlice,
  input  wire [31:0]   io_inputs_1_payload_pcTarget,
  input  wire          io_inputs_1_payload_taken,
  input  wire          io_inputs_1_payload_isBranch,
  input  wire          io_inputs_1_payload_isPush,
  input  wire          io_inputs_1_payload_isPop,
  input  wire          io_inputs_1_payload_wasWrong,
  input  wire          io_inputs_1_payload_badPredictedTarget,
  input  wire [11:0]   io_inputs_1_payload_history,
  input  wire [15:0]   io_inputs_1_payload_uopId,
  input  wire [1:0]    io_inputs_1_payload_ctx_GSharePlugin_GSHARE_COUNTER_0,
  input  wire [1:0]    io_inputs_1_payload_ctx_GSharePlugin_GSHARE_COUNTER_1,
  input  wire [1:0]    io_inputs_1_payload_ctx_GSharePlugin_GSHARE_COUNTER_2,
  input  wire [1:0]    io_inputs_1_payload_ctx_GSharePlugin_GSHARE_COUNTER_3,
  output wire          io_output_valid,
  input  wire          io_output_ready,
  output wire [31:0]   io_output_payload_pcOnLastSlice,
  output wire [31:0]   io_output_payload_pcTarget,
  output wire          io_output_payload_taken,
  output wire          io_output_payload_isBranch,
  output wire          io_output_payload_isPush,
  output wire          io_output_payload_isPop,
  output wire          io_output_payload_wasWrong,
  output wire          io_output_payload_badPredictedTarget,
  output wire [11:0]   io_output_payload_history,
  output wire [15:0]   io_output_payload_uopId,
  output wire [1:0]    io_output_payload_ctx_GSharePlugin_GSHARE_COUNTER_0,
  output wire [1:0]    io_output_payload_ctx_GSharePlugin_GSHARE_COUNTER_1,
  output wire [1:0]    io_output_payload_ctx_GSharePlugin_GSHARE_COUNTER_2,
  output wire [1:0]    io_output_payload_ctx_GSharePlugin_GSHARE_COUNTER_3,
  output wire [0:0]    io_chosen,
  output wire [1:0]    io_chosenOH,
  input  wire          clk_cpu,
  input  wire          reset_cpu
);

  wire       [3:0]    _zz__zz_maskProposal_0_2;
  wire       [3:0]    _zz__zz_maskProposal_0_2_1;
  wire       [1:0]    _zz__zz_maskProposal_0_2_2;
  wire                locked;
  wire                maskProposal_0;
  wire                maskProposal_1;
  reg                 maskLocked_0;
  reg                 maskLocked_1;
  wire                maskRouted_0;
  wire                maskRouted_1;
  wire       [1:0]    _zz_maskProposal_0;
  wire       [3:0]    _zz_maskProposal_0_1;
  wire       [3:0]    _zz_maskProposal_0_2;
  wire       [1:0]    _zz_maskProposal_0_3;
  wire                _zz_io_chosen;

  assign _zz__zz_maskProposal_0_2 = (_zz_maskProposal_0_1 - _zz__zz_maskProposal_0_2_1);
  assign _zz__zz_maskProposal_0_2_2 = {maskLocked_0,maskLocked_1};
  assign _zz__zz_maskProposal_0_2_1 = {2'd0, _zz__zz_maskProposal_0_2_2};
  assign locked = 1'b0;
  assign maskRouted_0 = (locked ? maskLocked_0 : maskProposal_0);
  assign maskRouted_1 = (locked ? maskLocked_1 : maskProposal_1);
  assign _zz_maskProposal_0 = {io_inputs_1_valid,io_inputs_0_valid};
  assign _zz_maskProposal_0_1 = {_zz_maskProposal_0,_zz_maskProposal_0};
  assign _zz_maskProposal_0_2 = (_zz_maskProposal_0_1 & (~ _zz__zz_maskProposal_0_2));
  assign _zz_maskProposal_0_3 = (_zz_maskProposal_0_2[3 : 2] | _zz_maskProposal_0_2[1 : 0]);
  assign maskProposal_0 = _zz_maskProposal_0_3[0];
  assign maskProposal_1 = _zz_maskProposal_0_3[1];
  assign io_output_valid = ((io_inputs_0_valid && maskRouted_0) || (io_inputs_1_valid && maskRouted_1));
  assign io_output_payload_pcOnLastSlice = (maskRouted_0 ? io_inputs_0_payload_pcOnLastSlice : io_inputs_1_payload_pcOnLastSlice);
  assign io_output_payload_pcTarget = (maskRouted_0 ? io_inputs_0_payload_pcTarget : io_inputs_1_payload_pcTarget);
  assign io_output_payload_taken = (maskRouted_0 ? io_inputs_0_payload_taken : io_inputs_1_payload_taken);
  assign io_output_payload_isBranch = (maskRouted_0 ? io_inputs_0_payload_isBranch : io_inputs_1_payload_isBranch);
  assign io_output_payload_isPush = (maskRouted_0 ? io_inputs_0_payload_isPush : io_inputs_1_payload_isPush);
  assign io_output_payload_isPop = (maskRouted_0 ? io_inputs_0_payload_isPop : io_inputs_1_payload_isPop);
  assign io_output_payload_wasWrong = (maskRouted_0 ? io_inputs_0_payload_wasWrong : io_inputs_1_payload_wasWrong);
  assign io_output_payload_badPredictedTarget = (maskRouted_0 ? io_inputs_0_payload_badPredictedTarget : io_inputs_1_payload_badPredictedTarget);
  assign io_output_payload_history = (maskRouted_0 ? io_inputs_0_payload_history : io_inputs_1_payload_history);
  assign io_output_payload_uopId = (maskRouted_0 ? io_inputs_0_payload_uopId : io_inputs_1_payload_uopId);
  assign io_output_payload_ctx_GSharePlugin_GSHARE_COUNTER_0 = (maskRouted_0 ? io_inputs_0_payload_ctx_GSharePlugin_GSHARE_COUNTER_0 : io_inputs_1_payload_ctx_GSharePlugin_GSHARE_COUNTER_0);
  assign io_output_payload_ctx_GSharePlugin_GSHARE_COUNTER_1 = (maskRouted_0 ? io_inputs_0_payload_ctx_GSharePlugin_GSHARE_COUNTER_1 : io_inputs_1_payload_ctx_GSharePlugin_GSHARE_COUNTER_1);
  assign io_output_payload_ctx_GSharePlugin_GSHARE_COUNTER_2 = (maskRouted_0 ? io_inputs_0_payload_ctx_GSharePlugin_GSHARE_COUNTER_2 : io_inputs_1_payload_ctx_GSharePlugin_GSHARE_COUNTER_2);
  assign io_output_payload_ctx_GSharePlugin_GSHARE_COUNTER_3 = (maskRouted_0 ? io_inputs_0_payload_ctx_GSharePlugin_GSHARE_COUNTER_3 : io_inputs_1_payload_ctx_GSharePlugin_GSHARE_COUNTER_3);
  assign io_inputs_0_ready = (maskRouted_0 && io_output_ready);
  assign io_inputs_1_ready = (maskRouted_1 && io_output_ready);
  assign io_chosenOH = {maskRouted_1,maskRouted_0};
  assign _zz_io_chosen = io_chosenOH[1];
  assign io_chosen = _zz_io_chosen;
  always @(posedge clk_cpu or posedge reset_cpu) begin
    if(reset_cpu) begin
      maskLocked_0 <= 1'b0;
      maskLocked_1 <= 1'b1;
    end else begin
      if(io_output_valid) begin
        maskLocked_0 <= maskRouted_0;
        maskLocked_1 <= maskRouted_1;
      end
    end
  end


endmodule

module StreamArbiter (
  input  wire          io_inputs_0_valid,
  output wire          io_inputs_0_ready,
  output wire          io_output_valid,
  input  wire          io_output_ready,
  output wire [0:0]    io_chosenOH,
  input  wire          clk_cpu,
  input  wire          reset_cpu
);

  reg                 locked;
  wire                maskProposal_0;
  reg                 maskLocked_0;
  wire                maskRouted_0;
  wire                io_output_fire;

  assign maskRouted_0 = (locked ? maskLocked_0 : maskProposal_0);
  assign maskProposal_0 = io_inputs_0_valid;
  assign io_output_fire = (io_output_valid && io_output_ready);
  assign io_output_valid = (io_inputs_0_valid && maskRouted_0);
  assign io_inputs_0_ready = (maskRouted_0 && io_output_ready);
  assign io_chosenOH = maskRouted_0;
  always @(posedge clk_cpu or posedge reset_cpu) begin
    if(reset_cpu) begin
      locked <= 1'b0;
    end else begin
      if(io_output_valid) begin
        locked <= 1'b1;
      end
      if(io_output_fire) begin
        locked <= 1'b0;
      end
    end
  end

  always @(posedge clk_cpu) begin
    if(io_output_valid) begin
      maskLocked_0 <= maskRouted_0;
    end
  end


endmodule

module DivRadix (
  input  wire          io_flush,
  input  wire          io_cmd_valid,
  output wire          io_cmd_ready,
  input  wire [31:0]   io_cmd_payload_a,
  input  wire [31:0]   io_cmd_payload_b,
  input  wire          io_cmd_payload_normalized,
  input  wire [4:0]    io_cmd_payload_iterations,
  output wire          io_rsp_valid,
  input  wire          io_rsp_ready,
  output wire [31:0]   io_rsp_payload_result,
  output wire [31:0]   io_rsp_payload_remain,
  input  wire          clk_cpu,
  input  wire          reset_cpu
);

  wire       [7:0]    _zz_shifter_1;
  wire       [15:0]   _zz_shifter_2;
  wire       [23:0]   _zz_shifter_3;
  wire       [30:0]   _zz_shifter_4;
  reg        [4:0]    counter;
  reg                 busy;
  wire                io_rsp_fire;
  reg                 done;
  wire                when_DivRadix_l41;
  reg        [31:0]   shifter;
  reg        [31:0]   numerator;
  reg        [31:0]   result;
  reg        [32:0]   div1;
  reg        [32:0]   div3;
  wire       [32:0]   div2;
  wire       [32:0]   shifted;
  wire       [33:0]   sub1;
  wire                when_DivRadix_l60;
  reg        [32:0]   _zz_shifter;
  wire                when_DivRadix_l64;
  wire                slicesZero_0;
  wire                slicesZero_1;
  wire                slicesZero_2;
  wire       [2:0]    shiftSel;
  wire       [3:0]    _zz_sel;
  wire                _zz_sel_1;
  wire                _zz_sel_2;
  wire                _zz_sel_3;
  reg        [3:0]    _zz_sel_4;
  wire       [3:0]    _zz_sel_5;
  wire                _zz_sel_6;
  wire                _zz_sel_7;
  wire                _zz_sel_8;
  wire       [1:0]    sel;
  reg                 wasBusy;
  wire                when_DivRadix_l89;

  assign _zz_shifter_1 = io_cmd_payload_a[31 : 24];
  assign _zz_shifter_2 = io_cmd_payload_a[31 : 16];
  assign _zz_shifter_3 = io_cmd_payload_a[31 : 8];
  assign _zz_shifter_4 = io_cmd_payload_a[31 : 1];
  assign io_rsp_fire = (io_rsp_valid && io_rsp_ready);
  assign when_DivRadix_l41 = (busy && (counter == 5'h1f));
  assign div2 = (div1 <<< 1);
  assign shifted = {shifter,numerator[31 : 31]};
  assign sub1 = ({1'b0,shifted} - {1'b0,div1});
  assign io_rsp_valid = done;
  assign io_rsp_payload_result = result;
  assign io_rsp_payload_remain = shifter;
  assign io_cmd_ready = (! busy);
  assign when_DivRadix_l60 = (! done);
  always @(*) begin
    _zz_shifter = shifted;
    if(when_DivRadix_l64) begin
      _zz_shifter = sub1[32:0];
    end
  end

  assign when_DivRadix_l64 = (! sub1[33]);
  assign slicesZero_0 = (io_cmd_payload_a[15 : 8] == 8'h0);
  assign slicesZero_1 = (io_cmd_payload_a[23 : 16] == 8'h0);
  assign slicesZero_2 = (io_cmd_payload_a[31 : 24] == 8'h0);
  assign shiftSel = {(&slicesZero_2),{(&{slicesZero_2,slicesZero_1}),(&{slicesZero_2,{slicesZero_1,slicesZero_0}})}};
  assign _zz_sel = {1'b1,shiftSel};
  assign _zz_sel_1 = _zz_sel[0];
  assign _zz_sel_2 = _zz_sel[1];
  assign _zz_sel_3 = _zz_sel[2];
  always @(*) begin
    _zz_sel_4[0] = (_zz_sel_1 && (! 1'b0));
    _zz_sel_4[1] = (_zz_sel_2 && (! _zz_sel_1));
    _zz_sel_4[2] = (_zz_sel_3 && (! (|{_zz_sel_2,_zz_sel_1})));
    _zz_sel_4[3] = (_zz_sel[3] && (! (|{_zz_sel_3,{_zz_sel_2,_zz_sel_1}})));
  end

  assign _zz_sel_5 = _zz_sel_4;
  assign _zz_sel_6 = _zz_sel_5[3];
  assign _zz_sel_7 = (_zz_sel_5[1] || _zz_sel_6);
  assign _zz_sel_8 = (_zz_sel_5[2] || _zz_sel_6);
  assign sel = {_zz_sel_8,_zz_sel_7};
  assign when_DivRadix_l89 = (! busy);
  always @(posedge clk_cpu or posedge reset_cpu) begin
    if(reset_cpu) begin
      busy <= 1'b0;
      done <= 1'b0;
      wasBusy <= 1'b0;
    end else begin
      if(io_rsp_fire) begin
        busy <= 1'b0;
      end
      if(when_DivRadix_l41) begin
        done <= 1'b1;
      end
      if(io_rsp_fire) begin
        done <= 1'b0;
      end
      wasBusy <= busy;
      if(when_DivRadix_l89) begin
        busy <= io_cmd_valid;
      end
      if(io_flush) begin
        done <= 1'b0;
        busy <= 1'b0;
      end
    end
  end

  always @(posedge clk_cpu) begin
    if(when_DivRadix_l60) begin
      counter <= (counter + 5'h01);
      result <= (result <<< 1);
      if(when_DivRadix_l64) begin
        result[0 : 0] <= 1'b1;
      end
      shifter <= _zz_shifter[31:0];
      numerator <= (numerator <<< 1);
    end
    if(when_DivRadix_l89) begin
      div1 <= {1'd0, io_cmd_payload_b};
      result <= ((io_cmd_payload_b == 32'h0) ? 32'hffffffff : 32'h0);
      case(sel)
        2'b11 : begin
          counter <= 5'h0;
          shifter <= 32'h0;
          numerator <= (io_cmd_payload_a <<< 0);
        end
        2'b10 : begin
          counter <= 5'h08;
          shifter <= {24'd0, _zz_shifter_1};
          numerator <= (io_cmd_payload_a <<< 8);
        end
        2'b01 : begin
          counter <= 5'h10;
          shifter <= {16'd0, _zz_shifter_2};
          numerator <= (io_cmd_payload_a <<< 16);
        end
        default : begin
          counter <= 5'h18;
          shifter <= {8'd0, _zz_shifter_3};
          numerator <= (io_cmd_payload_a <<< 24);
        end
      endcase
      if(io_cmd_payload_normalized) begin
        counter <= (5'h1f - io_cmd_payload_iterations);
        shifter <= {1'd0, _zz_shifter_4};
        numerator <= (io_cmd_payload_a <<< 31);
      end
    end
  end


endmodule

module BmbOnChipRamMultiPort (
  input  wire          io_buses_0_cmd_valid,
  output wire          io_buses_0_cmd_ready,
  input  wire          io_buses_0_cmd_payload_last,
  input  wire [0:0]    io_buses_0_cmd_payload_fragment_opcode,
  input  wire [11:0]   io_buses_0_cmd_payload_fragment_address,
  input  wire [5:0]    io_buses_0_cmd_payload_fragment_length,
  input  wire [31:0]   io_buses_0_cmd_payload_fragment_data,
  input  wire [3:0]    io_buses_0_cmd_payload_fragment_mask,
  output wire          io_buses_0_rsp_valid,
  input  wire          io_buses_0_rsp_ready,
  output wire          io_buses_0_rsp_payload_last,
  output wire [0:0]    io_buses_0_rsp_payload_fragment_opcode,
  output wire [31:0]   io_buses_0_rsp_payload_fragment_data,
  input  wire          io_buses_1_cmd_valid,
  output wire          io_buses_1_cmd_ready,
  input  wire          io_buses_1_cmd_payload_last,
  input  wire [0:0]    io_buses_1_cmd_payload_fragment_opcode,
  input  wire [11:0]   io_buses_1_cmd_payload_fragment_address,
  input  wire [1:0]    io_buses_1_cmd_payload_fragment_length,
  input  wire [31:0]   io_buses_1_cmd_payload_fragment_data,
  input  wire [3:0]    io_buses_1_cmd_payload_fragment_mask,
  output wire          io_buses_1_rsp_valid,
  input  wire          io_buses_1_rsp_ready,
  output wire          io_buses_1_rsp_payload_last,
  output wire [0:0]    io_buses_1_rsp_payload_fragment_opcode,
  output wire [31:0]   io_buses_1_rsp_payload_fragment_data,
  input  wire          clk_peripheral,
  input  wire          reset_peripheral
);

  reg        [31:0]   ram_1_spinal_port0;
  reg        [31:0]   ram_1_spinal_port2;
  wire                _zz_ram_1_port;
  wire                _zz_io_buses_0_rsp_payload_fragment_data_2;
  wire                _zz_ram_1_port_1;
  wire                _zz_ram_1_port_2;
  wire                _zz_io_buses_1_rsp_payload_fragment_data_2;
  wire                _zz_ram_1_port_3;
  reg        [9:0]    _zz_io_buses_0_rsp_payload_fragment_data;
  wire                io_buses_0_cmd_fire;
  reg        [9:0]    _zz_io_buses_0_rsp_payload_fragment_data_1;
  wire                io_buses_0_cmd_isStall;
  wire                io_buses_0_rsp_isStall;
  reg                 io_buses_0_cmd_valid_regNextWhen;
  reg        [9:0]    _zz_io_buses_1_rsp_payload_fragment_data;
  wire                io_buses_1_cmd_fire;
  reg        [9:0]    _zz_io_buses_1_rsp_payload_fragment_data_1;
  wire                io_buses_1_cmd_isStall;
  wire                io_buses_1_rsp_isStall;
  reg                 io_buses_1_cmd_valid_regNextWhen;
  reg [7:0] ram_1_symbol0 [0:1023];
  reg [7:0] ram_1_symbol1 [0:1023];
  reg [7:0] ram_1_symbol2 [0:1023];
  reg [7:0] ram_1_symbol3 [0:1023];
  reg [7:0] _zz_ram_1symbol_read;
  reg [7:0] _zz_ram_1symbol_read_1;
  reg [7:0] _zz_ram_1symbol_read_2;
  reg [7:0] _zz_ram_1symbol_read_3;
  reg [7:0] _zz_ram_1symbol_read_4;
  reg [7:0] _zz_ram_1symbol_read_5;
  reg [7:0] _zz_ram_1symbol_read_6;
  reg [7:0] _zz_ram_1symbol_read_7;

  assign _zz_io_buses_0_rsp_payload_fragment_data_2 = 1'b1;
  assign _zz_ram_1_port_1 = (io_buses_0_cmd_fire && (io_buses_0_cmd_payload_fragment_opcode == 1'b1));
  assign _zz_io_buses_1_rsp_payload_fragment_data_2 = 1'b1;
  assign _zz_ram_1_port_3 = (io_buses_1_cmd_fire && (io_buses_1_cmd_payload_fragment_opcode == 1'b1));
  always @(*) begin
    ram_1_spinal_port0 = {_zz_ram_1symbol_read_3, _zz_ram_1symbol_read_2, _zz_ram_1symbol_read_1, _zz_ram_1symbol_read};
  end
  always @(*) begin
    ram_1_spinal_port2 = {_zz_ram_1symbol_read_7, _zz_ram_1symbol_read_6, _zz_ram_1symbol_read_5, _zz_ram_1symbol_read_4};
  end
  always @(posedge clk_peripheral) begin
    if(_zz_io_buses_0_rsp_payload_fragment_data_2) begin
      _zz_ram_1symbol_read <= ram_1_symbol0[_zz_io_buses_0_rsp_payload_fragment_data];
      _zz_ram_1symbol_read_1 <= ram_1_symbol1[_zz_io_buses_0_rsp_payload_fragment_data];
      _zz_ram_1symbol_read_2 <= ram_1_symbol2[_zz_io_buses_0_rsp_payload_fragment_data];
      _zz_ram_1symbol_read_3 <= ram_1_symbol3[_zz_io_buses_0_rsp_payload_fragment_data];
    end
  end

  always @(posedge clk_peripheral) begin
    if(io_buses_0_cmd_payload_fragment_mask[0] && _zz_ram_1_port_1) begin
      ram_1_symbol0[_zz_io_buses_0_rsp_payload_fragment_data] <= io_buses_0_cmd_payload_fragment_data[7 : 0];
    end
    if(io_buses_0_cmd_payload_fragment_mask[1] && _zz_ram_1_port_1) begin
      ram_1_symbol1[_zz_io_buses_0_rsp_payload_fragment_data] <= io_buses_0_cmd_payload_fragment_data[15 : 8];
    end
    if(io_buses_0_cmd_payload_fragment_mask[2] && _zz_ram_1_port_1) begin
      ram_1_symbol2[_zz_io_buses_0_rsp_payload_fragment_data] <= io_buses_0_cmd_payload_fragment_data[23 : 16];
    end
    if(io_buses_0_cmd_payload_fragment_mask[3] && _zz_ram_1_port_1) begin
      ram_1_symbol3[_zz_io_buses_0_rsp_payload_fragment_data] <= io_buses_0_cmd_payload_fragment_data[31 : 24];
    end
  end

  always @(posedge clk_peripheral) begin
    if(_zz_io_buses_1_rsp_payload_fragment_data_2) begin
      _zz_ram_1symbol_read_4 <= ram_1_symbol0[_zz_io_buses_1_rsp_payload_fragment_data];
      _zz_ram_1symbol_read_5 <= ram_1_symbol1[_zz_io_buses_1_rsp_payload_fragment_data];
      _zz_ram_1symbol_read_6 <= ram_1_symbol2[_zz_io_buses_1_rsp_payload_fragment_data];
      _zz_ram_1symbol_read_7 <= ram_1_symbol3[_zz_io_buses_1_rsp_payload_fragment_data];
    end
  end

  always @(posedge clk_peripheral) begin
    if(io_buses_1_cmd_payload_fragment_mask[0] && _zz_ram_1_port_3) begin
      ram_1_symbol0[_zz_io_buses_1_rsp_payload_fragment_data] <= io_buses_1_cmd_payload_fragment_data[7 : 0];
    end
    if(io_buses_1_cmd_payload_fragment_mask[1] && _zz_ram_1_port_3) begin
      ram_1_symbol1[_zz_io_buses_1_rsp_payload_fragment_data] <= io_buses_1_cmd_payload_fragment_data[15 : 8];
    end
    if(io_buses_1_cmd_payload_fragment_mask[2] && _zz_ram_1_port_3) begin
      ram_1_symbol2[_zz_io_buses_1_rsp_payload_fragment_data] <= io_buses_1_cmd_payload_fragment_data[23 : 16];
    end
    if(io_buses_1_cmd_payload_fragment_mask[3] && _zz_ram_1_port_3) begin
      ram_1_symbol3[_zz_io_buses_1_rsp_payload_fragment_data] <= io_buses_1_cmd_payload_fragment_data[31 : 24];
    end
  end

  always @(*) begin
    _zz_io_buses_0_rsp_payload_fragment_data = (io_buses_0_cmd_payload_fragment_address >>> 2'd2);
    if(io_buses_0_cmd_isStall) begin
      _zz_io_buses_0_rsp_payload_fragment_data = _zz_io_buses_0_rsp_payload_fragment_data_1;
    end
  end

  assign io_buses_0_cmd_fire = (io_buses_0_cmd_valid && io_buses_0_cmd_ready);
  assign io_buses_0_cmd_isStall = (io_buses_0_cmd_valid && (! io_buses_0_cmd_ready));
  assign io_buses_0_rsp_isStall = (io_buses_0_rsp_valid && (! io_buses_0_rsp_ready));
  assign io_buses_0_cmd_ready = (! io_buses_0_rsp_isStall);
  assign io_buses_0_rsp_valid = io_buses_0_cmd_valid_regNextWhen;
  assign io_buses_0_rsp_payload_fragment_data = ram_1_spinal_port0;
  assign io_buses_0_rsp_payload_fragment_opcode = 1'b0;
  assign io_buses_0_rsp_payload_last = 1'b1;
  always @(*) begin
    _zz_io_buses_1_rsp_payload_fragment_data = (io_buses_1_cmd_payload_fragment_address >>> 2'd2);
    if(io_buses_1_cmd_isStall) begin
      _zz_io_buses_1_rsp_payload_fragment_data = _zz_io_buses_1_rsp_payload_fragment_data_1;
    end
  end

  assign io_buses_1_cmd_fire = (io_buses_1_cmd_valid && io_buses_1_cmd_ready);
  assign io_buses_1_cmd_isStall = (io_buses_1_cmd_valid && (! io_buses_1_cmd_ready));
  assign io_buses_1_rsp_isStall = (io_buses_1_rsp_valid && (! io_buses_1_rsp_ready));
  assign io_buses_1_cmd_ready = (! io_buses_1_rsp_isStall);
  assign io_buses_1_rsp_valid = io_buses_1_cmd_valid_regNextWhen;
  assign io_buses_1_rsp_payload_fragment_data = ram_1_spinal_port2;
  assign io_buses_1_rsp_payload_fragment_opcode = 1'b0;
  assign io_buses_1_rsp_payload_last = 1'b1;
  always @(posedge clk_peripheral) begin
    if(io_buses_0_cmd_fire) begin
      _zz_io_buses_0_rsp_payload_fragment_data_1 <= _zz_io_buses_0_rsp_payload_fragment_data;
    end
    if(io_buses_1_cmd_fire) begin
      _zz_io_buses_1_rsp_payload_fragment_data_1 <= _zz_io_buses_1_rsp_payload_fragment_data;
    end
  end

  always @(posedge clk_peripheral or posedge reset_peripheral) begin
    if(reset_peripheral) begin
      io_buses_0_cmd_valid_regNextWhen <= 1'b0;
      io_buses_1_cmd_valid_regNextWhen <= 1'b0;
    end else begin
      if(io_buses_0_cmd_ready) begin
        io_buses_0_cmd_valid_regNextWhen <= io_buses_0_cmd_valid;
      end
      if(io_buses_1_cmd_ready) begin
        io_buses_1_cmd_valid_regNextWhen <= io_buses_1_cmd_valid;
      end
    end
  end


endmodule

module UsbLsFsPhyModified (
  input  wire          io_ctrl_lowSpeed,
  input  wire          io_ctrl_tx_valid,
  output reg           io_ctrl_tx_ready,
  input  wire          io_ctrl_tx_payload_last,
  input  wire [7:0]    io_ctrl_tx_payload_fragment,
  output reg           io_ctrl_txEop,
  output reg           io_ctrl_rx_flow_valid,
  output reg           io_ctrl_rx_flow_payload_stuffingError,
  output reg  [7:0]    io_ctrl_rx_flow_payload_data,
  output reg           io_ctrl_rx_active,
  input  wire          io_ctrl_usbReset,
  input  wire          io_ctrl_usbResume,
  output wire          io_ctrl_overcurrent,
  output wire          io_ctrl_tick,
  input  wire          io_ctrl_ports_0_disable_valid,
  output wire          io_ctrl_ports_0_disable_ready,
  input  wire          io_ctrl_ports_0_removable,
  input  wire          io_ctrl_ports_0_power,
  input  wire          io_ctrl_ports_0_reset_valid,
  output reg           io_ctrl_ports_0_reset_ready,
  input  wire          io_ctrl_ports_0_suspend_valid,
  output wire          io_ctrl_ports_0_suspend_ready,
  input  wire          io_ctrl_ports_0_resume_valid,
  output wire          io_ctrl_ports_0_resume_ready,
  output reg           io_ctrl_ports_0_connect,
  output wire          io_ctrl_ports_0_disconnect,
  output wire          io_ctrl_ports_0_overcurrent,
  output wire          io_ctrl_ports_0_remoteResume,
  output wire          io_ctrl_ports_0_lowSpeed,
  input  wire          io_ctrl_ports_1_disable_valid,
  output wire          io_ctrl_ports_1_disable_ready,
  input  wire          io_ctrl_ports_1_removable,
  input  wire          io_ctrl_ports_1_power,
  input  wire          io_ctrl_ports_1_reset_valid,
  output reg           io_ctrl_ports_1_reset_ready,
  input  wire          io_ctrl_ports_1_suspend_valid,
  output wire          io_ctrl_ports_1_suspend_ready,
  input  wire          io_ctrl_ports_1_resume_valid,
  output wire          io_ctrl_ports_1_resume_ready,
  output reg           io_ctrl_ports_1_connect,
  output wire          io_ctrl_ports_1_disconnect,
  output wire          io_ctrl_ports_1_overcurrent,
  output wire          io_ctrl_ports_1_remoteResume,
  output wire          io_ctrl_ports_1_lowSpeed,
  output reg           io_usb_0_tx_enable,
  output reg           io_usb_0_tx_data,
  output reg           io_usb_0_tx_se0,
  input  wire          io_usb_0_rx_dp,
  input  wire          io_usb_0_rx_dm,
  output reg           io_usb_1_tx_enable,
  output reg           io_usb_1_tx_data,
  output reg           io_usb_1_tx_se0,
  input  wire          io_usb_1_rx_dp,
  input  wire          io_usb_1_rx_dm,
  input  wire          io_management_0_overcurrent,
  output wire          io_management_0_power,
  input  wire          io_management_1_overcurrent,
  output wire          io_management_1_power,
  input  wire          clk_peripheral,
  input  wire          reset_peripheral
);
  localparam txShared_frame_enumDef_BOOT = 4'd0;
  localparam txShared_frame_enumDef_IDLE = 4'd1;
  localparam txShared_frame_enumDef_TAKE_LINE = 4'd2;
  localparam txShared_frame_enumDef_PREAMBLE_SYNC = 4'd3;
  localparam txShared_frame_enumDef_PREAMBLE_PID = 4'd4;
  localparam txShared_frame_enumDef_PREAMBLE_DELAY = 4'd5;
  localparam txShared_frame_enumDef_SYNC = 4'd6;
  localparam txShared_frame_enumDef_DATA = 4'd7;
  localparam txShared_frame_enumDef_EOP_0 = 4'd8;
  localparam txShared_frame_enumDef_EOP_1 = 4'd9;
  localparam txShared_frame_enumDef_EOP_2 = 4'd10;
  localparam ports_0_fsm_enumDef_BOOT = 4'd0;
  localparam ports_0_fsm_enumDef_POWER_OFF = 4'd1;
  localparam ports_0_fsm_enumDef_DISCONNECTED = 4'd2;
  localparam ports_0_fsm_enumDef_DISABLED = 4'd3;
  localparam ports_0_fsm_enumDef_RESETTING = 4'd4;
  localparam ports_0_fsm_enumDef_RESETTING_DELAY = 4'd5;
  localparam ports_0_fsm_enumDef_RESETTING_SYNC = 4'd6;
  localparam ports_0_fsm_enumDef_ENABLED = 4'd7;
  localparam ports_0_fsm_enumDef_SUSPENDED = 4'd8;
  localparam ports_0_fsm_enumDef_RESUMING = 4'd9;
  localparam ports_0_fsm_enumDef_SEND_EOP_0 = 4'd10;
  localparam ports_0_fsm_enumDef_SEND_EOP_1 = 4'd11;
  localparam ports_0_fsm_enumDef_RESTART_S = 4'd12;
  localparam ports_0_fsm_enumDef_RESTART_E = 4'd13;
  localparam ports_1_fsm_enumDef_BOOT = 4'd0;
  localparam ports_1_fsm_enumDef_POWER_OFF = 4'd1;
  localparam ports_1_fsm_enumDef_DISCONNECTED = 4'd2;
  localparam ports_1_fsm_enumDef_DISABLED = 4'd3;
  localparam ports_1_fsm_enumDef_RESETTING = 4'd4;
  localparam ports_1_fsm_enumDef_RESETTING_DELAY = 4'd5;
  localparam ports_1_fsm_enumDef_RESETTING_SYNC = 4'd6;
  localparam ports_1_fsm_enumDef_ENABLED = 4'd7;
  localparam ports_1_fsm_enumDef_SUSPENDED = 4'd8;
  localparam ports_1_fsm_enumDef_RESUMING = 4'd9;
  localparam ports_1_fsm_enumDef_SEND_EOP_0 = 4'd10;
  localparam ports_1_fsm_enumDef_SEND_EOP_1 = 4'd11;
  localparam ports_1_fsm_enumDef_RESTART_S = 4'd12;
  localparam ports_1_fsm_enumDef_RESTART_E = 4'd13;
  localparam upstreamRx_enumDef_BOOT = 2'd0;
  localparam upstreamRx_enumDef_IDLE = 2'd1;
  localparam upstreamRx_enumDef_SUSPEND = 2'd2;
  localparam ports_0_rx_packet_enumDef_BOOT = 2'd0;
  localparam ports_0_rx_packet_enumDef_IDLE = 2'd1;
  localparam ports_0_rx_packet_enumDef_PACKET = 2'd2;
  localparam ports_0_rx_packet_enumDef_ERRORED = 2'd3;
  localparam ports_1_rx_packet_enumDef_BOOT = 2'd0;
  localparam ports_1_rx_packet_enumDef_IDLE = 2'd1;
  localparam ports_1_rx_packet_enumDef_PACKET = 2'd2;
  localparam ports_1_rx_packet_enumDef_ERRORED = 2'd3;

  wire                ports_0_filter_io_filtred_dp;
  wire                ports_0_filter_io_filtred_dm;
  wire                ports_0_filter_io_filtred_d;
  wire                ports_0_filter_io_filtred_se0;
  wire                ports_0_filter_io_filtred_sample;
  wire                ports_1_filter_io_filtred_dp;
  wire                ports_1_filter_io_filtred_dm;
  wire                ports_1_filter_io_filtred_d;
  wire                ports_1_filter_io_filtred_se0;
  wire                ports_1_filter_io_filtred_sample;
  wire       [1:0]    _zz_tickTimer_counter_valueNext;
  wire       [0:0]    _zz_tickTimer_counter_valueNext_1;
  wire       [9:0]    _zz_txShared_timer_oneCycle;
  wire       [4:0]    _zz_txShared_timer_oneCycle_1;
  wire       [9:0]    _zz_txShared_timer_twoCycle;
  wire       [5:0]    _zz_txShared_timer_twoCycle_1;
  wire       [9:0]    _zz_txShared_timer_fourCycle;
  wire       [7:0]    _zz_txShared_timer_fourCycle_1;
  wire       [8:0]    _zz_txShared_rxToTxDelay_twoCycle;
  wire       [6:0]    _zz_txShared_rxToTxDelay_twoCycle_1;
  wire       [1:0]    _zz_txShared_lowSpeedSof_state;
  wire       [0:0]    _zz_txShared_lowSpeedSof_state_1;
  wire       [6:0]    _zz_when_usbphy_l403;
  wire       [11:0]   _zz_ports_0_rx_packet_errorTimeout_trigger;
  wire       [9:0]    _zz_ports_0_rx_packet_errorTimeout_trigger_1;
  wire       [6:0]    _zz_ports_0_rx_disconnect_counter;
  wire       [0:0]    _zz_ports_0_rx_disconnect_counter_1;
  wire       [23:0]   _zz_ports_0_fsm_timer_ONE_BIT;
  wire       [4:0]    _zz_ports_0_fsm_timer_ONE_BIT_1;
  wire       [23:0]   _zz_ports_0_fsm_timer_TWO_BIT;
  wire       [5:0]    _zz_ports_0_fsm_timer_TWO_BIT_1;
  wire       [6:0]    _zz_when_usbphy_l403_1;
  wire       [11:0]   _zz_ports_1_rx_packet_errorTimeout_trigger;
  wire       [9:0]    _zz_ports_1_rx_packet_errorTimeout_trigger_1;
  wire       [6:0]    _zz_ports_1_rx_disconnect_counter;
  wire       [0:0]    _zz_ports_1_rx_disconnect_counter_1;
  wire       [23:0]   _zz_ports_1_fsm_timer_ONE_BIT;
  wire       [4:0]    _zz_ports_1_fsm_timer_ONE_BIT_1;
  wire       [23:0]   _zz_ports_1_fsm_timer_TWO_BIT;
  wire       [5:0]    _zz_ports_1_fsm_timer_TWO_BIT_1;
  wire                tickTimer_counter_willIncrement;
  wire                tickTimer_counter_willClear;
  reg        [1:0]    tickTimer_counter_valueNext;
  reg        [1:0]    tickTimer_counter_value;
  wire                tickTimer_counter_willOverflowIfInc;
  wire                tickTimer_counter_willOverflow;
  wire                tickTimer_tick;
  reg                 txShared_timer_lowSpeed;
  reg        [9:0]    txShared_timer_counter;
  reg                 txShared_timer_clear;
  wire                txShared_timer_inc;
  wire                txShared_timer_oneCycle;
  wire                txShared_timer_twoCycle;
  wire                txShared_timer_fourCycle;
  reg                 txShared_rxToTxDelay_lowSpeed;
  reg        [8:0]    txShared_rxToTxDelay_counter;
  reg                 txShared_rxToTxDelay_clear;
  wire                txShared_rxToTxDelay_inc;
  wire                txShared_rxToTxDelay_twoCycle;
  reg                 txShared_rxToTxDelay_active;
  reg                 txShared_encoder_input_valid;
  reg                 txShared_encoder_input_ready;
  reg                 txShared_encoder_input_data;
  reg                 txShared_encoder_input_lowSpeed;
  reg                 txShared_encoder_output_valid;
  reg                 txShared_encoder_output_se0;
  reg                 txShared_encoder_output_lowSpeed;
  reg                 txShared_encoder_output_data;
  reg        [2:0]    txShared_encoder_counter;
  reg                 txShared_encoder_state;
  wire                when_usbphy_l91;
  wire                when_usbphy_l96;
  wire                when_usbphy_l110;
  reg                 txShared_serialiser_input_valid;
  reg                 txShared_serialiser_input_ready;
  reg        [7:0]    txShared_serialiser_input_data;
  reg                 txShared_serialiser_input_lowSpeed;
  reg        [2:0]    txShared_serialiser_bitCounter;
  wire                when_usbphy_l136;
  wire                when_usbphy_l142;
  reg        [4:0]    txShared_lowSpeedSof_timer;
  reg        [1:0]    txShared_lowSpeedSof_state;
  reg                 txShared_lowSpeedSof_increment;
  reg                 txShared_lowSpeedSof_overrideEncoder;
  reg                 txShared_encoder_output_valid_regNext;
  wire                when_usbphy_l151;
  wire                when_usbphy_l153;
  wire                io_ctrl_tx_fire;
  reg                 io_ctrl_tx_payload_first;
  wire                when_usbphy_l154;
  wire                when_usbphy_l161;
  wire                txShared_lowSpeedSof_valid;
  wire                txShared_lowSpeedSof_data;
  wire                txShared_lowSpeedSof_se0;
  wire                txShared_frame_wantExit;
  reg                 txShared_frame_wantStart;
  wire                txShared_frame_wantKill;
  wire                txShared_frame_busy;
  reg                 txShared_frame_wasLowSpeed;
  wire                upstreamRx_wantExit;
  reg                 upstreamRx_wantStart;
  wire                upstreamRx_wantKill;
  wire                upstreamRx_timer_lowSpeed;
  reg        [19:0]   upstreamRx_timer_counter;
  reg                 upstreamRx_timer_clear;
  wire                upstreamRx_timer_inc;
  wire                upstreamRx_timer_IDLE_EOI;
  wire                Rx_Suspend;
  reg                 resumeFromPort;
  reg                 ports_0_portLowSpeed;
  reg                 ports_0_rx_enablePackets;
  wire                ports_0_rx_j;
  wire                ports_0_rx_k;
  reg                 ports_0_rx_stuffingError;
  reg                 ports_0_rx_waitSync;
  reg                 ports_0_rx_decoder_state;
  reg                 ports_0_rx_decoder_output_valid;
  reg                 ports_0_rx_decoder_output_payload;
  wire                when_usbphy_l347;
  reg        [2:0]    ports_0_rx_destuffer_counter;
  wire                ports_0_rx_destuffer_unstuffNext;
  wire                ports_0_rx_destuffer_output_valid;
  wire                ports_0_rx_destuffer_output_payload;
  wire                when_usbphy_l368;
  wire                ports_0_rx_history_updated;
  wire                _zz_ports_0_rx_history_value;
  reg                 _zz_ports_0_rx_history_value_1;
  reg                 _zz_ports_0_rx_history_value_2;
  reg                 _zz_ports_0_rx_history_value_3;
  reg                 _zz_ports_0_rx_history_value_4;
  reg                 _zz_ports_0_rx_history_value_5;
  reg                 _zz_ports_0_rx_history_value_6;
  reg                 _zz_ports_0_rx_history_value_7;
  wire       [7:0]    ports_0_rx_history_value;
  wire                ports_0_rx_history_sync_hit;
  wire       [6:0]    ports_0_rx_eop_maxThreshold;
  wire       [5:0]    ports_0_rx_eop_minThreshold;
  reg        [6:0]    ports_0_rx_eop_counter;
  wire                ports_0_rx_eop_maxHit;
  reg                 ports_0_rx_eop_hit;
  wire                when_usbphy_l395;
  wire                when_usbphy_l396;
  wire                when_usbphy_l403;
  wire                ports_0_rx_packet_wantExit;
  reg                 ports_0_rx_packet_wantStart;
  wire                ports_0_rx_packet_wantKill;
  reg        [2:0]    ports_0_rx_packet_counter;
  wire                ports_0_rx_packet_errorTimeout_lowSpeed;
  reg        [11:0]   ports_0_rx_packet_errorTimeout_counter;
  reg                 ports_0_rx_packet_errorTimeout_clear;
  wire                ports_0_rx_packet_errorTimeout_inc;
  wire                ports_0_rx_packet_errorTimeout_trigger;
  reg                 ports_0_rx_packet_errorTimeout_p;
  reg                 ports_0_rx_packet_errorTimeout_n;
  reg        [6:0]    ports_0_rx_disconnect_counter;
  reg                 ports_0_rx_disconnect_clear;
  wire                ports_0_rx_disconnect_hit;
  reg                 ports_0_rx_disconnect_hitLast;
  wire                ports_0_rx_disconnect_event;
  wire                when_usbphy_l475;
  wire                ports_0_fsm_wantExit;
  reg                 ports_0_fsm_wantStart;
  wire                ports_0_fsm_wantKill;
  reg                 ports_0_fsm_timer_lowSpeed;
  reg        [23:0]   ports_0_fsm_timer_counter;
  reg                 ports_0_fsm_timer_clear;
  wire                ports_0_fsm_timer_inc;
  wire                ports_0_fsm_timer_DISCONNECTED_EOI;
  wire                ports_0_fsm_timer_RESET_DELAY;
  wire                ports_0_fsm_timer_RESET_EOI;
  wire                ports_0_fsm_timer_RESUME_EOI;
  wire                ports_0_fsm_timer_RESTART_EOI;
  wire                ports_0_fsm_timer_ONE_BIT;
  wire                ports_0_fsm_timer_TWO_BIT;
  reg                 ports_0_fsm_resetInProgress;
  reg                 ports_0_fsm_lowSpeedEop;
  wire                ports_0_fsm_forceJ;
  wire                when_usbphy_l672;
  reg                 ports_1_portLowSpeed;
  reg                 ports_1_rx_enablePackets;
  wire                ports_1_rx_j;
  wire                ports_1_rx_k;
  reg                 ports_1_rx_stuffingError;
  reg                 ports_1_rx_waitSync;
  reg                 ports_1_rx_decoder_state;
  reg                 ports_1_rx_decoder_output_valid;
  reg                 ports_1_rx_decoder_output_payload;
  wire                when_usbphy_l347_1;
  reg        [2:0]    ports_1_rx_destuffer_counter;
  wire                ports_1_rx_destuffer_unstuffNext;
  wire                ports_1_rx_destuffer_output_valid;
  wire                ports_1_rx_destuffer_output_payload;
  wire                when_usbphy_l368_1;
  wire                ports_1_rx_history_updated;
  wire                _zz_ports_1_rx_history_value;
  reg                 _zz_ports_1_rx_history_value_1;
  reg                 _zz_ports_1_rx_history_value_2;
  reg                 _zz_ports_1_rx_history_value_3;
  reg                 _zz_ports_1_rx_history_value_4;
  reg                 _zz_ports_1_rx_history_value_5;
  reg                 _zz_ports_1_rx_history_value_6;
  reg                 _zz_ports_1_rx_history_value_7;
  wire       [7:0]    ports_1_rx_history_value;
  wire                ports_1_rx_history_sync_hit;
  wire       [6:0]    ports_1_rx_eop_maxThreshold;
  wire       [5:0]    ports_1_rx_eop_minThreshold;
  reg        [6:0]    ports_1_rx_eop_counter;
  wire                ports_1_rx_eop_maxHit;
  reg                 ports_1_rx_eop_hit;
  wire                when_usbphy_l395_1;
  wire                when_usbphy_l396_1;
  wire                when_usbphy_l403_1;
  wire                ports_1_rx_packet_wantExit;
  reg                 ports_1_rx_packet_wantStart;
  wire                ports_1_rx_packet_wantKill;
  reg        [2:0]    ports_1_rx_packet_counter;
  wire                ports_1_rx_packet_errorTimeout_lowSpeed;
  reg        [11:0]   ports_1_rx_packet_errorTimeout_counter;
  reg                 ports_1_rx_packet_errorTimeout_clear;
  wire                ports_1_rx_packet_errorTimeout_inc;
  wire                ports_1_rx_packet_errorTimeout_trigger;
  reg                 ports_1_rx_packet_errorTimeout_p;
  reg                 ports_1_rx_packet_errorTimeout_n;
  reg        [6:0]    ports_1_rx_disconnect_counter;
  reg                 ports_1_rx_disconnect_clear;
  wire                ports_1_rx_disconnect_hit;
  reg                 ports_1_rx_disconnect_hitLast;
  wire                ports_1_rx_disconnect_event;
  wire                when_usbphy_l475_1;
  wire                ports_1_fsm_wantExit;
  reg                 ports_1_fsm_wantStart;
  wire                ports_1_fsm_wantKill;
  reg                 ports_1_fsm_timer_lowSpeed;
  reg        [23:0]   ports_1_fsm_timer_counter;
  reg                 ports_1_fsm_timer_clear;
  wire                ports_1_fsm_timer_inc;
  wire                ports_1_fsm_timer_DISCONNECTED_EOI;
  wire                ports_1_fsm_timer_RESET_DELAY;
  wire                ports_1_fsm_timer_RESET_EOI;
  wire                ports_1_fsm_timer_RESUME_EOI;
  wire                ports_1_fsm_timer_RESTART_EOI;
  wire                ports_1_fsm_timer_ONE_BIT;
  wire                ports_1_fsm_timer_TWO_BIT;
  reg                 ports_1_fsm_resetInProgress;
  reg                 ports_1_fsm_lowSpeedEop;
  wire                ports_1_fsm_forceJ;
  wire                when_usbphy_l672_1;
  reg        [3:0]    txShared_frame_stateReg;
  reg        [3:0]    txShared_frame_stateNext;
  wire                when_usbphy_l191;
  reg        [1:0]    upstreamRx_stateReg;
  reg        [1:0]    upstreamRx_stateNext;
  reg        [1:0]    ports_0_rx_packet_stateReg;
  reg        [1:0]    ports_0_rx_packet_stateNext;
  wire                when_usbphy_l429;
  wire                when_usbphy_l451;
  wire                when_StateMachine_l253;
  wire                when_StateMachine_l253_1;
  reg        [3:0]    ports_0_fsm_stateReg;
  reg        [3:0]    ports_0_fsm_stateNext;
  wire                when_usbphy_l540;
  wire                when_usbphy_l547;
  wire                when_usbphy_l580;
  wire                when_usbphy_l593;
  wire                when_usbphy_l602;
  wire                when_usbphy_l610;
  wire                when_usbphy_l612;
  wire                when_usbphy_l653;
  wire                when_usbphy_l663;
  wire                when_StateMachine_l253_2;
  wire                when_StateMachine_l253_3;
  wire                when_StateMachine_l253_4;
  wire                when_StateMachine_l253_5;
  wire                when_StateMachine_l253_6;
  wire                when_StateMachine_l253_7;
  wire                when_StateMachine_l253_8;
  wire                when_StateMachine_l253_9;
  wire                when_usbphy_l512;
  wire                when_usbphy_l519;
  wire                when_usbphy_l520;
  reg        [1:0]    ports_1_rx_packet_stateReg;
  reg        [1:0]    ports_1_rx_packet_stateNext;
  wire                when_usbphy_l429_1;
  wire                when_usbphy_l451_1;
  wire                when_StateMachine_l253_10;
  wire                when_StateMachine_l253_11;
  reg        [3:0]    ports_1_fsm_stateReg;
  reg        [3:0]    ports_1_fsm_stateNext;
  wire                when_usbphy_l540_1;
  wire                when_usbphy_l547_1;
  wire                when_usbphy_l580_1;
  wire                when_usbphy_l593_1;
  wire                when_usbphy_l602_1;
  wire                when_usbphy_l610_1;
  wire                when_usbphy_l612_1;
  wire                when_usbphy_l653_1;
  wire                when_usbphy_l663_1;
  wire                when_StateMachine_l253_12;
  wire                when_StateMachine_l253_13;
  wire                when_StateMachine_l253_14;
  wire                when_StateMachine_l253_15;
  wire                when_StateMachine_l253_16;
  wire                when_StateMachine_l253_17;
  wire                when_StateMachine_l253_18;
  wire                when_StateMachine_l253_19;
  wire                when_usbphy_l512_1;
  wire                when_usbphy_l519_1;
  wire                when_usbphy_l520_1;
  `ifndef SYNTHESIS
  reg [111:0] txShared_frame_stateReg_string;
  reg [111:0] txShared_frame_stateNext_string;
  reg [55:0] upstreamRx_stateReg_string;
  reg [55:0] upstreamRx_stateNext_string;
  reg [55:0] ports_0_rx_packet_stateReg_string;
  reg [55:0] ports_0_rx_packet_stateNext_string;
  reg [119:0] ports_0_fsm_stateReg_string;
  reg [119:0] ports_0_fsm_stateNext_string;
  reg [55:0] ports_1_rx_packet_stateReg_string;
  reg [55:0] ports_1_rx_packet_stateNext_string;
  reg [119:0] ports_1_fsm_stateReg_string;
  reg [119:0] ports_1_fsm_stateNext_string;
  `endif


  assign _zz_tickTimer_counter_valueNext_1 = tickTimer_counter_willIncrement;
  assign _zz_tickTimer_counter_valueNext = {1'd0, _zz_tickTimer_counter_valueNext_1};
  assign _zz_txShared_timer_oneCycle_1 = (txShared_timer_lowSpeed ? 5'h1f : 5'h03);
  assign _zz_txShared_timer_oneCycle = {5'd0, _zz_txShared_timer_oneCycle_1};
  assign _zz_txShared_timer_twoCycle_1 = (txShared_timer_lowSpeed ? 6'h3f : 6'h07);
  assign _zz_txShared_timer_twoCycle = {4'd0, _zz_txShared_timer_twoCycle_1};
  assign _zz_txShared_timer_fourCycle_1 = (txShared_timer_lowSpeed ? 8'h9f : 8'h13);
  assign _zz_txShared_timer_fourCycle = {2'd0, _zz_txShared_timer_fourCycle_1};
  assign _zz_txShared_rxToTxDelay_twoCycle_1 = (txShared_rxToTxDelay_lowSpeed ? 7'h7f : 7'h0f);
  assign _zz_txShared_rxToTxDelay_twoCycle = {2'd0, _zz_txShared_rxToTxDelay_twoCycle_1};
  assign _zz_txShared_lowSpeedSof_state_1 = txShared_lowSpeedSof_increment;
  assign _zz_txShared_lowSpeedSof_state = {1'd0, _zz_txShared_lowSpeedSof_state_1};
  assign _zz_when_usbphy_l403 = {1'd0, ports_0_rx_eop_minThreshold};
  assign _zz_ports_0_rx_packet_errorTimeout_trigger_1 = (ports_0_rx_packet_errorTimeout_lowSpeed ? 10'h27f : 10'h04f);
  assign _zz_ports_0_rx_packet_errorTimeout_trigger = {2'd0, _zz_ports_0_rx_packet_errorTimeout_trigger_1};
  assign _zz_ports_0_rx_disconnect_counter_1 = (! ports_0_rx_disconnect_hit);
  assign _zz_ports_0_rx_disconnect_counter = {6'd0, _zz_ports_0_rx_disconnect_counter_1};
  assign _zz_ports_0_fsm_timer_ONE_BIT_1 = (ports_0_fsm_timer_lowSpeed ? 5'h1f : 5'h03);
  assign _zz_ports_0_fsm_timer_ONE_BIT = {19'd0, _zz_ports_0_fsm_timer_ONE_BIT_1};
  assign _zz_ports_0_fsm_timer_TWO_BIT_1 = (ports_0_fsm_timer_lowSpeed ? 6'h3f : 6'h07);
  assign _zz_ports_0_fsm_timer_TWO_BIT = {18'd0, _zz_ports_0_fsm_timer_TWO_BIT_1};
  assign _zz_when_usbphy_l403_1 = {1'd0, ports_1_rx_eop_minThreshold};
  assign _zz_ports_1_rx_packet_errorTimeout_trigger_1 = (ports_1_rx_packet_errorTimeout_lowSpeed ? 10'h27f : 10'h04f);
  assign _zz_ports_1_rx_packet_errorTimeout_trigger = {2'd0, _zz_ports_1_rx_packet_errorTimeout_trigger_1};
  assign _zz_ports_1_rx_disconnect_counter_1 = (! ports_1_rx_disconnect_hit);
  assign _zz_ports_1_rx_disconnect_counter = {6'd0, _zz_ports_1_rx_disconnect_counter_1};
  assign _zz_ports_1_fsm_timer_ONE_BIT_1 = (ports_1_fsm_timer_lowSpeed ? 5'h1f : 5'h03);
  assign _zz_ports_1_fsm_timer_ONE_BIT = {19'd0, _zz_ports_1_fsm_timer_ONE_BIT_1};
  assign _zz_ports_1_fsm_timer_TWO_BIT_1 = (ports_1_fsm_timer_lowSpeed ? 6'h3f : 6'h07);
  assign _zz_ports_1_fsm_timer_TWO_BIT = {18'd0, _zz_ports_1_fsm_timer_TWO_BIT_1};
  UsbLsFsPhyFilter ports_0_filter (
    .io_lowSpeed       (io_ctrl_lowSpeed                ), //i
    .io_usb_dp         (io_usb_0_rx_dp                  ), //i
    .io_usb_dm         (io_usb_0_rx_dm                  ), //i
    .io_filtred_dp     (ports_0_filter_io_filtred_dp    ), //o
    .io_filtred_dm     (ports_0_filter_io_filtred_dm    ), //o
    .io_filtred_d      (ports_0_filter_io_filtred_d     ), //o
    .io_filtred_se0    (ports_0_filter_io_filtred_se0   ), //o
    .io_filtred_sample (ports_0_filter_io_filtred_sample), //o
    .clk_peripheral    (clk_peripheral                  ), //i
    .reset_peripheral  (reset_peripheral                )  //i
  );
  UsbLsFsPhyFilter ports_1_filter (
    .io_lowSpeed       (io_ctrl_lowSpeed                ), //i
    .io_usb_dp         (io_usb_1_rx_dp                  ), //i
    .io_usb_dm         (io_usb_1_rx_dm                  ), //i
    .io_filtred_dp     (ports_1_filter_io_filtred_dp    ), //o
    .io_filtred_dm     (ports_1_filter_io_filtred_dm    ), //o
    .io_filtred_d      (ports_1_filter_io_filtred_d     ), //o
    .io_filtred_se0    (ports_1_filter_io_filtred_se0   ), //o
    .io_filtred_sample (ports_1_filter_io_filtred_sample), //o
    .clk_peripheral    (clk_peripheral                  ), //i
    .reset_peripheral  (reset_peripheral                )  //i
  );
  `ifndef SYNTHESIS
  always @(*) begin
    case(txShared_frame_stateReg)
      txShared_frame_enumDef_BOOT : txShared_frame_stateReg_string = "BOOT          ";
      txShared_frame_enumDef_IDLE : txShared_frame_stateReg_string = "IDLE          ";
      txShared_frame_enumDef_TAKE_LINE : txShared_frame_stateReg_string = "TAKE_LINE     ";
      txShared_frame_enumDef_PREAMBLE_SYNC : txShared_frame_stateReg_string = "PREAMBLE_SYNC ";
      txShared_frame_enumDef_PREAMBLE_PID : txShared_frame_stateReg_string = "PREAMBLE_PID  ";
      txShared_frame_enumDef_PREAMBLE_DELAY : txShared_frame_stateReg_string = "PREAMBLE_DELAY";
      txShared_frame_enumDef_SYNC : txShared_frame_stateReg_string = "SYNC          ";
      txShared_frame_enumDef_DATA : txShared_frame_stateReg_string = "DATA          ";
      txShared_frame_enumDef_EOP_0 : txShared_frame_stateReg_string = "EOP_0         ";
      txShared_frame_enumDef_EOP_1 : txShared_frame_stateReg_string = "EOP_1         ";
      txShared_frame_enumDef_EOP_2 : txShared_frame_stateReg_string = "EOP_2         ";
      default : txShared_frame_stateReg_string = "??????????????";
    endcase
  end
  always @(*) begin
    case(txShared_frame_stateNext)
      txShared_frame_enumDef_BOOT : txShared_frame_stateNext_string = "BOOT          ";
      txShared_frame_enumDef_IDLE : txShared_frame_stateNext_string = "IDLE          ";
      txShared_frame_enumDef_TAKE_LINE : txShared_frame_stateNext_string = "TAKE_LINE     ";
      txShared_frame_enumDef_PREAMBLE_SYNC : txShared_frame_stateNext_string = "PREAMBLE_SYNC ";
      txShared_frame_enumDef_PREAMBLE_PID : txShared_frame_stateNext_string = "PREAMBLE_PID  ";
      txShared_frame_enumDef_PREAMBLE_DELAY : txShared_frame_stateNext_string = "PREAMBLE_DELAY";
      txShared_frame_enumDef_SYNC : txShared_frame_stateNext_string = "SYNC          ";
      txShared_frame_enumDef_DATA : txShared_frame_stateNext_string = "DATA          ";
      txShared_frame_enumDef_EOP_0 : txShared_frame_stateNext_string = "EOP_0         ";
      txShared_frame_enumDef_EOP_1 : txShared_frame_stateNext_string = "EOP_1         ";
      txShared_frame_enumDef_EOP_2 : txShared_frame_stateNext_string = "EOP_2         ";
      default : txShared_frame_stateNext_string = "??????????????";
    endcase
  end
  always @(*) begin
    case(upstreamRx_stateReg)
      upstreamRx_enumDef_BOOT : upstreamRx_stateReg_string = "BOOT   ";
      upstreamRx_enumDef_IDLE : upstreamRx_stateReg_string = "IDLE   ";
      upstreamRx_enumDef_SUSPEND : upstreamRx_stateReg_string = "SUSPEND";
      default : upstreamRx_stateReg_string = "???????";
    endcase
  end
  always @(*) begin
    case(upstreamRx_stateNext)
      upstreamRx_enumDef_BOOT : upstreamRx_stateNext_string = "BOOT   ";
      upstreamRx_enumDef_IDLE : upstreamRx_stateNext_string = "IDLE   ";
      upstreamRx_enumDef_SUSPEND : upstreamRx_stateNext_string = "SUSPEND";
      default : upstreamRx_stateNext_string = "???????";
    endcase
  end
  always @(*) begin
    case(ports_0_rx_packet_stateReg)
      ports_0_rx_packet_enumDef_BOOT : ports_0_rx_packet_stateReg_string = "BOOT   ";
      ports_0_rx_packet_enumDef_IDLE : ports_0_rx_packet_stateReg_string = "IDLE   ";
      ports_0_rx_packet_enumDef_PACKET : ports_0_rx_packet_stateReg_string = "PACKET ";
      ports_0_rx_packet_enumDef_ERRORED : ports_0_rx_packet_stateReg_string = "ERRORED";
      default : ports_0_rx_packet_stateReg_string = "???????";
    endcase
  end
  always @(*) begin
    case(ports_0_rx_packet_stateNext)
      ports_0_rx_packet_enumDef_BOOT : ports_0_rx_packet_stateNext_string = "BOOT   ";
      ports_0_rx_packet_enumDef_IDLE : ports_0_rx_packet_stateNext_string = "IDLE   ";
      ports_0_rx_packet_enumDef_PACKET : ports_0_rx_packet_stateNext_string = "PACKET ";
      ports_0_rx_packet_enumDef_ERRORED : ports_0_rx_packet_stateNext_string = "ERRORED";
      default : ports_0_rx_packet_stateNext_string = "???????";
    endcase
  end
  always @(*) begin
    case(ports_0_fsm_stateReg)
      ports_0_fsm_enumDef_BOOT : ports_0_fsm_stateReg_string = "BOOT           ";
      ports_0_fsm_enumDef_POWER_OFF : ports_0_fsm_stateReg_string = "POWER_OFF      ";
      ports_0_fsm_enumDef_DISCONNECTED : ports_0_fsm_stateReg_string = "DISCONNECTED   ";
      ports_0_fsm_enumDef_DISABLED : ports_0_fsm_stateReg_string = "DISABLED       ";
      ports_0_fsm_enumDef_RESETTING : ports_0_fsm_stateReg_string = "RESETTING      ";
      ports_0_fsm_enumDef_RESETTING_DELAY : ports_0_fsm_stateReg_string = "RESETTING_DELAY";
      ports_0_fsm_enumDef_RESETTING_SYNC : ports_0_fsm_stateReg_string = "RESETTING_SYNC ";
      ports_0_fsm_enumDef_ENABLED : ports_0_fsm_stateReg_string = "ENABLED        ";
      ports_0_fsm_enumDef_SUSPENDED : ports_0_fsm_stateReg_string = "SUSPENDED      ";
      ports_0_fsm_enumDef_RESUMING : ports_0_fsm_stateReg_string = "RESUMING       ";
      ports_0_fsm_enumDef_SEND_EOP_0 : ports_0_fsm_stateReg_string = "SEND_EOP_0     ";
      ports_0_fsm_enumDef_SEND_EOP_1 : ports_0_fsm_stateReg_string = "SEND_EOP_1     ";
      ports_0_fsm_enumDef_RESTART_S : ports_0_fsm_stateReg_string = "RESTART_S      ";
      ports_0_fsm_enumDef_RESTART_E : ports_0_fsm_stateReg_string = "RESTART_E      ";
      default : ports_0_fsm_stateReg_string = "???????????????";
    endcase
  end
  always @(*) begin
    case(ports_0_fsm_stateNext)
      ports_0_fsm_enumDef_BOOT : ports_0_fsm_stateNext_string = "BOOT           ";
      ports_0_fsm_enumDef_POWER_OFF : ports_0_fsm_stateNext_string = "POWER_OFF      ";
      ports_0_fsm_enumDef_DISCONNECTED : ports_0_fsm_stateNext_string = "DISCONNECTED   ";
      ports_0_fsm_enumDef_DISABLED : ports_0_fsm_stateNext_string = "DISABLED       ";
      ports_0_fsm_enumDef_RESETTING : ports_0_fsm_stateNext_string = "RESETTING      ";
      ports_0_fsm_enumDef_RESETTING_DELAY : ports_0_fsm_stateNext_string = "RESETTING_DELAY";
      ports_0_fsm_enumDef_RESETTING_SYNC : ports_0_fsm_stateNext_string = "RESETTING_SYNC ";
      ports_0_fsm_enumDef_ENABLED : ports_0_fsm_stateNext_string = "ENABLED        ";
      ports_0_fsm_enumDef_SUSPENDED : ports_0_fsm_stateNext_string = "SUSPENDED      ";
      ports_0_fsm_enumDef_RESUMING : ports_0_fsm_stateNext_string = "RESUMING       ";
      ports_0_fsm_enumDef_SEND_EOP_0 : ports_0_fsm_stateNext_string = "SEND_EOP_0     ";
      ports_0_fsm_enumDef_SEND_EOP_1 : ports_0_fsm_stateNext_string = "SEND_EOP_1     ";
      ports_0_fsm_enumDef_RESTART_S : ports_0_fsm_stateNext_string = "RESTART_S      ";
      ports_0_fsm_enumDef_RESTART_E : ports_0_fsm_stateNext_string = "RESTART_E      ";
      default : ports_0_fsm_stateNext_string = "???????????????";
    endcase
  end
  always @(*) begin
    case(ports_1_rx_packet_stateReg)
      ports_1_rx_packet_enumDef_BOOT : ports_1_rx_packet_stateReg_string = "BOOT   ";
      ports_1_rx_packet_enumDef_IDLE : ports_1_rx_packet_stateReg_string = "IDLE   ";
      ports_1_rx_packet_enumDef_PACKET : ports_1_rx_packet_stateReg_string = "PACKET ";
      ports_1_rx_packet_enumDef_ERRORED : ports_1_rx_packet_stateReg_string = "ERRORED";
      default : ports_1_rx_packet_stateReg_string = "???????";
    endcase
  end
  always @(*) begin
    case(ports_1_rx_packet_stateNext)
      ports_1_rx_packet_enumDef_BOOT : ports_1_rx_packet_stateNext_string = "BOOT   ";
      ports_1_rx_packet_enumDef_IDLE : ports_1_rx_packet_stateNext_string = "IDLE   ";
      ports_1_rx_packet_enumDef_PACKET : ports_1_rx_packet_stateNext_string = "PACKET ";
      ports_1_rx_packet_enumDef_ERRORED : ports_1_rx_packet_stateNext_string = "ERRORED";
      default : ports_1_rx_packet_stateNext_string = "???????";
    endcase
  end
  always @(*) begin
    case(ports_1_fsm_stateReg)
      ports_1_fsm_enumDef_BOOT : ports_1_fsm_stateReg_string = "BOOT           ";
      ports_1_fsm_enumDef_POWER_OFF : ports_1_fsm_stateReg_string = "POWER_OFF      ";
      ports_1_fsm_enumDef_DISCONNECTED : ports_1_fsm_stateReg_string = "DISCONNECTED   ";
      ports_1_fsm_enumDef_DISABLED : ports_1_fsm_stateReg_string = "DISABLED       ";
      ports_1_fsm_enumDef_RESETTING : ports_1_fsm_stateReg_string = "RESETTING      ";
      ports_1_fsm_enumDef_RESETTING_DELAY : ports_1_fsm_stateReg_string = "RESETTING_DELAY";
      ports_1_fsm_enumDef_RESETTING_SYNC : ports_1_fsm_stateReg_string = "RESETTING_SYNC ";
      ports_1_fsm_enumDef_ENABLED : ports_1_fsm_stateReg_string = "ENABLED        ";
      ports_1_fsm_enumDef_SUSPENDED : ports_1_fsm_stateReg_string = "SUSPENDED      ";
      ports_1_fsm_enumDef_RESUMING : ports_1_fsm_stateReg_string = "RESUMING       ";
      ports_1_fsm_enumDef_SEND_EOP_0 : ports_1_fsm_stateReg_string = "SEND_EOP_0     ";
      ports_1_fsm_enumDef_SEND_EOP_1 : ports_1_fsm_stateReg_string = "SEND_EOP_1     ";
      ports_1_fsm_enumDef_RESTART_S : ports_1_fsm_stateReg_string = "RESTART_S      ";
      ports_1_fsm_enumDef_RESTART_E : ports_1_fsm_stateReg_string = "RESTART_E      ";
      default : ports_1_fsm_stateReg_string = "???????????????";
    endcase
  end
  always @(*) begin
    case(ports_1_fsm_stateNext)
      ports_1_fsm_enumDef_BOOT : ports_1_fsm_stateNext_string = "BOOT           ";
      ports_1_fsm_enumDef_POWER_OFF : ports_1_fsm_stateNext_string = "POWER_OFF      ";
      ports_1_fsm_enumDef_DISCONNECTED : ports_1_fsm_stateNext_string = "DISCONNECTED   ";
      ports_1_fsm_enumDef_DISABLED : ports_1_fsm_stateNext_string = "DISABLED       ";
      ports_1_fsm_enumDef_RESETTING : ports_1_fsm_stateNext_string = "RESETTING      ";
      ports_1_fsm_enumDef_RESETTING_DELAY : ports_1_fsm_stateNext_string = "RESETTING_DELAY";
      ports_1_fsm_enumDef_RESETTING_SYNC : ports_1_fsm_stateNext_string = "RESETTING_SYNC ";
      ports_1_fsm_enumDef_ENABLED : ports_1_fsm_stateNext_string = "ENABLED        ";
      ports_1_fsm_enumDef_SUSPENDED : ports_1_fsm_stateNext_string = "SUSPENDED      ";
      ports_1_fsm_enumDef_RESUMING : ports_1_fsm_stateNext_string = "RESUMING       ";
      ports_1_fsm_enumDef_SEND_EOP_0 : ports_1_fsm_stateNext_string = "SEND_EOP_0     ";
      ports_1_fsm_enumDef_SEND_EOP_1 : ports_1_fsm_stateNext_string = "SEND_EOP_1     ";
      ports_1_fsm_enumDef_RESTART_S : ports_1_fsm_stateNext_string = "RESTART_S      ";
      ports_1_fsm_enumDef_RESTART_E : ports_1_fsm_stateNext_string = "RESTART_E      ";
      default : ports_1_fsm_stateNext_string = "???????????????";
    endcase
  end
  `endif

  assign tickTimer_counter_willClear = 1'b0;
  assign tickTimer_counter_willOverflowIfInc = (tickTimer_counter_value == 2'b11);
  assign tickTimer_counter_willOverflow = (tickTimer_counter_willOverflowIfInc && tickTimer_counter_willIncrement);
  always @(*) begin
    tickTimer_counter_valueNext = (tickTimer_counter_value + _zz_tickTimer_counter_valueNext);
    if(tickTimer_counter_willClear) begin
      tickTimer_counter_valueNext = 2'b00;
    end
  end

  assign tickTimer_counter_willIncrement = 1'b1;
  assign tickTimer_tick = (tickTimer_counter_willOverflow == 1'b1);
  assign io_ctrl_tick = tickTimer_tick;
  always @(*) begin
    txShared_timer_clear = 1'b0;
    if(txShared_encoder_input_valid) begin
      if(txShared_encoder_input_data) begin
        if(txShared_timer_oneCycle) begin
          if(when_usbphy_l91) begin
            txShared_timer_clear = 1'b1;
          end
        end
      end
    end
    if(txShared_encoder_input_ready) begin
      txShared_timer_clear = 1'b1;
    end
    case(txShared_frame_stateReg)
      txShared_frame_enumDef_IDLE : begin
        txShared_timer_clear = 1'b1;
      end
      txShared_frame_enumDef_TAKE_LINE : begin
        if(txShared_timer_oneCycle) begin
          txShared_timer_clear = 1'b1;
        end
      end
      txShared_frame_enumDef_PREAMBLE_SYNC : begin
      end
      txShared_frame_enumDef_PREAMBLE_PID : begin
      end
      txShared_frame_enumDef_PREAMBLE_DELAY : begin
        if(txShared_timer_fourCycle) begin
          txShared_timer_clear = 1'b1;
        end
      end
      txShared_frame_enumDef_SYNC : begin
      end
      txShared_frame_enumDef_DATA : begin
      end
      txShared_frame_enumDef_EOP_0 : begin
        if(txShared_timer_twoCycle) begin
          txShared_timer_clear = 1'b1;
        end
      end
      txShared_frame_enumDef_EOP_1 : begin
        if(txShared_timer_oneCycle) begin
          txShared_timer_clear = 1'b1;
        end
      end
      txShared_frame_enumDef_EOP_2 : begin
        if(txShared_timer_twoCycle) begin
          txShared_timer_clear = 1'b1;
        end
      end
      default : begin
      end
    endcase
  end

  assign txShared_timer_inc = 1'b1;
  assign txShared_timer_oneCycle = (txShared_timer_counter == _zz_txShared_timer_oneCycle);
  assign txShared_timer_twoCycle = (txShared_timer_counter == _zz_txShared_timer_twoCycle);
  assign txShared_timer_fourCycle = (txShared_timer_counter == _zz_txShared_timer_fourCycle);
  always @(*) begin
    txShared_timer_lowSpeed = 1'b0;
    if(txShared_encoder_input_valid) begin
      txShared_timer_lowSpeed = txShared_encoder_input_lowSpeed;
    end
    case(txShared_frame_stateReg)
      txShared_frame_enumDef_IDLE : begin
      end
      txShared_frame_enumDef_TAKE_LINE : begin
        txShared_timer_lowSpeed = 1'b0;
      end
      txShared_frame_enumDef_PREAMBLE_SYNC : begin
      end
      txShared_frame_enumDef_PREAMBLE_PID : begin
      end
      txShared_frame_enumDef_PREAMBLE_DELAY : begin
        txShared_timer_lowSpeed = 1'b0;
      end
      txShared_frame_enumDef_SYNC : begin
      end
      txShared_frame_enumDef_DATA : begin
      end
      txShared_frame_enumDef_EOP_0 : begin
        txShared_timer_lowSpeed = txShared_frame_wasLowSpeed;
      end
      txShared_frame_enumDef_EOP_1 : begin
        txShared_timer_lowSpeed = txShared_frame_wasLowSpeed;
      end
      txShared_frame_enumDef_EOP_2 : begin
        txShared_timer_lowSpeed = txShared_frame_wasLowSpeed;
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    txShared_rxToTxDelay_clear = 1'b0;
    if(ports_0_rx_eop_hit) begin
      txShared_rxToTxDelay_clear = 1'b1;
    end
    if(ports_1_rx_eop_hit) begin
      txShared_rxToTxDelay_clear = 1'b1;
    end
  end

  assign txShared_rxToTxDelay_inc = 1'b1;
  assign txShared_rxToTxDelay_twoCycle = (txShared_rxToTxDelay_counter == _zz_txShared_rxToTxDelay_twoCycle);
  always @(*) begin
    txShared_encoder_input_valid = 1'b0;
    if(txShared_serialiser_input_valid) begin
      txShared_encoder_input_valid = 1'b1;
    end
  end

  always @(*) begin
    txShared_encoder_input_ready = 1'b0;
    if(txShared_encoder_input_valid) begin
      if(txShared_encoder_input_data) begin
        if(txShared_timer_oneCycle) begin
          txShared_encoder_input_ready = 1'b1;
          if(when_usbphy_l91) begin
            txShared_encoder_input_ready = 1'b0;
          end
        end
      end else begin
        if(txShared_timer_oneCycle) begin
          txShared_encoder_input_ready = 1'b1;
        end
      end
    end
  end

  always @(*) begin
    txShared_encoder_input_data = 1'bx;
    if(txShared_serialiser_input_valid) begin
      txShared_encoder_input_data = txShared_serialiser_input_data[txShared_serialiser_bitCounter];
    end
  end

  always @(*) begin
    txShared_encoder_input_lowSpeed = 1'bx;
    if(txShared_serialiser_input_valid) begin
      txShared_encoder_input_lowSpeed = txShared_serialiser_input_lowSpeed;
    end
  end

  always @(*) begin
    txShared_encoder_output_valid = 1'b0;
    if(txShared_encoder_input_valid) begin
      txShared_encoder_output_valid = txShared_encoder_input_valid;
    end
    case(txShared_frame_stateReg)
      txShared_frame_enumDef_IDLE : begin
      end
      txShared_frame_enumDef_TAKE_LINE : begin
        txShared_encoder_output_valid = 1'b1;
      end
      txShared_frame_enumDef_PREAMBLE_SYNC : begin
      end
      txShared_frame_enumDef_PREAMBLE_PID : begin
      end
      txShared_frame_enumDef_PREAMBLE_DELAY : begin
        txShared_encoder_output_valid = 1'b1;
      end
      txShared_frame_enumDef_SYNC : begin
      end
      txShared_frame_enumDef_DATA : begin
      end
      txShared_frame_enumDef_EOP_0 : begin
        txShared_encoder_output_valid = 1'b1;
      end
      txShared_frame_enumDef_EOP_1 : begin
        txShared_encoder_output_valid = 1'b1;
      end
      txShared_frame_enumDef_EOP_2 : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    txShared_encoder_output_se0 = 1'b0;
    case(txShared_frame_stateReg)
      txShared_frame_enumDef_IDLE : begin
      end
      txShared_frame_enumDef_TAKE_LINE : begin
      end
      txShared_frame_enumDef_PREAMBLE_SYNC : begin
      end
      txShared_frame_enumDef_PREAMBLE_PID : begin
      end
      txShared_frame_enumDef_PREAMBLE_DELAY : begin
      end
      txShared_frame_enumDef_SYNC : begin
      end
      txShared_frame_enumDef_DATA : begin
      end
      txShared_frame_enumDef_EOP_0 : begin
        txShared_encoder_output_se0 = 1'b1;
      end
      txShared_frame_enumDef_EOP_1 : begin
      end
      txShared_frame_enumDef_EOP_2 : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    txShared_encoder_output_lowSpeed = 1'bx;
    if(txShared_encoder_input_valid) begin
      txShared_encoder_output_lowSpeed = txShared_encoder_input_lowSpeed;
    end
    case(txShared_frame_stateReg)
      txShared_frame_enumDef_IDLE : begin
      end
      txShared_frame_enumDef_TAKE_LINE : begin
        txShared_encoder_output_lowSpeed = 1'b0;
      end
      txShared_frame_enumDef_PREAMBLE_SYNC : begin
      end
      txShared_frame_enumDef_PREAMBLE_PID : begin
      end
      txShared_frame_enumDef_PREAMBLE_DELAY : begin
        txShared_encoder_output_lowSpeed = 1'b0;
      end
      txShared_frame_enumDef_SYNC : begin
      end
      txShared_frame_enumDef_DATA : begin
      end
      txShared_frame_enumDef_EOP_0 : begin
        txShared_encoder_output_lowSpeed = txShared_frame_wasLowSpeed;
      end
      txShared_frame_enumDef_EOP_1 : begin
        txShared_encoder_output_lowSpeed = txShared_frame_wasLowSpeed;
      end
      txShared_frame_enumDef_EOP_2 : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    txShared_encoder_output_data = 1'bx;
    if(txShared_encoder_input_valid) begin
      if(txShared_encoder_input_data) begin
        txShared_encoder_output_data = txShared_encoder_state;
      end else begin
        txShared_encoder_output_data = (! txShared_encoder_state);
      end
    end
    case(txShared_frame_stateReg)
      txShared_frame_enumDef_IDLE : begin
      end
      txShared_frame_enumDef_TAKE_LINE : begin
        txShared_encoder_output_data = 1'b1;
      end
      txShared_frame_enumDef_PREAMBLE_SYNC : begin
      end
      txShared_frame_enumDef_PREAMBLE_PID : begin
      end
      txShared_frame_enumDef_PREAMBLE_DELAY : begin
        txShared_encoder_output_data = 1'b1;
      end
      txShared_frame_enumDef_SYNC : begin
      end
      txShared_frame_enumDef_DATA : begin
      end
      txShared_frame_enumDef_EOP_0 : begin
      end
      txShared_frame_enumDef_EOP_1 : begin
        txShared_encoder_output_data = 1'b1;
      end
      txShared_frame_enumDef_EOP_2 : begin
      end
      default : begin
      end
    endcase
  end

  assign when_usbphy_l91 = (txShared_encoder_counter == 3'b101);
  assign when_usbphy_l96 = (txShared_encoder_counter == 3'b110);
  assign when_usbphy_l110 = (! txShared_encoder_input_valid);
  always @(*) begin
    txShared_serialiser_input_valid = 1'b0;
    case(txShared_frame_stateReg)
      txShared_frame_enumDef_IDLE : begin
      end
      txShared_frame_enumDef_TAKE_LINE : begin
      end
      txShared_frame_enumDef_PREAMBLE_SYNC : begin
        txShared_serialiser_input_valid = 1'b1;
      end
      txShared_frame_enumDef_PREAMBLE_PID : begin
        txShared_serialiser_input_valid = 1'b1;
      end
      txShared_frame_enumDef_PREAMBLE_DELAY : begin
      end
      txShared_frame_enumDef_SYNC : begin
        txShared_serialiser_input_valid = 1'b1;
      end
      txShared_frame_enumDef_DATA : begin
        txShared_serialiser_input_valid = 1'b1;
      end
      txShared_frame_enumDef_EOP_0 : begin
      end
      txShared_frame_enumDef_EOP_1 : begin
      end
      txShared_frame_enumDef_EOP_2 : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    txShared_serialiser_input_ready = 1'b0;
    if(txShared_serialiser_input_valid) begin
      if(txShared_encoder_input_ready) begin
        if(when_usbphy_l136) begin
          txShared_serialiser_input_ready = 1'b1;
        end
      end
    end
  end

  always @(*) begin
    txShared_serialiser_input_data = 8'bxxxxxxxx;
    case(txShared_frame_stateReg)
      txShared_frame_enumDef_IDLE : begin
      end
      txShared_frame_enumDef_TAKE_LINE : begin
      end
      txShared_frame_enumDef_PREAMBLE_SYNC : begin
        txShared_serialiser_input_data = 8'h80;
      end
      txShared_frame_enumDef_PREAMBLE_PID : begin
        txShared_serialiser_input_data = 8'h3c;
      end
      txShared_frame_enumDef_PREAMBLE_DELAY : begin
      end
      txShared_frame_enumDef_SYNC : begin
        txShared_serialiser_input_data = 8'h80;
      end
      txShared_frame_enumDef_DATA : begin
        txShared_serialiser_input_data = io_ctrl_tx_payload_fragment;
      end
      txShared_frame_enumDef_EOP_0 : begin
      end
      txShared_frame_enumDef_EOP_1 : begin
      end
      txShared_frame_enumDef_EOP_2 : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    txShared_serialiser_input_lowSpeed = 1'bx;
    case(txShared_frame_stateReg)
      txShared_frame_enumDef_IDLE : begin
      end
      txShared_frame_enumDef_TAKE_LINE : begin
      end
      txShared_frame_enumDef_PREAMBLE_SYNC : begin
        txShared_serialiser_input_lowSpeed = 1'b0;
      end
      txShared_frame_enumDef_PREAMBLE_PID : begin
        txShared_serialiser_input_lowSpeed = 1'b0;
      end
      txShared_frame_enumDef_PREAMBLE_DELAY : begin
      end
      txShared_frame_enumDef_SYNC : begin
        txShared_serialiser_input_lowSpeed = txShared_frame_wasLowSpeed;
      end
      txShared_frame_enumDef_DATA : begin
        txShared_serialiser_input_lowSpeed = txShared_frame_wasLowSpeed;
      end
      txShared_frame_enumDef_EOP_0 : begin
      end
      txShared_frame_enumDef_EOP_1 : begin
      end
      txShared_frame_enumDef_EOP_2 : begin
      end
      default : begin
      end
    endcase
  end

  assign when_usbphy_l136 = (txShared_serialiser_bitCounter == 3'b111);
  assign when_usbphy_l142 = ((! txShared_serialiser_input_valid) || txShared_serialiser_input_ready);
  always @(*) begin
    txShared_lowSpeedSof_increment = 1'b0;
    if(when_usbphy_l153) begin
      if(when_usbphy_l154) begin
        txShared_lowSpeedSof_increment = 1'b1;
      end
    end
  end

  assign when_usbphy_l151 = ((! txShared_encoder_output_valid) && txShared_encoder_output_valid_regNext);
  assign when_usbphy_l153 = (txShared_lowSpeedSof_state == 2'b00);
  assign io_ctrl_tx_fire = (io_ctrl_tx_valid && io_ctrl_tx_ready);
  assign when_usbphy_l154 = ((io_ctrl_tx_valid && io_ctrl_tx_payload_first) && (io_ctrl_tx_payload_fragment == 8'ha5));
  assign when_usbphy_l161 = (txShared_lowSpeedSof_timer == 5'h1f);
  assign txShared_lowSpeedSof_valid = (txShared_lowSpeedSof_state != 2'b00);
  assign txShared_lowSpeedSof_data = 1'b0;
  assign txShared_lowSpeedSof_se0 = (txShared_lowSpeedSof_state != 2'b11);
  assign txShared_frame_wantExit = 1'b0;
  always @(*) begin
    txShared_frame_wantStart = 1'b0;
    case(txShared_frame_stateReg)
      txShared_frame_enumDef_IDLE : begin
      end
      txShared_frame_enumDef_TAKE_LINE : begin
      end
      txShared_frame_enumDef_PREAMBLE_SYNC : begin
      end
      txShared_frame_enumDef_PREAMBLE_PID : begin
      end
      txShared_frame_enumDef_PREAMBLE_DELAY : begin
      end
      txShared_frame_enumDef_SYNC : begin
      end
      txShared_frame_enumDef_DATA : begin
      end
      txShared_frame_enumDef_EOP_0 : begin
      end
      txShared_frame_enumDef_EOP_1 : begin
      end
      txShared_frame_enumDef_EOP_2 : begin
      end
      default : begin
        txShared_frame_wantStart = 1'b1;
      end
    endcase
  end

  assign txShared_frame_wantKill = 1'b0;
  assign txShared_frame_busy = (! (txShared_frame_stateReg == txShared_frame_enumDef_BOOT));
  always @(*) begin
    io_ctrl_tx_ready = 1'b0;
    case(txShared_frame_stateReg)
      txShared_frame_enumDef_IDLE : begin
      end
      txShared_frame_enumDef_TAKE_LINE : begin
      end
      txShared_frame_enumDef_PREAMBLE_SYNC : begin
      end
      txShared_frame_enumDef_PREAMBLE_PID : begin
      end
      txShared_frame_enumDef_PREAMBLE_DELAY : begin
      end
      txShared_frame_enumDef_SYNC : begin
      end
      txShared_frame_enumDef_DATA : begin
        if(txShared_serialiser_input_ready) begin
          io_ctrl_tx_ready = 1'b1;
        end
      end
      txShared_frame_enumDef_EOP_0 : begin
      end
      txShared_frame_enumDef_EOP_1 : begin
      end
      txShared_frame_enumDef_EOP_2 : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    io_ctrl_txEop = 1'b0;
    case(txShared_frame_stateReg)
      txShared_frame_enumDef_IDLE : begin
      end
      txShared_frame_enumDef_TAKE_LINE : begin
      end
      txShared_frame_enumDef_PREAMBLE_SYNC : begin
      end
      txShared_frame_enumDef_PREAMBLE_PID : begin
      end
      txShared_frame_enumDef_PREAMBLE_DELAY : begin
      end
      txShared_frame_enumDef_SYNC : begin
      end
      txShared_frame_enumDef_DATA : begin
      end
      txShared_frame_enumDef_EOP_0 : begin
        if(txShared_timer_twoCycle) begin
          io_ctrl_txEop = 1'b1;
        end
      end
      txShared_frame_enumDef_EOP_1 : begin
      end
      txShared_frame_enumDef_EOP_2 : begin
      end
      default : begin
      end
    endcase
  end

  assign upstreamRx_wantExit = 1'b0;
  always @(*) begin
    upstreamRx_wantStart = 1'b0;
    case(upstreamRx_stateReg)
      upstreamRx_enumDef_IDLE : begin
      end
      upstreamRx_enumDef_SUSPEND : begin
      end
      default : begin
        upstreamRx_wantStart = 1'b1;
      end
    endcase
  end

  assign upstreamRx_wantKill = 1'b0;
  always @(*) begin
    upstreamRx_timer_clear = 1'b0;
    if(txShared_encoder_output_valid) begin
      upstreamRx_timer_clear = 1'b1;
    end
  end

  assign upstreamRx_timer_inc = 1'b1;
  assign upstreamRx_timer_IDLE_EOI = (upstreamRx_timer_counter == 20'h2327f);
  assign io_ctrl_overcurrent = 1'b0;
  always @(*) begin
    io_ctrl_rx_flow_valid = 1'b0;
    case(ports_0_rx_packet_stateReg)
      ports_0_rx_packet_enumDef_IDLE : begin
      end
      ports_0_rx_packet_enumDef_PACKET : begin
        if(ports_0_rx_destuffer_output_valid) begin
          if(when_usbphy_l429) begin
            io_ctrl_rx_flow_valid = ports_0_rx_enablePackets;
          end
        end
      end
      ports_0_rx_packet_enumDef_ERRORED : begin
      end
      default : begin
      end
    endcase
    case(ports_1_rx_packet_stateReg)
      ports_1_rx_packet_enumDef_IDLE : begin
      end
      ports_1_rx_packet_enumDef_PACKET : begin
        if(ports_1_rx_destuffer_output_valid) begin
          if(when_usbphy_l429_1) begin
            io_ctrl_rx_flow_valid = ports_1_rx_enablePackets;
          end
        end
      end
      ports_1_rx_packet_enumDef_ERRORED : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    io_ctrl_rx_active = 1'b0;
    case(ports_0_rx_packet_stateReg)
      ports_0_rx_packet_enumDef_IDLE : begin
      end
      ports_0_rx_packet_enumDef_PACKET : begin
        io_ctrl_rx_active = 1'b1;
      end
      ports_0_rx_packet_enumDef_ERRORED : begin
        io_ctrl_rx_active = 1'b1;
      end
      default : begin
      end
    endcase
    case(ports_1_rx_packet_stateReg)
      ports_1_rx_packet_enumDef_IDLE : begin
      end
      ports_1_rx_packet_enumDef_PACKET : begin
        io_ctrl_rx_active = 1'b1;
      end
      ports_1_rx_packet_enumDef_ERRORED : begin
        io_ctrl_rx_active = 1'b1;
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    io_ctrl_rx_flow_payload_stuffingError = 1'b0;
    case(ports_0_rx_packet_stateReg)
      ports_0_rx_packet_enumDef_IDLE : begin
      end
      ports_0_rx_packet_enumDef_PACKET : begin
        io_ctrl_rx_flow_payload_stuffingError = ports_0_rx_stuffingError;
      end
      ports_0_rx_packet_enumDef_ERRORED : begin
      end
      default : begin
      end
    endcase
    case(ports_1_rx_packet_stateReg)
      ports_1_rx_packet_enumDef_IDLE : begin
      end
      ports_1_rx_packet_enumDef_PACKET : begin
        io_ctrl_rx_flow_payload_stuffingError = ports_1_rx_stuffingError;
      end
      ports_1_rx_packet_enumDef_ERRORED : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    io_ctrl_rx_flow_payload_data = 8'bxxxxxxxx;
    case(ports_0_rx_packet_stateReg)
      ports_0_rx_packet_enumDef_IDLE : begin
      end
      ports_0_rx_packet_enumDef_PACKET : begin
        io_ctrl_rx_flow_payload_data = ports_0_rx_history_value;
      end
      ports_0_rx_packet_enumDef_ERRORED : begin
      end
      default : begin
      end
    endcase
    case(ports_1_rx_packet_stateReg)
      ports_1_rx_packet_enumDef_IDLE : begin
      end
      ports_1_rx_packet_enumDef_PACKET : begin
        io_ctrl_rx_flow_payload_data = ports_1_rx_history_value;
      end
      ports_1_rx_packet_enumDef_ERRORED : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    resumeFromPort = 1'b0;
    case(ports_0_fsm_stateReg)
      ports_0_fsm_enumDef_POWER_OFF : begin
      end
      ports_0_fsm_enumDef_DISCONNECTED : begin
      end
      ports_0_fsm_enumDef_DISABLED : begin
      end
      ports_0_fsm_enumDef_RESETTING : begin
      end
      ports_0_fsm_enumDef_RESETTING_DELAY : begin
      end
      ports_0_fsm_enumDef_RESETTING_SYNC : begin
      end
      ports_0_fsm_enumDef_ENABLED : begin
      end
      ports_0_fsm_enumDef_SUSPENDED : begin
      end
      ports_0_fsm_enumDef_RESUMING : begin
      end
      ports_0_fsm_enumDef_SEND_EOP_0 : begin
      end
      ports_0_fsm_enumDef_SEND_EOP_1 : begin
      end
      ports_0_fsm_enumDef_RESTART_S : begin
        if(when_usbphy_l653) begin
          resumeFromPort = 1'b1;
        end
      end
      ports_0_fsm_enumDef_RESTART_E : begin
        if(when_usbphy_l663) begin
          resumeFromPort = 1'b1;
        end
      end
      default : begin
      end
    endcase
    case(ports_1_fsm_stateReg)
      ports_1_fsm_enumDef_POWER_OFF : begin
      end
      ports_1_fsm_enumDef_DISCONNECTED : begin
      end
      ports_1_fsm_enumDef_DISABLED : begin
      end
      ports_1_fsm_enumDef_RESETTING : begin
      end
      ports_1_fsm_enumDef_RESETTING_DELAY : begin
      end
      ports_1_fsm_enumDef_RESETTING_SYNC : begin
      end
      ports_1_fsm_enumDef_ENABLED : begin
      end
      ports_1_fsm_enumDef_SUSPENDED : begin
      end
      ports_1_fsm_enumDef_RESUMING : begin
      end
      ports_1_fsm_enumDef_SEND_EOP_0 : begin
      end
      ports_1_fsm_enumDef_SEND_EOP_1 : begin
      end
      ports_1_fsm_enumDef_RESTART_S : begin
        if(when_usbphy_l653_1) begin
          resumeFromPort = 1'b1;
        end
      end
      ports_1_fsm_enumDef_RESTART_E : begin
        if(when_usbphy_l663_1) begin
          resumeFromPort = 1'b1;
        end
      end
      default : begin
      end
    endcase
  end

  assign io_ctrl_ports_0_lowSpeed = ports_0_portLowSpeed;
  assign io_ctrl_ports_0_remoteResume = 1'b0;
  always @(*) begin
    ports_0_rx_enablePackets = 1'b0;
    case(ports_0_fsm_stateReg)
      ports_0_fsm_enumDef_POWER_OFF : begin
      end
      ports_0_fsm_enumDef_DISCONNECTED : begin
      end
      ports_0_fsm_enumDef_DISABLED : begin
      end
      ports_0_fsm_enumDef_RESETTING : begin
      end
      ports_0_fsm_enumDef_RESETTING_DELAY : begin
      end
      ports_0_fsm_enumDef_RESETTING_SYNC : begin
      end
      ports_0_fsm_enumDef_ENABLED : begin
        ports_0_rx_enablePackets = 1'b1;
      end
      ports_0_fsm_enumDef_SUSPENDED : begin
      end
      ports_0_fsm_enumDef_RESUMING : begin
      end
      ports_0_fsm_enumDef_SEND_EOP_0 : begin
      end
      ports_0_fsm_enumDef_SEND_EOP_1 : begin
      end
      ports_0_fsm_enumDef_RESTART_S : begin
      end
      ports_0_fsm_enumDef_RESTART_E : begin
      end
      default : begin
      end
    endcase
  end

  assign ports_0_rx_j = ((ports_0_filter_io_filtred_dp == (! ports_0_portLowSpeed)) && (ports_0_filter_io_filtred_dm == ports_0_portLowSpeed));
  assign ports_0_rx_k = ((ports_0_filter_io_filtred_dp == ports_0_portLowSpeed) && (ports_0_filter_io_filtred_dm == (! ports_0_portLowSpeed)));
  assign io_management_0_power = io_ctrl_ports_0_power;
  assign io_ctrl_ports_0_overcurrent = io_management_0_overcurrent;
  always @(*) begin
    ports_0_rx_waitSync = 1'b0;
    case(ports_0_rx_packet_stateReg)
      ports_0_rx_packet_enumDef_IDLE : begin
        ports_0_rx_waitSync = 1'b1;
      end
      ports_0_rx_packet_enumDef_PACKET : begin
      end
      ports_0_rx_packet_enumDef_ERRORED : begin
      end
      default : begin
      end
    endcase
    if(when_StateMachine_l253) begin
      ports_0_rx_waitSync = 1'b1;
    end
  end

  always @(*) begin
    ports_0_rx_decoder_output_valid = 1'b0;
    if(ports_0_filter_io_filtred_sample) begin
      ports_0_rx_decoder_output_valid = 1'b1;
    end
  end

  always @(*) begin
    ports_0_rx_decoder_output_payload = 1'bx;
    if(ports_0_filter_io_filtred_sample) begin
      if(when_usbphy_l347) begin
        ports_0_rx_decoder_output_payload = 1'b0;
      end else begin
        ports_0_rx_decoder_output_payload = 1'b1;
      end
    end
  end

  assign when_usbphy_l347 = ((ports_0_rx_decoder_state ^ ports_0_filter_io_filtred_d) ^ ports_0_portLowSpeed);
  assign ports_0_rx_destuffer_unstuffNext = (ports_0_rx_destuffer_counter == 3'b110);
  assign ports_0_rx_destuffer_output_valid = (ports_0_rx_decoder_output_valid && (! ports_0_rx_destuffer_unstuffNext));
  assign ports_0_rx_destuffer_output_payload = ports_0_rx_decoder_output_payload;
  assign when_usbphy_l368 = ((! ports_0_rx_decoder_output_payload) || ports_0_rx_destuffer_unstuffNext);
  assign ports_0_rx_history_updated = ports_0_rx_destuffer_output_valid;
  assign _zz_ports_0_rx_history_value = ports_0_rx_destuffer_output_payload;
  assign ports_0_rx_history_value = {_zz_ports_0_rx_history_value,{_zz_ports_0_rx_history_value_1,{_zz_ports_0_rx_history_value_2,{_zz_ports_0_rx_history_value_3,{_zz_ports_0_rx_history_value_4,{_zz_ports_0_rx_history_value_5,{_zz_ports_0_rx_history_value_6,_zz_ports_0_rx_history_value_7}}}}}}};
  assign ports_0_rx_history_sync_hit = (ports_0_rx_history_updated && (ports_0_rx_history_value == 8'hd5));
  assign ports_0_rx_eop_maxThreshold = (io_ctrl_lowSpeed ? 7'h60 : 7'h0c);
  assign ports_0_rx_eop_minThreshold = (io_ctrl_lowSpeed ? 6'h2a : 6'h05);
  assign ports_0_rx_eop_maxHit = (ports_0_rx_eop_counter == ports_0_rx_eop_maxThreshold);
  always @(*) begin
    ports_0_rx_eop_hit = 1'b0;
    if(ports_0_rx_j) begin
      if(when_usbphy_l403) begin
        ports_0_rx_eop_hit = 1'b1;
      end
    end
  end

  assign when_usbphy_l395 = ((! ports_0_filter_io_filtred_dp) && (! ports_0_filter_io_filtred_dm));
  assign when_usbphy_l396 = (! ports_0_rx_eop_maxHit);
  assign when_usbphy_l403 = ((_zz_when_usbphy_l403 <= ports_0_rx_eop_counter) && (! ports_0_rx_eop_maxHit));
  assign ports_0_rx_packet_wantExit = 1'b0;
  always @(*) begin
    ports_0_rx_packet_wantStart = 1'b0;
    case(ports_0_rx_packet_stateReg)
      ports_0_rx_packet_enumDef_IDLE : begin
      end
      ports_0_rx_packet_enumDef_PACKET : begin
      end
      ports_0_rx_packet_enumDef_ERRORED : begin
      end
      default : begin
        ports_0_rx_packet_wantStart = 1'b1;
      end
    endcase
  end

  assign ports_0_rx_packet_wantKill = 1'b0;
  always @(*) begin
    ports_0_rx_packet_errorTimeout_clear = 1'b0;
    case(ports_0_rx_packet_stateReg)
      ports_0_rx_packet_enumDef_IDLE : begin
      end
      ports_0_rx_packet_enumDef_PACKET : begin
      end
      ports_0_rx_packet_enumDef_ERRORED : begin
        if(when_usbphy_l451) begin
          ports_0_rx_packet_errorTimeout_clear = 1'b1;
        end
      end
      default : begin
      end
    endcase
    if(when_StateMachine_l253_1) begin
      ports_0_rx_packet_errorTimeout_clear = 1'b1;
    end
  end

  assign ports_0_rx_packet_errorTimeout_inc = 1'b1;
  assign ports_0_rx_packet_errorTimeout_lowSpeed = io_ctrl_lowSpeed;
  assign ports_0_rx_packet_errorTimeout_trigger = (ports_0_rx_packet_errorTimeout_counter == _zz_ports_0_rx_packet_errorTimeout_trigger);
  always @(*) begin
    ports_0_rx_disconnect_clear = 1'b0;
    if(when_usbphy_l475) begin
      ports_0_rx_disconnect_clear = 1'b1;
    end
    if(when_usbphy_l672) begin
      ports_0_rx_disconnect_clear = 1'b1;
    end
  end

  assign ports_0_rx_disconnect_hit = (ports_0_rx_disconnect_counter == 7'h68);
  assign ports_0_rx_disconnect_event = (ports_0_rx_disconnect_hit && (! ports_0_rx_disconnect_hitLast));
  assign when_usbphy_l475 = ((! ports_0_filter_io_filtred_se0) || io_usb_0_tx_enable);
  assign io_ctrl_ports_0_disconnect = ports_0_rx_disconnect_event;
  assign ports_0_fsm_wantExit = 1'b0;
  always @(*) begin
    ports_0_fsm_wantStart = 1'b0;
    case(ports_0_fsm_stateReg)
      ports_0_fsm_enumDef_POWER_OFF : begin
      end
      ports_0_fsm_enumDef_DISCONNECTED : begin
      end
      ports_0_fsm_enumDef_DISABLED : begin
      end
      ports_0_fsm_enumDef_RESETTING : begin
      end
      ports_0_fsm_enumDef_RESETTING_DELAY : begin
      end
      ports_0_fsm_enumDef_RESETTING_SYNC : begin
      end
      ports_0_fsm_enumDef_ENABLED : begin
      end
      ports_0_fsm_enumDef_SUSPENDED : begin
      end
      ports_0_fsm_enumDef_RESUMING : begin
      end
      ports_0_fsm_enumDef_SEND_EOP_0 : begin
      end
      ports_0_fsm_enumDef_SEND_EOP_1 : begin
      end
      ports_0_fsm_enumDef_RESTART_S : begin
      end
      ports_0_fsm_enumDef_RESTART_E : begin
      end
      default : begin
        ports_0_fsm_wantStart = 1'b1;
      end
    endcase
  end

  assign ports_0_fsm_wantKill = 1'b0;
  always @(*) begin
    ports_0_fsm_timer_clear = 1'b0;
    case(ports_0_fsm_stateReg)
      ports_0_fsm_enumDef_POWER_OFF : begin
      end
      ports_0_fsm_enumDef_DISCONNECTED : begin
        if(when_usbphy_l540) begin
          ports_0_fsm_timer_clear = 1'b1;
        end
      end
      ports_0_fsm_enumDef_DISABLED : begin
      end
      ports_0_fsm_enumDef_RESETTING : begin
      end
      ports_0_fsm_enumDef_RESETTING_DELAY : begin
      end
      ports_0_fsm_enumDef_RESETTING_SYNC : begin
      end
      ports_0_fsm_enumDef_ENABLED : begin
      end
      ports_0_fsm_enumDef_SUSPENDED : begin
      end
      ports_0_fsm_enumDef_RESUMING : begin
      end
      ports_0_fsm_enumDef_SEND_EOP_0 : begin
      end
      ports_0_fsm_enumDef_SEND_EOP_1 : begin
      end
      ports_0_fsm_enumDef_RESTART_S : begin
      end
      ports_0_fsm_enumDef_RESTART_E : begin
      end
      default : begin
      end
    endcase
    if(when_StateMachine_l253_2) begin
      ports_0_fsm_timer_clear = 1'b1;
    end
    if(when_StateMachine_l253_3) begin
      ports_0_fsm_timer_clear = 1'b1;
    end
    if(when_StateMachine_l253_4) begin
      ports_0_fsm_timer_clear = 1'b1;
    end
    if(when_StateMachine_l253_5) begin
      ports_0_fsm_timer_clear = 1'b1;
    end
    if(when_StateMachine_l253_6) begin
      ports_0_fsm_timer_clear = 1'b1;
    end
    if(when_StateMachine_l253_7) begin
      ports_0_fsm_timer_clear = 1'b1;
    end
    if(when_StateMachine_l253_8) begin
      ports_0_fsm_timer_clear = 1'b1;
    end
    if(when_StateMachine_l253_9) begin
      ports_0_fsm_timer_clear = 1'b1;
    end
  end

  assign ports_0_fsm_timer_inc = 1'b1;
  assign ports_0_fsm_timer_DISCONNECTED_EOI = (ports_0_fsm_timer_counter == 24'h005dbf);
  assign ports_0_fsm_timer_RESET_DELAY = (ports_0_fsm_timer_counter == 24'h00095f);
  assign ports_0_fsm_timer_RESET_EOI = (ports_0_fsm_timer_counter == 24'h249eff);
  assign ports_0_fsm_timer_RESUME_EOI = (ports_0_fsm_timer_counter == 24'h0f617f);
  assign ports_0_fsm_timer_RESTART_EOI = (ports_0_fsm_timer_counter == 24'h0012bf);
  assign ports_0_fsm_timer_ONE_BIT = (ports_0_fsm_timer_counter == _zz_ports_0_fsm_timer_ONE_BIT);
  assign ports_0_fsm_timer_TWO_BIT = (ports_0_fsm_timer_counter == _zz_ports_0_fsm_timer_TWO_BIT);
  always @(*) begin
    ports_0_fsm_timer_lowSpeed = ports_0_portLowSpeed;
    case(ports_0_fsm_stateReg)
      ports_0_fsm_enumDef_POWER_OFF : begin
      end
      ports_0_fsm_enumDef_DISCONNECTED : begin
      end
      ports_0_fsm_enumDef_DISABLED : begin
      end
      ports_0_fsm_enumDef_RESETTING : begin
      end
      ports_0_fsm_enumDef_RESETTING_DELAY : begin
      end
      ports_0_fsm_enumDef_RESETTING_SYNC : begin
      end
      ports_0_fsm_enumDef_ENABLED : begin
      end
      ports_0_fsm_enumDef_SUSPENDED : begin
      end
      ports_0_fsm_enumDef_RESUMING : begin
      end
      ports_0_fsm_enumDef_SEND_EOP_0 : begin
        if(ports_0_fsm_lowSpeedEop) begin
          ports_0_fsm_timer_lowSpeed = 1'b1;
        end
      end
      ports_0_fsm_enumDef_SEND_EOP_1 : begin
        if(ports_0_fsm_lowSpeedEop) begin
          ports_0_fsm_timer_lowSpeed = 1'b1;
        end
      end
      ports_0_fsm_enumDef_RESTART_S : begin
      end
      ports_0_fsm_enumDef_RESTART_E : begin
      end
      default : begin
      end
    endcase
  end

  assign io_ctrl_ports_0_disable_ready = 1'b1;
  always @(*) begin
    io_ctrl_ports_0_reset_ready = 1'b0;
    case(ports_0_fsm_stateReg)
      ports_0_fsm_enumDef_POWER_OFF : begin
      end
      ports_0_fsm_enumDef_DISCONNECTED : begin
      end
      ports_0_fsm_enumDef_DISABLED : begin
      end
      ports_0_fsm_enumDef_RESETTING : begin
      end
      ports_0_fsm_enumDef_RESETTING_DELAY : begin
      end
      ports_0_fsm_enumDef_RESETTING_SYNC : begin
        if(when_usbphy_l580) begin
          io_ctrl_ports_0_reset_ready = 1'b1;
        end
      end
      ports_0_fsm_enumDef_ENABLED : begin
      end
      ports_0_fsm_enumDef_SUSPENDED : begin
      end
      ports_0_fsm_enumDef_RESUMING : begin
      end
      ports_0_fsm_enumDef_SEND_EOP_0 : begin
      end
      ports_0_fsm_enumDef_SEND_EOP_1 : begin
      end
      ports_0_fsm_enumDef_RESTART_S : begin
      end
      ports_0_fsm_enumDef_RESTART_E : begin
      end
      default : begin
      end
    endcase
  end

  assign io_ctrl_ports_0_resume_ready = 1'b1;
  assign io_ctrl_ports_0_suspend_ready = 1'b1;
  always @(*) begin
    io_ctrl_ports_0_connect = 1'b0;
    case(ports_0_fsm_stateReg)
      ports_0_fsm_enumDef_POWER_OFF : begin
      end
      ports_0_fsm_enumDef_DISCONNECTED : begin
        if(ports_0_fsm_timer_DISCONNECTED_EOI) begin
          io_ctrl_ports_0_connect = 1'b1;
        end
      end
      ports_0_fsm_enumDef_DISABLED : begin
      end
      ports_0_fsm_enumDef_RESETTING : begin
      end
      ports_0_fsm_enumDef_RESETTING_DELAY : begin
      end
      ports_0_fsm_enumDef_RESETTING_SYNC : begin
      end
      ports_0_fsm_enumDef_ENABLED : begin
      end
      ports_0_fsm_enumDef_SUSPENDED : begin
      end
      ports_0_fsm_enumDef_RESUMING : begin
      end
      ports_0_fsm_enumDef_SEND_EOP_0 : begin
      end
      ports_0_fsm_enumDef_SEND_EOP_1 : begin
      end
      ports_0_fsm_enumDef_RESTART_S : begin
      end
      ports_0_fsm_enumDef_RESTART_E : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    io_usb_0_tx_enable = 1'b0;
    case(ports_0_fsm_stateReg)
      ports_0_fsm_enumDef_POWER_OFF : begin
        io_usb_0_tx_enable = 1'b1;
      end
      ports_0_fsm_enumDef_DISCONNECTED : begin
      end
      ports_0_fsm_enumDef_DISABLED : begin
      end
      ports_0_fsm_enumDef_RESETTING : begin
        io_usb_0_tx_enable = 1'b1;
      end
      ports_0_fsm_enumDef_RESETTING_DELAY : begin
      end
      ports_0_fsm_enumDef_RESETTING_SYNC : begin
      end
      ports_0_fsm_enumDef_ENABLED : begin
        io_usb_0_tx_enable = txShared_encoder_output_valid;
        if(when_usbphy_l593) begin
          io_usb_0_tx_enable = txShared_lowSpeedSof_valid;
        end
      end
      ports_0_fsm_enumDef_SUSPENDED : begin
      end
      ports_0_fsm_enumDef_RESUMING : begin
        io_usb_0_tx_enable = 1'b1;
      end
      ports_0_fsm_enumDef_SEND_EOP_0 : begin
        io_usb_0_tx_enable = 1'b1;
      end
      ports_0_fsm_enumDef_SEND_EOP_1 : begin
        io_usb_0_tx_enable = 1'b1;
      end
      ports_0_fsm_enumDef_RESTART_S : begin
      end
      ports_0_fsm_enumDef_RESTART_E : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    io_usb_0_tx_data = 1'bx;
    case(ports_0_fsm_stateReg)
      ports_0_fsm_enumDef_POWER_OFF : begin
      end
      ports_0_fsm_enumDef_DISCONNECTED : begin
      end
      ports_0_fsm_enumDef_DISABLED : begin
      end
      ports_0_fsm_enumDef_RESETTING : begin
      end
      ports_0_fsm_enumDef_RESETTING_DELAY : begin
      end
      ports_0_fsm_enumDef_RESETTING_SYNC : begin
      end
      ports_0_fsm_enumDef_ENABLED : begin
        io_usb_0_tx_data = ((txShared_encoder_output_data || ports_0_fsm_forceJ) ^ ports_0_portLowSpeed);
        if(when_usbphy_l593) begin
          io_usb_0_tx_data = txShared_lowSpeedSof_data;
        end
      end
      ports_0_fsm_enumDef_SUSPENDED : begin
      end
      ports_0_fsm_enumDef_RESUMING : begin
        io_usb_0_tx_data = ports_0_portLowSpeed;
      end
      ports_0_fsm_enumDef_SEND_EOP_0 : begin
      end
      ports_0_fsm_enumDef_SEND_EOP_1 : begin
        io_usb_0_tx_data = (! ports_0_portLowSpeed);
      end
      ports_0_fsm_enumDef_RESTART_S : begin
      end
      ports_0_fsm_enumDef_RESTART_E : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    io_usb_0_tx_se0 = 1'bx;
    case(ports_0_fsm_stateReg)
      ports_0_fsm_enumDef_POWER_OFF : begin
        io_usb_0_tx_se0 = 1'b1;
      end
      ports_0_fsm_enumDef_DISCONNECTED : begin
      end
      ports_0_fsm_enumDef_DISABLED : begin
      end
      ports_0_fsm_enumDef_RESETTING : begin
        io_usb_0_tx_se0 = 1'b1;
      end
      ports_0_fsm_enumDef_RESETTING_DELAY : begin
      end
      ports_0_fsm_enumDef_RESETTING_SYNC : begin
      end
      ports_0_fsm_enumDef_ENABLED : begin
        io_usb_0_tx_se0 = (txShared_encoder_output_se0 && (! ports_0_fsm_forceJ));
        if(when_usbphy_l593) begin
          io_usb_0_tx_se0 = txShared_lowSpeedSof_se0;
        end
      end
      ports_0_fsm_enumDef_SUSPENDED : begin
      end
      ports_0_fsm_enumDef_RESUMING : begin
        io_usb_0_tx_se0 = 1'b0;
      end
      ports_0_fsm_enumDef_SEND_EOP_0 : begin
        io_usb_0_tx_se0 = 1'b1;
      end
      ports_0_fsm_enumDef_SEND_EOP_1 : begin
        io_usb_0_tx_se0 = 1'b0;
      end
      ports_0_fsm_enumDef_RESTART_S : begin
      end
      ports_0_fsm_enumDef_RESTART_E : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    ports_0_fsm_resetInProgress = 1'b0;
    case(ports_0_fsm_stateReg)
      ports_0_fsm_enumDef_POWER_OFF : begin
      end
      ports_0_fsm_enumDef_DISCONNECTED : begin
      end
      ports_0_fsm_enumDef_DISABLED : begin
      end
      ports_0_fsm_enumDef_RESETTING : begin
        ports_0_fsm_resetInProgress = 1'b1;
      end
      ports_0_fsm_enumDef_RESETTING_DELAY : begin
        ports_0_fsm_resetInProgress = 1'b1;
      end
      ports_0_fsm_enumDef_RESETTING_SYNC : begin
        ports_0_fsm_resetInProgress = 1'b1;
      end
      ports_0_fsm_enumDef_ENABLED : begin
      end
      ports_0_fsm_enumDef_SUSPENDED : begin
      end
      ports_0_fsm_enumDef_RESUMING : begin
      end
      ports_0_fsm_enumDef_SEND_EOP_0 : begin
      end
      ports_0_fsm_enumDef_SEND_EOP_1 : begin
      end
      ports_0_fsm_enumDef_RESTART_S : begin
      end
      ports_0_fsm_enumDef_RESTART_E : begin
      end
      default : begin
      end
    endcase
  end

  assign ports_0_fsm_forceJ = (ports_0_portLowSpeed && (! txShared_encoder_output_lowSpeed));
  assign when_usbphy_l672 = (&{(! (ports_0_fsm_stateReg == ports_0_fsm_enumDef_DISABLED)),{(! (ports_0_fsm_stateReg == ports_0_fsm_enumDef_SUSPENDED)),(! (ports_0_fsm_stateReg == ports_0_fsm_enumDef_ENABLED))}});
  assign io_ctrl_ports_1_lowSpeed = ports_1_portLowSpeed;
  assign io_ctrl_ports_1_remoteResume = 1'b0;
  always @(*) begin
    ports_1_rx_enablePackets = 1'b0;
    case(ports_1_fsm_stateReg)
      ports_1_fsm_enumDef_POWER_OFF : begin
      end
      ports_1_fsm_enumDef_DISCONNECTED : begin
      end
      ports_1_fsm_enumDef_DISABLED : begin
      end
      ports_1_fsm_enumDef_RESETTING : begin
      end
      ports_1_fsm_enumDef_RESETTING_DELAY : begin
      end
      ports_1_fsm_enumDef_RESETTING_SYNC : begin
      end
      ports_1_fsm_enumDef_ENABLED : begin
        ports_1_rx_enablePackets = 1'b1;
      end
      ports_1_fsm_enumDef_SUSPENDED : begin
      end
      ports_1_fsm_enumDef_RESUMING : begin
      end
      ports_1_fsm_enumDef_SEND_EOP_0 : begin
      end
      ports_1_fsm_enumDef_SEND_EOP_1 : begin
      end
      ports_1_fsm_enumDef_RESTART_S : begin
      end
      ports_1_fsm_enumDef_RESTART_E : begin
      end
      default : begin
      end
    endcase
  end

  assign ports_1_rx_j = ((ports_1_filter_io_filtred_dp == (! ports_1_portLowSpeed)) && (ports_1_filter_io_filtred_dm == ports_1_portLowSpeed));
  assign ports_1_rx_k = ((ports_1_filter_io_filtred_dp == ports_1_portLowSpeed) && (ports_1_filter_io_filtred_dm == (! ports_1_portLowSpeed)));
  assign io_management_1_power = io_ctrl_ports_1_power;
  assign io_ctrl_ports_1_overcurrent = io_management_1_overcurrent;
  always @(*) begin
    ports_1_rx_waitSync = 1'b0;
    case(ports_1_rx_packet_stateReg)
      ports_1_rx_packet_enumDef_IDLE : begin
        ports_1_rx_waitSync = 1'b1;
      end
      ports_1_rx_packet_enumDef_PACKET : begin
      end
      ports_1_rx_packet_enumDef_ERRORED : begin
      end
      default : begin
      end
    endcase
    if(when_StateMachine_l253_10) begin
      ports_1_rx_waitSync = 1'b1;
    end
  end

  always @(*) begin
    ports_1_rx_decoder_output_valid = 1'b0;
    if(ports_1_filter_io_filtred_sample) begin
      ports_1_rx_decoder_output_valid = 1'b1;
    end
  end

  always @(*) begin
    ports_1_rx_decoder_output_payload = 1'bx;
    if(ports_1_filter_io_filtred_sample) begin
      if(when_usbphy_l347_1) begin
        ports_1_rx_decoder_output_payload = 1'b0;
      end else begin
        ports_1_rx_decoder_output_payload = 1'b1;
      end
    end
  end

  assign when_usbphy_l347_1 = ((ports_1_rx_decoder_state ^ ports_1_filter_io_filtred_d) ^ ports_1_portLowSpeed);
  assign ports_1_rx_destuffer_unstuffNext = (ports_1_rx_destuffer_counter == 3'b110);
  assign ports_1_rx_destuffer_output_valid = (ports_1_rx_decoder_output_valid && (! ports_1_rx_destuffer_unstuffNext));
  assign ports_1_rx_destuffer_output_payload = ports_1_rx_decoder_output_payload;
  assign when_usbphy_l368_1 = ((! ports_1_rx_decoder_output_payload) || ports_1_rx_destuffer_unstuffNext);
  assign ports_1_rx_history_updated = ports_1_rx_destuffer_output_valid;
  assign _zz_ports_1_rx_history_value = ports_1_rx_destuffer_output_payload;
  assign ports_1_rx_history_value = {_zz_ports_1_rx_history_value,{_zz_ports_1_rx_history_value_1,{_zz_ports_1_rx_history_value_2,{_zz_ports_1_rx_history_value_3,{_zz_ports_1_rx_history_value_4,{_zz_ports_1_rx_history_value_5,{_zz_ports_1_rx_history_value_6,_zz_ports_1_rx_history_value_7}}}}}}};
  assign ports_1_rx_history_sync_hit = (ports_1_rx_history_updated && (ports_1_rx_history_value == 8'hd5));
  assign ports_1_rx_eop_maxThreshold = (io_ctrl_lowSpeed ? 7'h60 : 7'h0c);
  assign ports_1_rx_eop_minThreshold = (io_ctrl_lowSpeed ? 6'h2a : 6'h05);
  assign ports_1_rx_eop_maxHit = (ports_1_rx_eop_counter == ports_1_rx_eop_maxThreshold);
  always @(*) begin
    ports_1_rx_eop_hit = 1'b0;
    if(ports_1_rx_j) begin
      if(when_usbphy_l403_1) begin
        ports_1_rx_eop_hit = 1'b1;
      end
    end
  end

  assign when_usbphy_l395_1 = ((! ports_1_filter_io_filtred_dp) && (! ports_1_filter_io_filtred_dm));
  assign when_usbphy_l396_1 = (! ports_1_rx_eop_maxHit);
  assign when_usbphy_l403_1 = ((_zz_when_usbphy_l403_1 <= ports_1_rx_eop_counter) && (! ports_1_rx_eop_maxHit));
  assign ports_1_rx_packet_wantExit = 1'b0;
  always @(*) begin
    ports_1_rx_packet_wantStart = 1'b0;
    case(ports_1_rx_packet_stateReg)
      ports_1_rx_packet_enumDef_IDLE : begin
      end
      ports_1_rx_packet_enumDef_PACKET : begin
      end
      ports_1_rx_packet_enumDef_ERRORED : begin
      end
      default : begin
        ports_1_rx_packet_wantStart = 1'b1;
      end
    endcase
  end

  assign ports_1_rx_packet_wantKill = 1'b0;
  always @(*) begin
    ports_1_rx_packet_errorTimeout_clear = 1'b0;
    case(ports_1_rx_packet_stateReg)
      ports_1_rx_packet_enumDef_IDLE : begin
      end
      ports_1_rx_packet_enumDef_PACKET : begin
      end
      ports_1_rx_packet_enumDef_ERRORED : begin
        if(when_usbphy_l451_1) begin
          ports_1_rx_packet_errorTimeout_clear = 1'b1;
        end
      end
      default : begin
      end
    endcase
    if(when_StateMachine_l253_11) begin
      ports_1_rx_packet_errorTimeout_clear = 1'b1;
    end
  end

  assign ports_1_rx_packet_errorTimeout_inc = 1'b1;
  assign ports_1_rx_packet_errorTimeout_lowSpeed = io_ctrl_lowSpeed;
  assign ports_1_rx_packet_errorTimeout_trigger = (ports_1_rx_packet_errorTimeout_counter == _zz_ports_1_rx_packet_errorTimeout_trigger);
  always @(*) begin
    ports_1_rx_disconnect_clear = 1'b0;
    if(when_usbphy_l475_1) begin
      ports_1_rx_disconnect_clear = 1'b1;
    end
    if(when_usbphy_l672_1) begin
      ports_1_rx_disconnect_clear = 1'b1;
    end
  end

  assign ports_1_rx_disconnect_hit = (ports_1_rx_disconnect_counter == 7'h68);
  assign ports_1_rx_disconnect_event = (ports_1_rx_disconnect_hit && (! ports_1_rx_disconnect_hitLast));
  assign when_usbphy_l475_1 = ((! ports_1_filter_io_filtred_se0) || io_usb_1_tx_enable);
  assign io_ctrl_ports_1_disconnect = ports_1_rx_disconnect_event;
  assign ports_1_fsm_wantExit = 1'b0;
  always @(*) begin
    ports_1_fsm_wantStart = 1'b0;
    case(ports_1_fsm_stateReg)
      ports_1_fsm_enumDef_POWER_OFF : begin
      end
      ports_1_fsm_enumDef_DISCONNECTED : begin
      end
      ports_1_fsm_enumDef_DISABLED : begin
      end
      ports_1_fsm_enumDef_RESETTING : begin
      end
      ports_1_fsm_enumDef_RESETTING_DELAY : begin
      end
      ports_1_fsm_enumDef_RESETTING_SYNC : begin
      end
      ports_1_fsm_enumDef_ENABLED : begin
      end
      ports_1_fsm_enumDef_SUSPENDED : begin
      end
      ports_1_fsm_enumDef_RESUMING : begin
      end
      ports_1_fsm_enumDef_SEND_EOP_0 : begin
      end
      ports_1_fsm_enumDef_SEND_EOP_1 : begin
      end
      ports_1_fsm_enumDef_RESTART_S : begin
      end
      ports_1_fsm_enumDef_RESTART_E : begin
      end
      default : begin
        ports_1_fsm_wantStart = 1'b1;
      end
    endcase
  end

  assign ports_1_fsm_wantKill = 1'b0;
  always @(*) begin
    ports_1_fsm_timer_clear = 1'b0;
    case(ports_1_fsm_stateReg)
      ports_1_fsm_enumDef_POWER_OFF : begin
      end
      ports_1_fsm_enumDef_DISCONNECTED : begin
        if(when_usbphy_l540_1) begin
          ports_1_fsm_timer_clear = 1'b1;
        end
      end
      ports_1_fsm_enumDef_DISABLED : begin
      end
      ports_1_fsm_enumDef_RESETTING : begin
      end
      ports_1_fsm_enumDef_RESETTING_DELAY : begin
      end
      ports_1_fsm_enumDef_RESETTING_SYNC : begin
      end
      ports_1_fsm_enumDef_ENABLED : begin
      end
      ports_1_fsm_enumDef_SUSPENDED : begin
      end
      ports_1_fsm_enumDef_RESUMING : begin
      end
      ports_1_fsm_enumDef_SEND_EOP_0 : begin
      end
      ports_1_fsm_enumDef_SEND_EOP_1 : begin
      end
      ports_1_fsm_enumDef_RESTART_S : begin
      end
      ports_1_fsm_enumDef_RESTART_E : begin
      end
      default : begin
      end
    endcase
    if(when_StateMachine_l253_12) begin
      ports_1_fsm_timer_clear = 1'b1;
    end
    if(when_StateMachine_l253_13) begin
      ports_1_fsm_timer_clear = 1'b1;
    end
    if(when_StateMachine_l253_14) begin
      ports_1_fsm_timer_clear = 1'b1;
    end
    if(when_StateMachine_l253_15) begin
      ports_1_fsm_timer_clear = 1'b1;
    end
    if(when_StateMachine_l253_16) begin
      ports_1_fsm_timer_clear = 1'b1;
    end
    if(when_StateMachine_l253_17) begin
      ports_1_fsm_timer_clear = 1'b1;
    end
    if(when_StateMachine_l253_18) begin
      ports_1_fsm_timer_clear = 1'b1;
    end
    if(when_StateMachine_l253_19) begin
      ports_1_fsm_timer_clear = 1'b1;
    end
  end

  assign ports_1_fsm_timer_inc = 1'b1;
  assign ports_1_fsm_timer_DISCONNECTED_EOI = (ports_1_fsm_timer_counter == 24'h005dbf);
  assign ports_1_fsm_timer_RESET_DELAY = (ports_1_fsm_timer_counter == 24'h00095f);
  assign ports_1_fsm_timer_RESET_EOI = (ports_1_fsm_timer_counter == 24'h249eff);
  assign ports_1_fsm_timer_RESUME_EOI = (ports_1_fsm_timer_counter == 24'h0f617f);
  assign ports_1_fsm_timer_RESTART_EOI = (ports_1_fsm_timer_counter == 24'h0012bf);
  assign ports_1_fsm_timer_ONE_BIT = (ports_1_fsm_timer_counter == _zz_ports_1_fsm_timer_ONE_BIT);
  assign ports_1_fsm_timer_TWO_BIT = (ports_1_fsm_timer_counter == _zz_ports_1_fsm_timer_TWO_BIT);
  always @(*) begin
    ports_1_fsm_timer_lowSpeed = ports_1_portLowSpeed;
    case(ports_1_fsm_stateReg)
      ports_1_fsm_enumDef_POWER_OFF : begin
      end
      ports_1_fsm_enumDef_DISCONNECTED : begin
      end
      ports_1_fsm_enumDef_DISABLED : begin
      end
      ports_1_fsm_enumDef_RESETTING : begin
      end
      ports_1_fsm_enumDef_RESETTING_DELAY : begin
      end
      ports_1_fsm_enumDef_RESETTING_SYNC : begin
      end
      ports_1_fsm_enumDef_ENABLED : begin
      end
      ports_1_fsm_enumDef_SUSPENDED : begin
      end
      ports_1_fsm_enumDef_RESUMING : begin
      end
      ports_1_fsm_enumDef_SEND_EOP_0 : begin
        if(ports_1_fsm_lowSpeedEop) begin
          ports_1_fsm_timer_lowSpeed = 1'b1;
        end
      end
      ports_1_fsm_enumDef_SEND_EOP_1 : begin
        if(ports_1_fsm_lowSpeedEop) begin
          ports_1_fsm_timer_lowSpeed = 1'b1;
        end
      end
      ports_1_fsm_enumDef_RESTART_S : begin
      end
      ports_1_fsm_enumDef_RESTART_E : begin
      end
      default : begin
      end
    endcase
  end

  assign io_ctrl_ports_1_disable_ready = 1'b1;
  always @(*) begin
    io_ctrl_ports_1_reset_ready = 1'b0;
    case(ports_1_fsm_stateReg)
      ports_1_fsm_enumDef_POWER_OFF : begin
      end
      ports_1_fsm_enumDef_DISCONNECTED : begin
      end
      ports_1_fsm_enumDef_DISABLED : begin
      end
      ports_1_fsm_enumDef_RESETTING : begin
      end
      ports_1_fsm_enumDef_RESETTING_DELAY : begin
      end
      ports_1_fsm_enumDef_RESETTING_SYNC : begin
        if(when_usbphy_l580_1) begin
          io_ctrl_ports_1_reset_ready = 1'b1;
        end
      end
      ports_1_fsm_enumDef_ENABLED : begin
      end
      ports_1_fsm_enumDef_SUSPENDED : begin
      end
      ports_1_fsm_enumDef_RESUMING : begin
      end
      ports_1_fsm_enumDef_SEND_EOP_0 : begin
      end
      ports_1_fsm_enumDef_SEND_EOP_1 : begin
      end
      ports_1_fsm_enumDef_RESTART_S : begin
      end
      ports_1_fsm_enumDef_RESTART_E : begin
      end
      default : begin
      end
    endcase
  end

  assign io_ctrl_ports_1_resume_ready = 1'b1;
  assign io_ctrl_ports_1_suspend_ready = 1'b1;
  always @(*) begin
    io_ctrl_ports_1_connect = 1'b0;
    case(ports_1_fsm_stateReg)
      ports_1_fsm_enumDef_POWER_OFF : begin
      end
      ports_1_fsm_enumDef_DISCONNECTED : begin
        if(ports_1_fsm_timer_DISCONNECTED_EOI) begin
          io_ctrl_ports_1_connect = 1'b1;
        end
      end
      ports_1_fsm_enumDef_DISABLED : begin
      end
      ports_1_fsm_enumDef_RESETTING : begin
      end
      ports_1_fsm_enumDef_RESETTING_DELAY : begin
      end
      ports_1_fsm_enumDef_RESETTING_SYNC : begin
      end
      ports_1_fsm_enumDef_ENABLED : begin
      end
      ports_1_fsm_enumDef_SUSPENDED : begin
      end
      ports_1_fsm_enumDef_RESUMING : begin
      end
      ports_1_fsm_enumDef_SEND_EOP_0 : begin
      end
      ports_1_fsm_enumDef_SEND_EOP_1 : begin
      end
      ports_1_fsm_enumDef_RESTART_S : begin
      end
      ports_1_fsm_enumDef_RESTART_E : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    io_usb_1_tx_enable = 1'b0;
    case(ports_1_fsm_stateReg)
      ports_1_fsm_enumDef_POWER_OFF : begin
        io_usb_1_tx_enable = 1'b1;
      end
      ports_1_fsm_enumDef_DISCONNECTED : begin
      end
      ports_1_fsm_enumDef_DISABLED : begin
      end
      ports_1_fsm_enumDef_RESETTING : begin
        io_usb_1_tx_enable = 1'b1;
      end
      ports_1_fsm_enumDef_RESETTING_DELAY : begin
      end
      ports_1_fsm_enumDef_RESETTING_SYNC : begin
      end
      ports_1_fsm_enumDef_ENABLED : begin
        io_usb_1_tx_enable = txShared_encoder_output_valid;
        if(when_usbphy_l593_1) begin
          io_usb_1_tx_enable = txShared_lowSpeedSof_valid;
        end
      end
      ports_1_fsm_enumDef_SUSPENDED : begin
      end
      ports_1_fsm_enumDef_RESUMING : begin
        io_usb_1_tx_enable = 1'b1;
      end
      ports_1_fsm_enumDef_SEND_EOP_0 : begin
        io_usb_1_tx_enable = 1'b1;
      end
      ports_1_fsm_enumDef_SEND_EOP_1 : begin
        io_usb_1_tx_enable = 1'b1;
      end
      ports_1_fsm_enumDef_RESTART_S : begin
      end
      ports_1_fsm_enumDef_RESTART_E : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    io_usb_1_tx_data = 1'bx;
    case(ports_1_fsm_stateReg)
      ports_1_fsm_enumDef_POWER_OFF : begin
      end
      ports_1_fsm_enumDef_DISCONNECTED : begin
      end
      ports_1_fsm_enumDef_DISABLED : begin
      end
      ports_1_fsm_enumDef_RESETTING : begin
      end
      ports_1_fsm_enumDef_RESETTING_DELAY : begin
      end
      ports_1_fsm_enumDef_RESETTING_SYNC : begin
      end
      ports_1_fsm_enumDef_ENABLED : begin
        io_usb_1_tx_data = ((txShared_encoder_output_data || ports_1_fsm_forceJ) ^ ports_1_portLowSpeed);
        if(when_usbphy_l593_1) begin
          io_usb_1_tx_data = txShared_lowSpeedSof_data;
        end
      end
      ports_1_fsm_enumDef_SUSPENDED : begin
      end
      ports_1_fsm_enumDef_RESUMING : begin
        io_usb_1_tx_data = ports_1_portLowSpeed;
      end
      ports_1_fsm_enumDef_SEND_EOP_0 : begin
      end
      ports_1_fsm_enumDef_SEND_EOP_1 : begin
        io_usb_1_tx_data = (! ports_1_portLowSpeed);
      end
      ports_1_fsm_enumDef_RESTART_S : begin
      end
      ports_1_fsm_enumDef_RESTART_E : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    io_usb_1_tx_se0 = 1'bx;
    case(ports_1_fsm_stateReg)
      ports_1_fsm_enumDef_POWER_OFF : begin
        io_usb_1_tx_se0 = 1'b1;
      end
      ports_1_fsm_enumDef_DISCONNECTED : begin
      end
      ports_1_fsm_enumDef_DISABLED : begin
      end
      ports_1_fsm_enumDef_RESETTING : begin
        io_usb_1_tx_se0 = 1'b1;
      end
      ports_1_fsm_enumDef_RESETTING_DELAY : begin
      end
      ports_1_fsm_enumDef_RESETTING_SYNC : begin
      end
      ports_1_fsm_enumDef_ENABLED : begin
        io_usb_1_tx_se0 = (txShared_encoder_output_se0 && (! ports_1_fsm_forceJ));
        if(when_usbphy_l593_1) begin
          io_usb_1_tx_se0 = txShared_lowSpeedSof_se0;
        end
      end
      ports_1_fsm_enumDef_SUSPENDED : begin
      end
      ports_1_fsm_enumDef_RESUMING : begin
        io_usb_1_tx_se0 = 1'b0;
      end
      ports_1_fsm_enumDef_SEND_EOP_0 : begin
        io_usb_1_tx_se0 = 1'b1;
      end
      ports_1_fsm_enumDef_SEND_EOP_1 : begin
        io_usb_1_tx_se0 = 1'b0;
      end
      ports_1_fsm_enumDef_RESTART_S : begin
      end
      ports_1_fsm_enumDef_RESTART_E : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    ports_1_fsm_resetInProgress = 1'b0;
    case(ports_1_fsm_stateReg)
      ports_1_fsm_enumDef_POWER_OFF : begin
      end
      ports_1_fsm_enumDef_DISCONNECTED : begin
      end
      ports_1_fsm_enumDef_DISABLED : begin
      end
      ports_1_fsm_enumDef_RESETTING : begin
        ports_1_fsm_resetInProgress = 1'b1;
      end
      ports_1_fsm_enumDef_RESETTING_DELAY : begin
        ports_1_fsm_resetInProgress = 1'b1;
      end
      ports_1_fsm_enumDef_RESETTING_SYNC : begin
        ports_1_fsm_resetInProgress = 1'b1;
      end
      ports_1_fsm_enumDef_ENABLED : begin
      end
      ports_1_fsm_enumDef_SUSPENDED : begin
      end
      ports_1_fsm_enumDef_RESUMING : begin
      end
      ports_1_fsm_enumDef_SEND_EOP_0 : begin
      end
      ports_1_fsm_enumDef_SEND_EOP_1 : begin
      end
      ports_1_fsm_enumDef_RESTART_S : begin
      end
      ports_1_fsm_enumDef_RESTART_E : begin
      end
      default : begin
      end
    endcase
  end

  assign ports_1_fsm_forceJ = (ports_1_portLowSpeed && (! txShared_encoder_output_lowSpeed));
  assign when_usbphy_l672_1 = (&{(! (ports_1_fsm_stateReg == ports_1_fsm_enumDef_DISABLED)),{(! (ports_1_fsm_stateReg == ports_1_fsm_enumDef_SUSPENDED)),(! (ports_1_fsm_stateReg == ports_1_fsm_enumDef_ENABLED))}});
  always @(*) begin
    txShared_frame_stateNext = txShared_frame_stateReg;
    case(txShared_frame_stateReg)
      txShared_frame_enumDef_IDLE : begin
        if(when_usbphy_l191) begin
          txShared_frame_stateNext = txShared_frame_enumDef_TAKE_LINE;
        end
      end
      txShared_frame_enumDef_TAKE_LINE : begin
        if(txShared_timer_oneCycle) begin
          if(io_ctrl_lowSpeed) begin
            txShared_frame_stateNext = txShared_frame_enumDef_PREAMBLE_SYNC;
          end else begin
            txShared_frame_stateNext = txShared_frame_enumDef_SYNC;
          end
        end
      end
      txShared_frame_enumDef_PREAMBLE_SYNC : begin
        if(txShared_serialiser_input_ready) begin
          txShared_frame_stateNext = txShared_frame_enumDef_PREAMBLE_PID;
        end
      end
      txShared_frame_enumDef_PREAMBLE_PID : begin
        if(txShared_serialiser_input_ready) begin
          txShared_frame_stateNext = txShared_frame_enumDef_PREAMBLE_DELAY;
        end
      end
      txShared_frame_enumDef_PREAMBLE_DELAY : begin
        if(txShared_timer_fourCycle) begin
          txShared_frame_stateNext = txShared_frame_enumDef_SYNC;
        end
      end
      txShared_frame_enumDef_SYNC : begin
        if(txShared_serialiser_input_ready) begin
          txShared_frame_stateNext = txShared_frame_enumDef_DATA;
        end
      end
      txShared_frame_enumDef_DATA : begin
        if(txShared_serialiser_input_ready) begin
          if(io_ctrl_tx_payload_last) begin
            txShared_frame_stateNext = txShared_frame_enumDef_EOP_0;
          end
        end
      end
      txShared_frame_enumDef_EOP_0 : begin
        if(txShared_timer_twoCycle) begin
          txShared_frame_stateNext = txShared_frame_enumDef_EOP_1;
        end
      end
      txShared_frame_enumDef_EOP_1 : begin
        if(txShared_timer_oneCycle) begin
          txShared_frame_stateNext = txShared_frame_enumDef_EOP_2;
        end
      end
      txShared_frame_enumDef_EOP_2 : begin
        if(txShared_timer_twoCycle) begin
          txShared_frame_stateNext = txShared_frame_enumDef_IDLE;
        end
      end
      default : begin
      end
    endcase
    if(txShared_frame_wantStart) begin
      txShared_frame_stateNext = txShared_frame_enumDef_IDLE;
    end
    if(txShared_frame_wantKill) begin
      txShared_frame_stateNext = txShared_frame_enumDef_BOOT;
    end
  end

  assign when_usbphy_l191 = (io_ctrl_tx_valid && (! txShared_rxToTxDelay_active));
  always @(*) begin
    upstreamRx_stateNext = upstreamRx_stateReg;
    case(upstreamRx_stateReg)
      upstreamRx_enumDef_IDLE : begin
        if(upstreamRx_timer_IDLE_EOI) begin
          upstreamRx_stateNext = upstreamRx_enumDef_SUSPEND;
        end
      end
      upstreamRx_enumDef_SUSPEND : begin
        if(txShared_encoder_output_valid) begin
          upstreamRx_stateNext = upstreamRx_enumDef_IDLE;
        end
      end
      default : begin
      end
    endcase
    if(upstreamRx_wantStart) begin
      upstreamRx_stateNext = upstreamRx_enumDef_IDLE;
    end
    if(upstreamRx_wantKill) begin
      upstreamRx_stateNext = upstreamRx_enumDef_BOOT;
    end
  end

  assign Rx_Suspend = (upstreamRx_stateReg == upstreamRx_enumDef_SUSPEND);
  always @(*) begin
    ports_0_rx_packet_stateNext = ports_0_rx_packet_stateReg;
    case(ports_0_rx_packet_stateReg)
      ports_0_rx_packet_enumDef_IDLE : begin
        if(ports_0_rx_history_sync_hit) begin
          ports_0_rx_packet_stateNext = ports_0_rx_packet_enumDef_PACKET;
        end
      end
      ports_0_rx_packet_enumDef_PACKET : begin
        if(ports_0_rx_destuffer_output_valid) begin
          if(when_usbphy_l429) begin
            if(ports_0_rx_stuffingError) begin
              ports_0_rx_packet_stateNext = ports_0_rx_packet_enumDef_ERRORED;
            end
          end
        end
      end
      ports_0_rx_packet_enumDef_ERRORED : begin
        if(ports_0_rx_packet_errorTimeout_trigger) begin
          ports_0_rx_packet_stateNext = ports_0_rx_packet_enumDef_IDLE;
        end
      end
      default : begin
      end
    endcase
    if(ports_0_rx_eop_hit) begin
      ports_0_rx_packet_stateNext = ports_0_rx_packet_enumDef_IDLE;
    end
    if(txShared_encoder_output_valid) begin
      ports_0_rx_packet_stateNext = ports_0_rx_packet_enumDef_IDLE;
    end
    if(ports_0_rx_packet_wantStart) begin
      ports_0_rx_packet_stateNext = ports_0_rx_packet_enumDef_IDLE;
    end
    if(ports_0_rx_packet_wantKill) begin
      ports_0_rx_packet_stateNext = ports_0_rx_packet_enumDef_BOOT;
    end
  end

  assign when_usbphy_l429 = (ports_0_rx_packet_counter == 3'b111);
  assign when_usbphy_l451 = ((ports_0_rx_packet_errorTimeout_p != ports_0_filter_io_filtred_dp) || (ports_0_rx_packet_errorTimeout_n != ports_0_filter_io_filtred_dm));
  assign when_StateMachine_l253 = ((! (ports_0_rx_packet_stateReg == ports_0_rx_packet_enumDef_IDLE)) && (ports_0_rx_packet_stateNext == ports_0_rx_packet_enumDef_IDLE));
  assign when_StateMachine_l253_1 = ((! (ports_0_rx_packet_stateReg == ports_0_rx_packet_enumDef_ERRORED)) && (ports_0_rx_packet_stateNext == ports_0_rx_packet_enumDef_ERRORED));
  always @(*) begin
    ports_0_fsm_stateNext = ports_0_fsm_stateReg;
    case(ports_0_fsm_stateReg)
      ports_0_fsm_enumDef_POWER_OFF : begin
        if(io_ctrl_ports_0_power) begin
          ports_0_fsm_stateNext = ports_0_fsm_enumDef_DISCONNECTED;
        end
      end
      ports_0_fsm_enumDef_DISCONNECTED : begin
        if(ports_0_fsm_timer_DISCONNECTED_EOI) begin
          ports_0_fsm_stateNext = ports_0_fsm_enumDef_DISABLED;
        end
      end
      ports_0_fsm_enumDef_DISABLED : begin
      end
      ports_0_fsm_enumDef_RESETTING : begin
        if(ports_0_fsm_timer_RESET_EOI) begin
          ports_0_fsm_stateNext = ports_0_fsm_enumDef_RESETTING_DELAY;
        end
      end
      ports_0_fsm_enumDef_RESETTING_DELAY : begin
        if(ports_0_fsm_timer_RESET_DELAY) begin
          ports_0_fsm_stateNext = ports_0_fsm_enumDef_RESETTING_SYNC;
        end
      end
      ports_0_fsm_enumDef_RESETTING_SYNC : begin
        if(when_usbphy_l580) begin
          ports_0_fsm_stateNext = ports_0_fsm_enumDef_ENABLED;
        end
      end
      ports_0_fsm_enumDef_ENABLED : begin
        if(io_ctrl_ports_0_suspend_valid) begin
          ports_0_fsm_stateNext = ports_0_fsm_enumDef_SUSPENDED;
        end else begin
          if(when_usbphy_l602) begin
            ports_0_fsm_stateNext = ports_0_fsm_enumDef_RESTART_E;
          end else begin
            if(io_ctrl_usbResume) begin
              ports_0_fsm_stateNext = ports_0_fsm_enumDef_RESUMING;
            end
          end
        end
      end
      ports_0_fsm_enumDef_SUSPENDED : begin
        if(when_usbphy_l610) begin
          ports_0_fsm_stateNext = ports_0_fsm_enumDef_RESUMING;
        end else begin
          if(when_usbphy_l612) begin
            ports_0_fsm_stateNext = ports_0_fsm_enumDef_RESTART_S;
          end
        end
      end
      ports_0_fsm_enumDef_RESUMING : begin
        if(ports_0_fsm_timer_RESUME_EOI) begin
          ports_0_fsm_stateNext = ports_0_fsm_enumDef_SEND_EOP_0;
        end
      end
      ports_0_fsm_enumDef_SEND_EOP_0 : begin
        if(ports_0_fsm_timer_TWO_BIT) begin
          ports_0_fsm_stateNext = ports_0_fsm_enumDef_SEND_EOP_1;
        end
      end
      ports_0_fsm_enumDef_SEND_EOP_1 : begin
        if(ports_0_fsm_timer_ONE_BIT) begin
          ports_0_fsm_stateNext = ports_0_fsm_enumDef_ENABLED;
        end
      end
      ports_0_fsm_enumDef_RESTART_S : begin
        if(when_usbphy_l653) begin
          ports_0_fsm_stateNext = ports_0_fsm_enumDef_RESUMING;
        end
        if(ports_0_fsm_timer_RESTART_EOI) begin
          ports_0_fsm_stateNext = ports_0_fsm_enumDef_DISCONNECTED;
        end
      end
      ports_0_fsm_enumDef_RESTART_E : begin
        if(when_usbphy_l663) begin
          ports_0_fsm_stateNext = ports_0_fsm_enumDef_RESUMING;
        end
        if(ports_0_fsm_timer_RESTART_EOI) begin
          ports_0_fsm_stateNext = ports_0_fsm_enumDef_DISCONNECTED;
        end
      end
      default : begin
      end
    endcase
    if(when_usbphy_l512) begin
      ports_0_fsm_stateNext = ports_0_fsm_enumDef_POWER_OFF;
    end else begin
      if(ports_0_rx_disconnect_event) begin
        ports_0_fsm_stateNext = ports_0_fsm_enumDef_DISCONNECTED;
      end else begin
        if(io_ctrl_ports_0_disable_valid) begin
          ports_0_fsm_stateNext = ports_0_fsm_enumDef_DISABLED;
        end else begin
          if(io_ctrl_ports_0_reset_valid) begin
            if(when_usbphy_l519) begin
              if(when_usbphy_l520) begin
                ports_0_fsm_stateNext = ports_0_fsm_enumDef_RESETTING;
              end
            end
          end
        end
      end
    end
    if(ports_0_fsm_wantStart) begin
      ports_0_fsm_stateNext = ports_0_fsm_enumDef_POWER_OFF;
    end
    if(ports_0_fsm_wantKill) begin
      ports_0_fsm_stateNext = ports_0_fsm_enumDef_BOOT;
    end
  end

  assign when_usbphy_l540 = ((! ports_0_filter_io_filtred_dp) && (! ports_0_filter_io_filtred_dm));
  assign when_usbphy_l547 = ((! io_ctrl_ports_0_reset_valid) && (ports_0_filter_io_filtred_dm != ports_0_filter_io_filtred_dp));
  assign when_usbphy_l580 = (! txShared_encoder_output_valid);
  assign when_usbphy_l593 = (ports_0_portLowSpeed && txShared_lowSpeedSof_overrideEncoder);
  assign when_usbphy_l602 = (Rx_Suspend && (ports_0_filter_io_filtred_se0 || ((! ports_0_filter_io_filtred_se0) && ((! ports_0_filter_io_filtred_d) ^ ports_0_portLowSpeed))));
  assign when_usbphy_l610 = (io_ctrl_ports_0_resume_valid || ((! Rx_Suspend) && ((! ports_0_filter_io_filtred_se0) && ((! ports_0_filter_io_filtred_d) ^ ports_0_portLowSpeed))));
  assign when_usbphy_l612 = (Rx_Suspend && (ports_0_filter_io_filtred_se0 || ((! ports_0_filter_io_filtred_se0) && ((! ports_0_filter_io_filtred_d) ^ ports_0_portLowSpeed))));
  assign when_usbphy_l653 = ((! ports_0_filter_io_filtred_se0) && ((! ports_0_filter_io_filtred_d) ^ ports_0_portLowSpeed));
  assign when_usbphy_l663 = ((! ports_0_filter_io_filtred_se0) && ((! ports_0_filter_io_filtred_d) ^ ports_0_portLowSpeed));
  assign when_StateMachine_l253_2 = ((! (ports_0_fsm_stateReg == ports_0_fsm_enumDef_DISCONNECTED)) && (ports_0_fsm_stateNext == ports_0_fsm_enumDef_DISCONNECTED));
  assign when_StateMachine_l253_3 = ((! (ports_0_fsm_stateReg == ports_0_fsm_enumDef_RESETTING)) && (ports_0_fsm_stateNext == ports_0_fsm_enumDef_RESETTING));
  assign when_StateMachine_l253_4 = ((! (ports_0_fsm_stateReg == ports_0_fsm_enumDef_RESETTING_DELAY)) && (ports_0_fsm_stateNext == ports_0_fsm_enumDef_RESETTING_DELAY));
  assign when_StateMachine_l253_5 = ((! (ports_0_fsm_stateReg == ports_0_fsm_enumDef_RESUMING)) && (ports_0_fsm_stateNext == ports_0_fsm_enumDef_RESUMING));
  assign when_StateMachine_l253_6 = ((! (ports_0_fsm_stateReg == ports_0_fsm_enumDef_SEND_EOP_0)) && (ports_0_fsm_stateNext == ports_0_fsm_enumDef_SEND_EOP_0));
  assign when_StateMachine_l253_7 = ((! (ports_0_fsm_stateReg == ports_0_fsm_enumDef_SEND_EOP_1)) && (ports_0_fsm_stateNext == ports_0_fsm_enumDef_SEND_EOP_1));
  assign when_StateMachine_l253_8 = ((! (ports_0_fsm_stateReg == ports_0_fsm_enumDef_RESTART_S)) && (ports_0_fsm_stateNext == ports_0_fsm_enumDef_RESTART_S));
  assign when_StateMachine_l253_9 = ((! (ports_0_fsm_stateReg == ports_0_fsm_enumDef_RESTART_E)) && (ports_0_fsm_stateNext == ports_0_fsm_enumDef_RESTART_E));
  assign when_usbphy_l512 = ((! io_ctrl_ports_0_power) || io_ctrl_usbReset);
  assign when_usbphy_l519 = (! ports_0_fsm_resetInProgress);
  assign when_usbphy_l520 = (ports_0_filter_io_filtred_dm != ports_0_filter_io_filtred_dp);
  always @(*) begin
    ports_1_rx_packet_stateNext = ports_1_rx_packet_stateReg;
    case(ports_1_rx_packet_stateReg)
      ports_1_rx_packet_enumDef_IDLE : begin
        if(ports_1_rx_history_sync_hit) begin
          ports_1_rx_packet_stateNext = ports_1_rx_packet_enumDef_PACKET;
        end
      end
      ports_1_rx_packet_enumDef_PACKET : begin
        if(ports_1_rx_destuffer_output_valid) begin
          if(when_usbphy_l429_1) begin
            if(ports_1_rx_stuffingError) begin
              ports_1_rx_packet_stateNext = ports_1_rx_packet_enumDef_ERRORED;
            end
          end
        end
      end
      ports_1_rx_packet_enumDef_ERRORED : begin
        if(ports_1_rx_packet_errorTimeout_trigger) begin
          ports_1_rx_packet_stateNext = ports_1_rx_packet_enumDef_IDLE;
        end
      end
      default : begin
      end
    endcase
    if(ports_1_rx_eop_hit) begin
      ports_1_rx_packet_stateNext = ports_1_rx_packet_enumDef_IDLE;
    end
    if(txShared_encoder_output_valid) begin
      ports_1_rx_packet_stateNext = ports_1_rx_packet_enumDef_IDLE;
    end
    if(ports_1_rx_packet_wantStart) begin
      ports_1_rx_packet_stateNext = ports_1_rx_packet_enumDef_IDLE;
    end
    if(ports_1_rx_packet_wantKill) begin
      ports_1_rx_packet_stateNext = ports_1_rx_packet_enumDef_BOOT;
    end
  end

  assign when_usbphy_l429_1 = (ports_1_rx_packet_counter == 3'b111);
  assign when_usbphy_l451_1 = ((ports_1_rx_packet_errorTimeout_p != ports_1_filter_io_filtred_dp) || (ports_1_rx_packet_errorTimeout_n != ports_1_filter_io_filtred_dm));
  assign when_StateMachine_l253_10 = ((! (ports_1_rx_packet_stateReg == ports_1_rx_packet_enumDef_IDLE)) && (ports_1_rx_packet_stateNext == ports_1_rx_packet_enumDef_IDLE));
  assign when_StateMachine_l253_11 = ((! (ports_1_rx_packet_stateReg == ports_1_rx_packet_enumDef_ERRORED)) && (ports_1_rx_packet_stateNext == ports_1_rx_packet_enumDef_ERRORED));
  always @(*) begin
    ports_1_fsm_stateNext = ports_1_fsm_stateReg;
    case(ports_1_fsm_stateReg)
      ports_1_fsm_enumDef_POWER_OFF : begin
        if(io_ctrl_ports_1_power) begin
          ports_1_fsm_stateNext = ports_1_fsm_enumDef_DISCONNECTED;
        end
      end
      ports_1_fsm_enumDef_DISCONNECTED : begin
        if(ports_1_fsm_timer_DISCONNECTED_EOI) begin
          ports_1_fsm_stateNext = ports_1_fsm_enumDef_DISABLED;
        end
      end
      ports_1_fsm_enumDef_DISABLED : begin
      end
      ports_1_fsm_enumDef_RESETTING : begin
        if(ports_1_fsm_timer_RESET_EOI) begin
          ports_1_fsm_stateNext = ports_1_fsm_enumDef_RESETTING_DELAY;
        end
      end
      ports_1_fsm_enumDef_RESETTING_DELAY : begin
        if(ports_1_fsm_timer_RESET_DELAY) begin
          ports_1_fsm_stateNext = ports_1_fsm_enumDef_RESETTING_SYNC;
        end
      end
      ports_1_fsm_enumDef_RESETTING_SYNC : begin
        if(when_usbphy_l580_1) begin
          ports_1_fsm_stateNext = ports_1_fsm_enumDef_ENABLED;
        end
      end
      ports_1_fsm_enumDef_ENABLED : begin
        if(io_ctrl_ports_1_suspend_valid) begin
          ports_1_fsm_stateNext = ports_1_fsm_enumDef_SUSPENDED;
        end else begin
          if(when_usbphy_l602_1) begin
            ports_1_fsm_stateNext = ports_1_fsm_enumDef_RESTART_E;
          end else begin
            if(io_ctrl_usbResume) begin
              ports_1_fsm_stateNext = ports_1_fsm_enumDef_RESUMING;
            end
          end
        end
      end
      ports_1_fsm_enumDef_SUSPENDED : begin
        if(when_usbphy_l610_1) begin
          ports_1_fsm_stateNext = ports_1_fsm_enumDef_RESUMING;
        end else begin
          if(when_usbphy_l612_1) begin
            ports_1_fsm_stateNext = ports_1_fsm_enumDef_RESTART_S;
          end
        end
      end
      ports_1_fsm_enumDef_RESUMING : begin
        if(ports_1_fsm_timer_RESUME_EOI) begin
          ports_1_fsm_stateNext = ports_1_fsm_enumDef_SEND_EOP_0;
        end
      end
      ports_1_fsm_enumDef_SEND_EOP_0 : begin
        if(ports_1_fsm_timer_TWO_BIT) begin
          ports_1_fsm_stateNext = ports_1_fsm_enumDef_SEND_EOP_1;
        end
      end
      ports_1_fsm_enumDef_SEND_EOP_1 : begin
        if(ports_1_fsm_timer_ONE_BIT) begin
          ports_1_fsm_stateNext = ports_1_fsm_enumDef_ENABLED;
        end
      end
      ports_1_fsm_enumDef_RESTART_S : begin
        if(when_usbphy_l653_1) begin
          ports_1_fsm_stateNext = ports_1_fsm_enumDef_RESUMING;
        end
        if(ports_1_fsm_timer_RESTART_EOI) begin
          ports_1_fsm_stateNext = ports_1_fsm_enumDef_DISCONNECTED;
        end
      end
      ports_1_fsm_enumDef_RESTART_E : begin
        if(when_usbphy_l663_1) begin
          ports_1_fsm_stateNext = ports_1_fsm_enumDef_RESUMING;
        end
        if(ports_1_fsm_timer_RESTART_EOI) begin
          ports_1_fsm_stateNext = ports_1_fsm_enumDef_DISCONNECTED;
        end
      end
      default : begin
      end
    endcase
    if(when_usbphy_l512_1) begin
      ports_1_fsm_stateNext = ports_1_fsm_enumDef_POWER_OFF;
    end else begin
      if(ports_1_rx_disconnect_event) begin
        ports_1_fsm_stateNext = ports_1_fsm_enumDef_DISCONNECTED;
      end else begin
        if(io_ctrl_ports_1_disable_valid) begin
          ports_1_fsm_stateNext = ports_1_fsm_enumDef_DISABLED;
        end else begin
          if(io_ctrl_ports_1_reset_valid) begin
            if(when_usbphy_l519_1) begin
              if(when_usbphy_l520_1) begin
                ports_1_fsm_stateNext = ports_1_fsm_enumDef_RESETTING;
              end
            end
          end
        end
      end
    end
    if(ports_1_fsm_wantStart) begin
      ports_1_fsm_stateNext = ports_1_fsm_enumDef_POWER_OFF;
    end
    if(ports_1_fsm_wantKill) begin
      ports_1_fsm_stateNext = ports_1_fsm_enumDef_BOOT;
    end
  end

  assign when_usbphy_l540_1 = ((! ports_1_filter_io_filtred_dp) && (! ports_1_filter_io_filtred_dm));
  assign when_usbphy_l547_1 = ((! io_ctrl_ports_1_reset_valid) && (ports_1_filter_io_filtred_dm != ports_1_filter_io_filtred_dp));
  assign when_usbphy_l580_1 = (! txShared_encoder_output_valid);
  assign when_usbphy_l593_1 = (ports_1_portLowSpeed && txShared_lowSpeedSof_overrideEncoder);
  assign when_usbphy_l602_1 = (Rx_Suspend && (ports_1_filter_io_filtred_se0 || ((! ports_1_filter_io_filtred_se0) && ((! ports_1_filter_io_filtred_d) ^ ports_1_portLowSpeed))));
  assign when_usbphy_l610_1 = (io_ctrl_ports_1_resume_valid || ((! Rx_Suspend) && ((! ports_1_filter_io_filtred_se0) && ((! ports_1_filter_io_filtred_d) ^ ports_1_portLowSpeed))));
  assign when_usbphy_l612_1 = (Rx_Suspend && (ports_1_filter_io_filtred_se0 || ((! ports_1_filter_io_filtred_se0) && ((! ports_1_filter_io_filtred_d) ^ ports_1_portLowSpeed))));
  assign when_usbphy_l653_1 = ((! ports_1_filter_io_filtred_se0) && ((! ports_1_filter_io_filtred_d) ^ ports_1_portLowSpeed));
  assign when_usbphy_l663_1 = ((! ports_1_filter_io_filtred_se0) && ((! ports_1_filter_io_filtred_d) ^ ports_1_portLowSpeed));
  assign when_StateMachine_l253_12 = ((! (ports_1_fsm_stateReg == ports_1_fsm_enumDef_DISCONNECTED)) && (ports_1_fsm_stateNext == ports_1_fsm_enumDef_DISCONNECTED));
  assign when_StateMachine_l253_13 = ((! (ports_1_fsm_stateReg == ports_1_fsm_enumDef_RESETTING)) && (ports_1_fsm_stateNext == ports_1_fsm_enumDef_RESETTING));
  assign when_StateMachine_l253_14 = ((! (ports_1_fsm_stateReg == ports_1_fsm_enumDef_RESETTING_DELAY)) && (ports_1_fsm_stateNext == ports_1_fsm_enumDef_RESETTING_DELAY));
  assign when_StateMachine_l253_15 = ((! (ports_1_fsm_stateReg == ports_1_fsm_enumDef_RESUMING)) && (ports_1_fsm_stateNext == ports_1_fsm_enumDef_RESUMING));
  assign when_StateMachine_l253_16 = ((! (ports_1_fsm_stateReg == ports_1_fsm_enumDef_SEND_EOP_0)) && (ports_1_fsm_stateNext == ports_1_fsm_enumDef_SEND_EOP_0));
  assign when_StateMachine_l253_17 = ((! (ports_1_fsm_stateReg == ports_1_fsm_enumDef_SEND_EOP_1)) && (ports_1_fsm_stateNext == ports_1_fsm_enumDef_SEND_EOP_1));
  assign when_StateMachine_l253_18 = ((! (ports_1_fsm_stateReg == ports_1_fsm_enumDef_RESTART_S)) && (ports_1_fsm_stateNext == ports_1_fsm_enumDef_RESTART_S));
  assign when_StateMachine_l253_19 = ((! (ports_1_fsm_stateReg == ports_1_fsm_enumDef_RESTART_E)) && (ports_1_fsm_stateNext == ports_1_fsm_enumDef_RESTART_E));
  assign when_usbphy_l512_1 = ((! io_ctrl_ports_1_power) || io_ctrl_usbReset);
  assign when_usbphy_l519_1 = (! ports_1_fsm_resetInProgress);
  assign when_usbphy_l520_1 = (ports_1_filter_io_filtred_dm != ports_1_filter_io_filtred_dp);
  always @(posedge clk_peripheral or posedge reset_peripheral) begin
    if(reset_peripheral) begin
      tickTimer_counter_value <= 2'b00;
      txShared_rxToTxDelay_active <= 1'b0;
      txShared_lowSpeedSof_state <= 2'b00;
      txShared_lowSpeedSof_overrideEncoder <= 1'b0;
      ports_0_portLowSpeed <= 1'b0;
      ports_0_rx_eop_counter <= 7'h0;
      ports_0_rx_disconnect_counter <= 7'h0;
      ports_1_portLowSpeed <= 1'b0;
      ports_1_rx_eop_counter <= 7'h0;
      ports_1_rx_disconnect_counter <= 7'h0;
      txShared_frame_stateReg <= txShared_frame_enumDef_BOOT;
      upstreamRx_stateReg <= upstreamRx_enumDef_BOOT;
      ports_0_rx_packet_stateReg <= ports_0_rx_packet_enumDef_BOOT;
      ports_0_fsm_stateReg <= ports_0_fsm_enumDef_BOOT;
      ports_1_rx_packet_stateReg <= ports_1_rx_packet_enumDef_BOOT;
      ports_1_fsm_stateReg <= ports_1_fsm_enumDef_BOOT;
    end else begin
      tickTimer_counter_value <= tickTimer_counter_valueNext;
      if(txShared_rxToTxDelay_twoCycle) begin
        txShared_rxToTxDelay_active <= 1'b0;
      end
      if(when_usbphy_l151) begin
        txShared_lowSpeedSof_overrideEncoder <= 1'b0;
      end
      txShared_lowSpeedSof_state <= (txShared_lowSpeedSof_state + _zz_txShared_lowSpeedSof_state);
      if(when_usbphy_l153) begin
        if(when_usbphy_l154) begin
          txShared_lowSpeedSof_overrideEncoder <= 1'b1;
        end
      end else begin
        if(when_usbphy_l161) begin
          txShared_lowSpeedSof_state <= (txShared_lowSpeedSof_state + 2'b01);
        end
      end
      if(when_usbphy_l395) begin
        if(when_usbphy_l396) begin
          ports_0_rx_eop_counter <= (ports_0_rx_eop_counter + 7'h01);
        end
      end else begin
        ports_0_rx_eop_counter <= 7'h0;
      end
      ports_0_rx_disconnect_counter <= (ports_0_rx_disconnect_counter + _zz_ports_0_rx_disconnect_counter);
      if(ports_0_rx_disconnect_clear) begin
        ports_0_rx_disconnect_counter <= 7'h0;
      end
      if(when_usbphy_l395_1) begin
        if(when_usbphy_l396_1) begin
          ports_1_rx_eop_counter <= (ports_1_rx_eop_counter + 7'h01);
        end
      end else begin
        ports_1_rx_eop_counter <= 7'h0;
      end
      ports_1_rx_disconnect_counter <= (ports_1_rx_disconnect_counter + _zz_ports_1_rx_disconnect_counter);
      if(ports_1_rx_disconnect_clear) begin
        ports_1_rx_disconnect_counter <= 7'h0;
      end
      txShared_frame_stateReg <= txShared_frame_stateNext;
      upstreamRx_stateReg <= upstreamRx_stateNext;
      ports_0_rx_packet_stateReg <= ports_0_rx_packet_stateNext;
      if(ports_0_rx_eop_hit) begin
        txShared_rxToTxDelay_active <= 1'b1;
      end
      ports_0_fsm_stateReg <= ports_0_fsm_stateNext;
      case(ports_0_fsm_stateReg)
        ports_0_fsm_enumDef_POWER_OFF : begin
        end
        ports_0_fsm_enumDef_DISCONNECTED : begin
          if(when_usbphy_l547) begin
            ports_0_portLowSpeed <= (! ports_0_filter_io_filtred_d);
          end
        end
        ports_0_fsm_enumDef_DISABLED : begin
        end
        ports_0_fsm_enumDef_RESETTING : begin
        end
        ports_0_fsm_enumDef_RESETTING_DELAY : begin
        end
        ports_0_fsm_enumDef_RESETTING_SYNC : begin
        end
        ports_0_fsm_enumDef_ENABLED : begin
        end
        ports_0_fsm_enumDef_SUSPENDED : begin
        end
        ports_0_fsm_enumDef_RESUMING : begin
        end
        ports_0_fsm_enumDef_SEND_EOP_0 : begin
        end
        ports_0_fsm_enumDef_SEND_EOP_1 : begin
        end
        ports_0_fsm_enumDef_RESTART_S : begin
        end
        ports_0_fsm_enumDef_RESTART_E : begin
        end
        default : begin
        end
      endcase
      if(!when_usbphy_l512) begin
        if(!ports_0_rx_disconnect_event) begin
          if(!io_ctrl_ports_0_disable_valid) begin
            if(io_ctrl_ports_0_reset_valid) begin
              if(when_usbphy_l519) begin
                if(when_usbphy_l520) begin
                  ports_0_portLowSpeed <= (! ports_0_filter_io_filtred_d);
                end
              end
            end
          end
        end
      end
      ports_1_rx_packet_stateReg <= ports_1_rx_packet_stateNext;
      if(ports_1_rx_eop_hit) begin
        txShared_rxToTxDelay_active <= 1'b1;
      end
      ports_1_fsm_stateReg <= ports_1_fsm_stateNext;
      case(ports_1_fsm_stateReg)
        ports_1_fsm_enumDef_POWER_OFF : begin
        end
        ports_1_fsm_enumDef_DISCONNECTED : begin
          if(when_usbphy_l547_1) begin
            ports_1_portLowSpeed <= (! ports_1_filter_io_filtred_d);
          end
        end
        ports_1_fsm_enumDef_DISABLED : begin
        end
        ports_1_fsm_enumDef_RESETTING : begin
        end
        ports_1_fsm_enumDef_RESETTING_DELAY : begin
        end
        ports_1_fsm_enumDef_RESETTING_SYNC : begin
        end
        ports_1_fsm_enumDef_ENABLED : begin
        end
        ports_1_fsm_enumDef_SUSPENDED : begin
        end
        ports_1_fsm_enumDef_RESUMING : begin
        end
        ports_1_fsm_enumDef_SEND_EOP_0 : begin
        end
        ports_1_fsm_enumDef_SEND_EOP_1 : begin
        end
        ports_1_fsm_enumDef_RESTART_S : begin
        end
        ports_1_fsm_enumDef_RESTART_E : begin
        end
        default : begin
        end
      endcase
      if(!when_usbphy_l512_1) begin
        if(!ports_1_rx_disconnect_event) begin
          if(!io_ctrl_ports_1_disable_valid) begin
            if(io_ctrl_ports_1_reset_valid) begin
              if(when_usbphy_l519_1) begin
                if(when_usbphy_l520_1) begin
                  ports_1_portLowSpeed <= (! ports_1_filter_io_filtred_d);
                end
              end
            end
          end
        end
      end
    end
  end

  always @(posedge clk_peripheral) begin
    if(txShared_timer_inc) begin
      txShared_timer_counter <= (txShared_timer_counter + 10'h001);
    end
    if(txShared_timer_clear) begin
      txShared_timer_counter <= 10'h0;
    end
    if(txShared_rxToTxDelay_inc) begin
      txShared_rxToTxDelay_counter <= (txShared_rxToTxDelay_counter + 9'h001);
    end
    if(txShared_rxToTxDelay_clear) begin
      txShared_rxToTxDelay_counter <= 9'h0;
    end
    if(txShared_encoder_input_valid) begin
      if(txShared_encoder_input_data) begin
        if(txShared_timer_oneCycle) begin
          txShared_encoder_counter <= (txShared_encoder_counter + 3'b001);
          if(when_usbphy_l91) begin
            txShared_encoder_state <= (! txShared_encoder_state);
          end
          if(when_usbphy_l96) begin
            txShared_encoder_counter <= 3'b000;
          end
        end
      end else begin
        if(txShared_timer_oneCycle) begin
          txShared_encoder_counter <= 3'b000;
          txShared_encoder_state <= (! txShared_encoder_state);
        end
      end
    end
    if(when_usbphy_l110) begin
      txShared_encoder_counter <= 3'b000;
      txShared_encoder_state <= 1'b1;
    end
    if(txShared_serialiser_input_valid) begin
      if(txShared_encoder_input_ready) begin
        txShared_serialiser_bitCounter <= (txShared_serialiser_bitCounter + 3'b001);
      end
    end
    if(when_usbphy_l142) begin
      txShared_serialiser_bitCounter <= 3'b000;
    end
    txShared_encoder_output_valid_regNext <= txShared_encoder_output_valid;
    if(when_usbphy_l153) begin
      if(when_usbphy_l154) begin
        txShared_lowSpeedSof_timer <= 5'h0;
      end
    end else begin
      txShared_lowSpeedSof_timer <= (txShared_lowSpeedSof_timer + 5'h01);
    end
    if(upstreamRx_timer_inc) begin
      upstreamRx_timer_counter <= (upstreamRx_timer_counter + 20'h00001);
    end
    if(upstreamRx_timer_clear) begin
      upstreamRx_timer_counter <= 20'h0;
    end
    if(ports_0_filter_io_filtred_sample) begin
      if(when_usbphy_l347) begin
        ports_0_rx_decoder_state <= (! ports_0_rx_decoder_state);
      end
    end
    if(ports_0_rx_waitSync) begin
      ports_0_rx_decoder_state <= 1'b0;
    end
    if(ports_0_rx_decoder_output_valid) begin
      ports_0_rx_destuffer_counter <= (ports_0_rx_destuffer_counter + 3'b001);
      if(when_usbphy_l368) begin
        ports_0_rx_destuffer_counter <= 3'b000;
        if(ports_0_rx_decoder_output_payload) begin
          ports_0_rx_stuffingError <= 1'b1;
        end
      end
    end
    if(ports_0_rx_waitSync) begin
      ports_0_rx_destuffer_counter <= 3'b000;
    end
    if(ports_0_rx_history_updated) begin
      _zz_ports_0_rx_history_value_1 <= _zz_ports_0_rx_history_value;
    end
    if(ports_0_rx_history_updated) begin
      _zz_ports_0_rx_history_value_2 <= _zz_ports_0_rx_history_value_1;
    end
    if(ports_0_rx_history_updated) begin
      _zz_ports_0_rx_history_value_3 <= _zz_ports_0_rx_history_value_2;
    end
    if(ports_0_rx_history_updated) begin
      _zz_ports_0_rx_history_value_4 <= _zz_ports_0_rx_history_value_3;
    end
    if(ports_0_rx_history_updated) begin
      _zz_ports_0_rx_history_value_5 <= _zz_ports_0_rx_history_value_4;
    end
    if(ports_0_rx_history_updated) begin
      _zz_ports_0_rx_history_value_6 <= _zz_ports_0_rx_history_value_5;
    end
    if(ports_0_rx_history_updated) begin
      _zz_ports_0_rx_history_value_7 <= _zz_ports_0_rx_history_value_6;
    end
    if(ports_0_rx_packet_errorTimeout_inc) begin
      ports_0_rx_packet_errorTimeout_counter <= (ports_0_rx_packet_errorTimeout_counter + 12'h001);
    end
    if(ports_0_rx_packet_errorTimeout_clear) begin
      ports_0_rx_packet_errorTimeout_counter <= 12'h0;
    end
    ports_0_rx_disconnect_hitLast <= ports_0_rx_disconnect_hit;
    if(ports_0_fsm_timer_inc) begin
      ports_0_fsm_timer_counter <= (ports_0_fsm_timer_counter + 24'h000001);
    end
    if(ports_0_fsm_timer_clear) begin
      ports_0_fsm_timer_counter <= 24'h0;
    end
    if(ports_1_filter_io_filtred_sample) begin
      if(when_usbphy_l347_1) begin
        ports_1_rx_decoder_state <= (! ports_1_rx_decoder_state);
      end
    end
    if(ports_1_rx_waitSync) begin
      ports_1_rx_decoder_state <= 1'b0;
    end
    if(ports_1_rx_decoder_output_valid) begin
      ports_1_rx_destuffer_counter <= (ports_1_rx_destuffer_counter + 3'b001);
      if(when_usbphy_l368_1) begin
        ports_1_rx_destuffer_counter <= 3'b000;
        if(ports_1_rx_decoder_output_payload) begin
          ports_1_rx_stuffingError <= 1'b1;
        end
      end
    end
    if(ports_1_rx_waitSync) begin
      ports_1_rx_destuffer_counter <= 3'b000;
    end
    if(ports_1_rx_history_updated) begin
      _zz_ports_1_rx_history_value_1 <= _zz_ports_1_rx_history_value;
    end
    if(ports_1_rx_history_updated) begin
      _zz_ports_1_rx_history_value_2 <= _zz_ports_1_rx_history_value_1;
    end
    if(ports_1_rx_history_updated) begin
      _zz_ports_1_rx_history_value_3 <= _zz_ports_1_rx_history_value_2;
    end
    if(ports_1_rx_history_updated) begin
      _zz_ports_1_rx_history_value_4 <= _zz_ports_1_rx_history_value_3;
    end
    if(ports_1_rx_history_updated) begin
      _zz_ports_1_rx_history_value_5 <= _zz_ports_1_rx_history_value_4;
    end
    if(ports_1_rx_history_updated) begin
      _zz_ports_1_rx_history_value_6 <= _zz_ports_1_rx_history_value_5;
    end
    if(ports_1_rx_history_updated) begin
      _zz_ports_1_rx_history_value_7 <= _zz_ports_1_rx_history_value_6;
    end
    if(ports_1_rx_packet_errorTimeout_inc) begin
      ports_1_rx_packet_errorTimeout_counter <= (ports_1_rx_packet_errorTimeout_counter + 12'h001);
    end
    if(ports_1_rx_packet_errorTimeout_clear) begin
      ports_1_rx_packet_errorTimeout_counter <= 12'h0;
    end
    ports_1_rx_disconnect_hitLast <= ports_1_rx_disconnect_hit;
    if(ports_1_fsm_timer_inc) begin
      ports_1_fsm_timer_counter <= (ports_1_fsm_timer_counter + 24'h000001);
    end
    if(ports_1_fsm_timer_clear) begin
      ports_1_fsm_timer_counter <= 24'h0;
    end
    case(txShared_frame_stateReg)
      txShared_frame_enumDef_IDLE : begin
        txShared_frame_wasLowSpeed <= io_ctrl_lowSpeed;
      end
      txShared_frame_enumDef_TAKE_LINE : begin
      end
      txShared_frame_enumDef_PREAMBLE_SYNC : begin
      end
      txShared_frame_enumDef_PREAMBLE_PID : begin
      end
      txShared_frame_enumDef_PREAMBLE_DELAY : begin
      end
      txShared_frame_enumDef_SYNC : begin
      end
      txShared_frame_enumDef_DATA : begin
      end
      txShared_frame_enumDef_EOP_0 : begin
      end
      txShared_frame_enumDef_EOP_1 : begin
      end
      txShared_frame_enumDef_EOP_2 : begin
      end
      default : begin
      end
    endcase
    case(ports_0_rx_packet_stateReg)
      ports_0_rx_packet_enumDef_IDLE : begin
        ports_0_rx_packet_counter <= 3'b000;
        ports_0_rx_stuffingError <= 1'b0;
      end
      ports_0_rx_packet_enumDef_PACKET : begin
        if(ports_0_rx_destuffer_output_valid) begin
          ports_0_rx_packet_counter <= (ports_0_rx_packet_counter + 3'b001);
        end
      end
      ports_0_rx_packet_enumDef_ERRORED : begin
        ports_0_rx_packet_errorTimeout_p <= ports_0_filter_io_filtred_dp;
        ports_0_rx_packet_errorTimeout_n <= ports_0_filter_io_filtred_dm;
      end
      default : begin
      end
    endcase
    if(ports_0_rx_eop_hit) begin
      txShared_rxToTxDelay_lowSpeed <= io_ctrl_lowSpeed;
    end
    case(ports_0_fsm_stateReg)
      ports_0_fsm_enumDef_POWER_OFF : begin
      end
      ports_0_fsm_enumDef_DISCONNECTED : begin
      end
      ports_0_fsm_enumDef_DISABLED : begin
      end
      ports_0_fsm_enumDef_RESETTING : begin
      end
      ports_0_fsm_enumDef_RESETTING_DELAY : begin
      end
      ports_0_fsm_enumDef_RESETTING_SYNC : begin
      end
      ports_0_fsm_enumDef_ENABLED : begin
      end
      ports_0_fsm_enumDef_SUSPENDED : begin
      end
      ports_0_fsm_enumDef_RESUMING : begin
        if(ports_0_fsm_timer_RESUME_EOI) begin
          ports_0_fsm_lowSpeedEop <= 1'b1;
        end
      end
      ports_0_fsm_enumDef_SEND_EOP_0 : begin
      end
      ports_0_fsm_enumDef_SEND_EOP_1 : begin
      end
      ports_0_fsm_enumDef_RESTART_S : begin
      end
      ports_0_fsm_enumDef_RESTART_E : begin
      end
      default : begin
      end
    endcase
    case(ports_1_rx_packet_stateReg)
      ports_1_rx_packet_enumDef_IDLE : begin
        ports_1_rx_packet_counter <= 3'b000;
        ports_1_rx_stuffingError <= 1'b0;
      end
      ports_1_rx_packet_enumDef_PACKET : begin
        if(ports_1_rx_destuffer_output_valid) begin
          ports_1_rx_packet_counter <= (ports_1_rx_packet_counter + 3'b001);
        end
      end
      ports_1_rx_packet_enumDef_ERRORED : begin
        ports_1_rx_packet_errorTimeout_p <= ports_1_filter_io_filtred_dp;
        ports_1_rx_packet_errorTimeout_n <= ports_1_filter_io_filtred_dm;
      end
      default : begin
      end
    endcase
    if(ports_1_rx_eop_hit) begin
      txShared_rxToTxDelay_lowSpeed <= io_ctrl_lowSpeed;
    end
    case(ports_1_fsm_stateReg)
      ports_1_fsm_enumDef_POWER_OFF : begin
      end
      ports_1_fsm_enumDef_DISCONNECTED : begin
      end
      ports_1_fsm_enumDef_DISABLED : begin
      end
      ports_1_fsm_enumDef_RESETTING : begin
      end
      ports_1_fsm_enumDef_RESETTING_DELAY : begin
      end
      ports_1_fsm_enumDef_RESETTING_SYNC : begin
      end
      ports_1_fsm_enumDef_ENABLED : begin
      end
      ports_1_fsm_enumDef_SUSPENDED : begin
      end
      ports_1_fsm_enumDef_RESUMING : begin
        if(ports_1_fsm_timer_RESUME_EOI) begin
          ports_1_fsm_lowSpeedEop <= 1'b1;
        end
      end
      ports_1_fsm_enumDef_SEND_EOP_0 : begin
      end
      ports_1_fsm_enumDef_SEND_EOP_1 : begin
      end
      ports_1_fsm_enumDef_RESTART_S : begin
      end
      ports_1_fsm_enumDef_RESTART_E : begin
      end
      default : begin
      end
    endcase
  end

  always @(posedge clk_peripheral or posedge reset_peripheral) begin
    if(reset_peripheral) begin
      io_ctrl_tx_payload_first <= 1'b1;
    end else begin
      if(io_ctrl_tx_fire) begin
        io_ctrl_tx_payload_first <= io_ctrl_tx_payload_last;
      end
    end
  end


endmodule

module UsbOhci (
  input  wire          io_ctrl_cmd_valid,
  output wire          io_ctrl_cmd_ready,
  input  wire          io_ctrl_cmd_payload_last,
  input  wire [0:0]    io_ctrl_cmd_payload_fragment_opcode,
  input  wire [11:0]   io_ctrl_cmd_payload_fragment_address,
  input  wire [1:0]    io_ctrl_cmd_payload_fragment_length,
  input  wire [31:0]   io_ctrl_cmd_payload_fragment_data,
  input  wire [3:0]    io_ctrl_cmd_payload_fragment_mask,
  output wire          io_ctrl_rsp_valid,
  input  wire          io_ctrl_rsp_ready,
  output wire          io_ctrl_rsp_payload_last,
  output wire [0:0]    io_ctrl_rsp_payload_fragment_opcode,
  output wire [31:0]   io_ctrl_rsp_payload_fragment_data,
  output reg           io_phy_lowSpeed,
  output reg           io_phy_tx_valid,
  input  wire          io_phy_tx_ready,
  output reg           io_phy_tx_payload_last,
  output reg  [7:0]    io_phy_tx_payload_fragment,
  input  wire          io_phy_txEop,
  input  wire          io_phy_rx_flow_valid,
  input  wire          io_phy_rx_flow_payload_stuffingError,
  input  wire [7:0]    io_phy_rx_flow_payload_data,
  input  wire          io_phy_rx_active,
  output wire          io_phy_usbReset,
  output wire          io_phy_usbResume,
  input  wire          io_phy_overcurrent,
  input  wire          io_phy_tick,
  output wire          io_phy_ports_0_disable_valid,
  input  wire          io_phy_ports_0_disable_ready,
  output wire          io_phy_ports_0_removable,
  output wire          io_phy_ports_0_power,
  output wire          io_phy_ports_0_reset_valid,
  input  wire          io_phy_ports_0_reset_ready,
  output wire          io_phy_ports_0_suspend_valid,
  input  wire          io_phy_ports_0_suspend_ready,
  output wire          io_phy_ports_0_resume_valid,
  input  wire          io_phy_ports_0_resume_ready,
  input  wire          io_phy_ports_0_connect,
  input  wire          io_phy_ports_0_disconnect,
  input  wire          io_phy_ports_0_overcurrent,
  input  wire          io_phy_ports_0_remoteResume,
  input  wire          io_phy_ports_0_lowSpeed,
  output wire          io_phy_ports_1_disable_valid,
  input  wire          io_phy_ports_1_disable_ready,
  output wire          io_phy_ports_1_removable,
  output wire          io_phy_ports_1_power,
  output wire          io_phy_ports_1_reset_valid,
  input  wire          io_phy_ports_1_reset_ready,
  output wire          io_phy_ports_1_suspend_valid,
  input  wire          io_phy_ports_1_suspend_ready,
  output wire          io_phy_ports_1_resume_valid,
  input  wire          io_phy_ports_1_resume_ready,
  input  wire          io_phy_ports_1_connect,
  input  wire          io_phy_ports_1_disconnect,
  input  wire          io_phy_ports_1_overcurrent,
  input  wire          io_phy_ports_1_remoteResume,
  input  wire          io_phy_ports_1_lowSpeed,
  output wire          io_dma_cmd_valid,
  input  wire          io_dma_cmd_ready,
  output wire          io_dma_cmd_payload_last,
  output wire [0:0]    io_dma_cmd_payload_fragment_opcode,
  output wire [31:0]   io_dma_cmd_payload_fragment_address,
  output wire [5:0]    io_dma_cmd_payload_fragment_length,
  output wire [31:0]   io_dma_cmd_payload_fragment_data,
  output wire [3:0]    io_dma_cmd_payload_fragment_mask,
  input  wire          io_dma_rsp_valid,
  output wire          io_dma_rsp_ready,
  input  wire          io_dma_rsp_payload_last,
  input  wire [0:0]    io_dma_rsp_payload_fragment_opcode,
  input  wire [31:0]   io_dma_rsp_payload_fragment_data,
  output wire          io_interrupt,
  output wire          io_interruptBios,
  input  wire          clk_peripheral,
  input  wire          reset_peripheral
);
  localparam MainState_RESET = 2'd0;
  localparam MainState_RESUME = 2'd1;
  localparam MainState_OPERATIONAL = 2'd2;
  localparam MainState_SUSPEND = 2'd3;
  localparam FlowType_BULK = 2'd0;
  localparam FlowType_CONTROL = 2'd1;
  localparam FlowType_PERIODIC = 2'd2;
  localparam endpoint_Status_OK = 1'd0;
  localparam endpoint_Status_FRAME_TIME = 1'd1;
  localparam endpoint_enumDef_BOOT = 5'd0;
  localparam endpoint_enumDef_ED_READ_CMD = 5'd1;
  localparam endpoint_enumDef_ED_READ_RSP = 5'd2;
  localparam endpoint_enumDef_ED_ANALYSE = 5'd3;
  localparam endpoint_enumDef_TD_READ_CMD = 5'd4;
  localparam endpoint_enumDef_TD_READ_RSP = 5'd5;
  localparam endpoint_enumDef_TD_READ_DELAY = 5'd6;
  localparam endpoint_enumDef_TD_ANALYSE = 5'd7;
  localparam endpoint_enumDef_TD_CHECK_TIME = 5'd8;
  localparam endpoint_enumDef_BUFFER_READ = 5'd9;
  localparam endpoint_enumDef_TOKEN = 5'd10;
  localparam endpoint_enumDef_DATA_TX = 5'd11;
  localparam endpoint_enumDef_DATA_RX = 5'd12;
  localparam endpoint_enumDef_DATA_RX_VALIDATE = 5'd13;
  localparam endpoint_enumDef_ACK_RX = 5'd14;
  localparam endpoint_enumDef_ACK_TX_0 = 5'd15;
  localparam endpoint_enumDef_ACK_TX_1 = 5'd16;
  localparam endpoint_enumDef_ACK_TX_EOP = 5'd17;
  localparam endpoint_enumDef_DATA_RX_WAIT_DMA = 5'd18;
  localparam endpoint_enumDef_UPDATE_TD_PROCESS = 5'd19;
  localparam endpoint_enumDef_UPDATE_TD_CMD = 5'd20;
  localparam endpoint_enumDef_UPDATE_ED_CMD = 5'd21;
  localparam endpoint_enumDef_UPDATE_SYNC = 5'd22;
  localparam endpoint_enumDef_ABORD = 5'd23;
  localparam endpoint_dmaLogic_enumDef_BOOT = 3'd0;
  localparam endpoint_dmaLogic_enumDef_INIT = 3'd1;
  localparam endpoint_dmaLogic_enumDef_TO_USB = 3'd2;
  localparam endpoint_dmaLogic_enumDef_FROM_USB = 3'd3;
  localparam endpoint_dmaLogic_enumDef_VALIDATION = 3'd4;
  localparam endpoint_dmaLogic_enumDef_CALC_CMD = 3'd5;
  localparam endpoint_dmaLogic_enumDef_READ_CMD = 3'd6;
  localparam endpoint_dmaLogic_enumDef_WRITE_CMD = 3'd7;
  localparam token_enumDef_BOOT = 3'd0;
  localparam token_enumDef_INIT = 3'd1;
  localparam token_enumDef_PID = 3'd2;
  localparam token_enumDef_B1 = 3'd3;
  localparam token_enumDef_B2 = 3'd4;
  localparam token_enumDef_EOP = 3'd5;
  localparam dataTx_enumDef_BOOT = 3'd0;
  localparam dataTx_enumDef_PID = 3'd1;
  localparam dataTx_enumDef_DATA = 3'd2;
  localparam dataTx_enumDef_CRC_0 = 3'd3;
  localparam dataTx_enumDef_CRC_1 = 3'd4;
  localparam dataTx_enumDef_EOP = 3'd5;
  localparam dataRx_enumDef_BOOT = 2'd0;
  localparam dataRx_enumDef_IDLE = 2'd1;
  localparam dataRx_enumDef_PID = 2'd2;
  localparam dataRx_enumDef_DATA = 2'd3;
  localparam sof_enumDef_BOOT = 2'd0;
  localparam sof_enumDef_FRAME_TX = 2'd1;
  localparam sof_enumDef_FRAME_NUMBER_CMD = 2'd2;
  localparam sof_enumDef_FRAME_NUMBER_RSP = 2'd3;
  localparam operational_enumDef_BOOT = 3'd0;
  localparam operational_enumDef_SOF = 3'd1;
  localparam operational_enumDef_ARBITER = 3'd2;
  localparam operational_enumDef_END_POINT = 3'd3;
  localparam operational_enumDef_PERIODIC_HEAD_CMD = 3'd4;
  localparam operational_enumDef_PERIODIC_HEAD_RSP = 3'd5;
  localparam operational_enumDef_WAIT_SOF = 3'd6;
  localparam hc_enumDef_BOOT = 3'd0;
  localparam hc_enumDef_RESET = 3'd1;
  localparam hc_enumDef_RESUME = 3'd2;
  localparam hc_enumDef_OPERATIONAL = 3'd3;
  localparam hc_enumDef_SUSPEND = 3'd4;
  localparam hc_enumDef_ANY_TO_RESET = 3'd5;
  localparam hc_enumDef_ANY_TO_SUSPEND = 3'd6;

  reg                 token_crc5_io_flush;
  reg                 token_crc5_io_input_valid;
  reg                 dataTx_crc16_io_flush;
  reg                 dataRx_crc16_io_flush;
  reg                 dataRx_crc16_io_input_valid;
  reg        [31:0]   endpoint_dmaLogic_storage_ram_spinal_port0;
  wire       [4:0]    token_crc5_io_result;
  wire       [4:0]    token_crc5_io_resultNext;
  wire       [15:0]   dataTx_crc16_io_result;
  wire       [15:0]   dataTx_crc16_io_resultNext;
  wire       [15:0]   dataRx_crc16_io_result;
  wire       [15:0]   dataRx_crc16_io_resultNext;
  wire       [3:0]    _zz_dmaCtx_pendingCounter;
  wire       [3:0]    _zz_dmaCtx_pendingCounter_1;
  wire       [0:0]    _zz_dmaCtx_pendingCounter_2;
  wire       [3:0]    _zz_dmaCtx_pendingCounter_3;
  wire       [0:0]    _zz_dmaCtx_pendingCounter_4;
  wire       [0:0]    _zz_reg_hcCommandStatus_startSoftReset;
  wire       [0:0]    _zz_reg_hcCommandStatus_CLF;
  wire       [0:0]    _zz_reg_hcCommandStatus_BLF;
  wire       [0:0]    _zz_reg_hcCommandStatus_OCR;
  wire       [0:0]    _zz_reg_hcInterrupt_MIE;
  wire       [0:0]    _zz_reg_hcInterrupt_MIE_1;
  wire       [0:0]    _zz_reg_hcInterrupt_SO_status;
  wire       [0:0]    _zz_reg_hcInterrupt_SO_enable;
  wire       [0:0]    _zz_reg_hcInterrupt_SO_enable_1;
  wire       [0:0]    _zz_reg_hcInterrupt_WDH_status;
  wire       [0:0]    _zz_reg_hcInterrupt_WDH_enable;
  wire       [0:0]    _zz_reg_hcInterrupt_WDH_enable_1;
  wire       [0:0]    _zz_reg_hcInterrupt_SF_status;
  wire       [0:0]    _zz_reg_hcInterrupt_SF_enable;
  wire       [0:0]    _zz_reg_hcInterrupt_SF_enable_1;
  wire       [0:0]    _zz_reg_hcInterrupt_RD_status;
  wire       [0:0]    _zz_reg_hcInterrupt_RD_enable;
  wire       [0:0]    _zz_reg_hcInterrupt_RD_enable_1;
  wire       [0:0]    _zz_reg_hcInterrupt_UE_status;
  wire       [0:0]    _zz_reg_hcInterrupt_UE_enable;
  wire       [0:0]    _zz_reg_hcInterrupt_UE_enable_1;
  wire       [0:0]    _zz_reg_hcInterrupt_FNO_status;
  wire       [0:0]    _zz_reg_hcInterrupt_FNO_enable;
  wire       [0:0]    _zz_reg_hcInterrupt_FNO_enable_1;
  wire       [0:0]    _zz_reg_hcInterrupt_RHSC_status;
  wire       [0:0]    _zz_reg_hcInterrupt_RHSC_enable;
  wire       [0:0]    _zz_reg_hcInterrupt_RHSC_enable_1;
  wire       [0:0]    _zz_reg_hcInterrupt_OC_status;
  wire       [0:0]    _zz_reg_hcInterrupt_OC_enable;
  wire       [0:0]    _zz_reg_hcInterrupt_OC_enable_1;
  wire       [13:0]   _zz_reg_hcLSThreshold_hit;
  wire       [0:0]    _zz_reg_hcRhStatus_CCIC;
  wire       [0:0]    _zz_reg_hcRhStatus_clearGlobalPower;
  wire       [0:0]    _zz_reg_hcRhStatus_setRemoteWakeupEnable;
  wire       [0:0]    _zz_reg_hcRhStatus_setGlobalPower;
  wire       [0:0]    _zz_reg_hcRhStatus_clearRemoteWakeupEnable;
  wire       [0:0]    _zz_reg_hcRhPortStatus_0_clearPortEnable;
  wire       [0:0]    _zz_reg_hcRhPortStatus_0_setPortEnable;
  wire       [0:0]    _zz_reg_hcRhPortStatus_0_setPortSuspend;
  wire       [0:0]    _zz_reg_hcRhPortStatus_0_clearSuspendStatus;
  wire       [0:0]    _zz_reg_hcRhPortStatus_0_setPortReset;
  wire       [0:0]    _zz_reg_hcRhPortStatus_0_setPortPower;
  wire       [0:0]    _zz_reg_hcRhPortStatus_0_clearPortPower;
  wire       [0:0]    _zz_reg_hcRhPortStatus_0_CSC_clear;
  wire       [0:0]    _zz_reg_hcRhPortStatus_0_PESC_clear;
  wire       [0:0]    _zz_reg_hcRhPortStatus_0_PSSC_clear;
  wire       [0:0]    _zz_reg_hcRhPortStatus_0_OCIC_clear;
  wire       [0:0]    _zz_reg_hcRhPortStatus_0_PRSC_clear;
  wire       [0:0]    _zz_reg_hcRhPortStatus_1_clearPortEnable;
  wire       [0:0]    _zz_reg_hcRhPortStatus_1_setPortEnable;
  wire       [0:0]    _zz_reg_hcRhPortStatus_1_setPortSuspend;
  wire       [0:0]    _zz_reg_hcRhPortStatus_1_clearSuspendStatus;
  wire       [0:0]    _zz_reg_hcRhPortStatus_1_setPortReset;
  wire       [0:0]    _zz_reg_hcRhPortStatus_1_setPortPower;
  wire       [0:0]    _zz_reg_hcRhPortStatus_1_clearPortPower;
  wire       [0:0]    _zz_reg_hcRhPortStatus_1_CSC_clear;
  wire       [0:0]    _zz_reg_hcRhPortStatus_1_PESC_clear;
  wire       [0:0]    _zz_reg_hcRhPortStatus_1_PSSC_clear;
  wire       [0:0]    _zz_reg_hcRhPortStatus_1_OCIC_clear;
  wire       [0:0]    _zz_reg_hcRhPortStatus_1_PRSC_clear;
  wire       [7:0]    _zz_rxTimer_ackTx;
  wire       [3:0]    _zz_rxTimer_ackTx_1;
  wire       [15:0]   _zz_endpoint_TD_isoOverrun;
  wire       [12:0]   _zz_endpoint_TD_firstOffset;
  wire       [11:0]   _zz_endpoint_TD_firstOffset_1;
  wire       [12:0]   _zz_endpoint_TD_lastOffset;
  wire       [12:0]   _zz_endpoint_TD_lastOffset_1;
  wire       [0:0]    _zz_endpoint_TD_lastOffset_2;
  wire       [25:0]   _zz_endpoint_currentAddressBmb;
  wire       [13:0]   _zz_endpoint_transactionSizeMinusOne;
  wire       [13:0]   _zz_endpoint_dataDone;
  wire       [2:0]    _zz_endpoint_dmaLogic_storage_full_1;
  wire       [7:0]    _zz_endpoint_dmaLogic_storage_full_2;
  wire       [5:0]    _zz_endpoint_dmaLogic_lengthMax;
  wire       [13:0]   _zz_endpoint_dmaLogic_lengthCalc;
  wire       [13:0]   _zz_endpoint_dmaLogic_lengthCalc_1;
  wire       [13:0]   _zz_endpoint_dmaLogic_lengthCalc_2;
  wire       [6:0]    _zz_endpoint_dmaLogic_beatCount;
  wire       [6:0]    _zz_endpoint_dmaLogic_beatCount_1;
  wire       [1:0]    _zz_endpoint_dmaLogic_beatCount_2;
  wire       [6:0]    _zz_endpoint_dmaLogic_fromUsb_dmaReady;
  wire       [13:0]   _zz_when_UsbOhci_l1011;
  wire       [13:0]   _zz_endpoint_dmaLogic_overflow;
  wire       [12:0]   _zz_endpoint_lastAddress_1;
  wire       [12:0]   _zz_endpoint_lastAddress_2;
  wire       [10:0]   _zz_endpoint_dmaLogic_fromUsbCounter;
  wire       [0:0]    _zz_endpoint_dmaLogic_fromUsbCounter_1;
  wire       [13:0]   _zz_endpoint_dmaLogic_lastMask;
  wire       [13:0]   _zz_endpoint_dmaLogic_lastMask_1;
  wire       [13:0]   _zz_endpoint_dmaLogic_lastMask_2;
  wire       [13:0]   _zz_endpoint_dmaLogic_lastMask_3;
  wire       [13:0]   _zz_endpoint_dmaLogic_lastMask_4;
  wire       [13:0]   _zz_endpoint_dmaLogic_lastMask_5;
  wire       [13:0]   _zz_endpoint_dmaLogic_lastMask_6;
  wire       [13:0]   _zz_endpoint_dmaLogic_lastMask_7;
  wire       [3:0]    _zz_endpoint_dmaLogic_headHit;
  wire       [11:0]   _zz_endpoint_dmaLogic_headHit_1;
  wire       [3:0]    _zz_endpoint_dmaLogic_lastHit;
  wire       [11:0]   _zz_endpoint_dmaLogic_lastHit_1;
  wire       [13:0]   _zz_endpoint_dmaLogic_lastHit_2;
  wire       [13:0]   _zz_endpoint_dmaLogic_lastHit_3;
  wire       [13:0]   _zz_endpoint_byteCountCalc;
  wire       [13:0]   _zz_endpoint_byteCountCalc_1;
  wire       [16:0]   _zz_endpoint_fsTimeCheck;
  wire       [16:0]   _zz_endpoint_fsTimeCheck_1;
  wire       [15:0]   _zz_token_data;
  wire       [4:0]    _zz_ioDma_cmd_payload_fragment_length;
  wire       [13:0]   _zz__zz_endpoint_lastAddress;
  wire       [13:0]   _zz__zz_endpoint_lastAddress_1;
  wire       [11:0]   _zz__zz_endpoint_lastAddress_2;
  wire       [13:0]   _zz_endpoint_lastAddress_3;
  wire       [13:0]   _zz_endpoint_lastAddress_4;
  wire       [13:0]   _zz_endpoint_lastAddress_5;
  wire       [13:0]   _zz_endpoint_lastAddress_6;
  wire       [13:0]   _zz_when_UsbOhci_l1386;
  wire       [1:0]    _zz_endpoint_TD_words_0;
  wire       [4:0]    _zz_ioDma_cmd_payload_fragment_length_1;
  wire       [3:0]    _zz_ioDma_cmd_payload_last;
  wire       [2:0]    _zz_ioDma_cmd_payload_last_1;
  wire       [11:0]   _zz__zz_ioDma_cmd_payload_fragment_data;
  wire       [13:0]   _zz__zz_ioDma_cmd_payload_fragment_data_1;
  wire       [13:0]   _zz__zz_ioDma_cmd_payload_fragment_data_2;
  wire       [13:0]   _zz__zz_ioDma_cmd_payload_fragment_data_3;
  wire       [11:0]   _zz_endpoint_dmaLogic_storage_writePtr;
  wire       [11:0]   _zz_endpoint_dmaLogic_storage_readPtr;
  wire       [13:0]   _zz_endpoint_dmaLogic_storage_readPtr_1;
  wire       [7:0]    _zz_endpoint_dmaLogic_storage_readPtr_2;
  wire       [11:0]   _zz_endpoint_dmaLogic_storage_writePtr_1;
  wire       [13:0]   _zz_endpoint_dmaLogic_storage_writePtr_2;
  wire       [7:0]    _zz_endpoint_dmaLogic_storage_writePtr_3;
  wire       [11:0]   _zz_endpoint_dmaLogic_storage_readPtr_3;
  wire       [13:0]   _zz_endpoint_dmaLogic_fromUsb_transactionSizeMax;
  wire       [13:0]   _zz_endpoint_dmaLogic_fromUsb_transactionSizeMax_1;
  wire       [13:0]   _zz_endpoint_currentAddress;
  wire       [13:0]   _zz_endpoint_currentAddress_1;
  wire       [13:0]   _zz_endpoint_currentAddress_2;
  wire       [13:0]   _zz_endpoint_currentAddress_3;
  reg        [7:0]    _zz_dataTx_data_payload_fragment;
  wire       [31:0]   _zz_ioDma_cmd_payload_fragment_address;
  wire       [6:0]    _zz_ioDma_cmd_payload_fragment_address_1;
  reg                 _zz_1;
  reg                 unscheduleAll_valid;
  reg                 unscheduleAll_ready;
  reg                 ioDma_cmd_valid;
  wire                ioDma_cmd_ready;
  reg                 ioDma_cmd_payload_last;
  reg        [0:0]    ioDma_cmd_payload_fragment_opcode;
  reg        [31:0]   ioDma_cmd_payload_fragment_address;
  reg        [5:0]    ioDma_cmd_payload_fragment_length;
  reg        [31:0]   ioDma_cmd_payload_fragment_data;
  reg        [3:0]    ioDma_cmd_payload_fragment_mask;
  wire                ioDma_rsp_valid;
  wire                ioDma_rsp_ready;
  wire                ioDma_rsp_payload_last;
  wire       [0:0]    ioDma_rsp_payload_fragment_opcode;
  wire       [31:0]   ioDma_rsp_payload_fragment_data;
  reg        [3:0]    dmaCtx_pendingCounter;
  wire                ioDma_cmd_fire;
  wire                ioDma_rsp_fire;
  wire                dmaCtx_pendingFull;
  wire                dmaCtx_pendingEmpty;
  reg        [3:0]    dmaCtx_beatCounter;
  wire                when_UsbOhci_l158;
  wire                io_dma_cmd_fire;
  reg                 io_dma_cmd_payload_first;
  wire                _zz_io_dma_cmd_valid;
  wire       [31:0]   dmaRspMux_vec_0;
  wire       [31:0]   dmaRspMux_data;
  reg        [3:0]    dmaReadCtx_counter;
  reg        [3:0]    dmaWriteCtx_counter;
  reg                 ctrlHalt;
  wire                ctrl_readErrorFlag;
  wire                ctrl_writeErrorFlag;
  wire                ctrl_readHaltTrigger;
  reg                 ctrl_writeHaltTrigger;
  wire                ctrl_rsp_valid;
  wire                ctrl_rsp_ready;
  wire                ctrl_rsp_payload_last;
  reg        [0:0]    ctrl_rsp_payload_fragment_opcode;
  reg        [31:0]   ctrl_rsp_payload_fragment_data;
  wire                _zz_ctrl_rsp_ready;
  reg                 _zz_ctrl_rsp_ready_1;
  wire                _zz_io_ctrl_rsp_valid;
  reg                 _zz_io_ctrl_rsp_valid_1;
  reg                 _zz_io_ctrl_rsp_payload_last;
  reg        [0:0]    _zz_io_ctrl_rsp_payload_fragment_opcode;
  reg        [31:0]   _zz_io_ctrl_rsp_payload_fragment_data;
  wire                when_Stream_l393;
  wire                ctrl_askWrite;
  wire                ctrl_askRead;
  wire                io_ctrl_cmd_fire;
  wire                ctrl_doWrite;
  wire                ctrl_doRead;
  wire                when_BmbSlaveFactory_l33;
  wire                when_BmbSlaveFactory_l35;
  reg                 doUnschedule;
  reg                 doSoftReset;
  wire                when_UsbOhci_l224;
  wire       [4:0]    reg_hcRevision_REV;
  reg        [1:0]    reg_hcControl_CBSR;
  reg                 reg_hcControl_PLE;
  reg                 reg_hcControl_IE;
  reg                 reg_hcControl_CLE;
  reg                 reg_hcControl_BLE;
  reg        [1:0]    reg_hcControl_HCFS;
  reg                 reg_hcControl_IR;
  reg                 reg_hcControl_RWC;
  reg                 reg_hcControl_RWE;
  reg                 reg_hcControl_HCFSWrite_valid;
  wire       [1:0]    reg_hcControl_HCFSWrite_payload;
  reg                 reg_hcCommandStatus_startSoftReset;
  reg                 when_BusSlaveFactory_l377;
  wire                when_BusSlaveFactory_l379;
  reg                 reg_hcCommandStatus_CLF;
  reg                 when_BusSlaveFactory_l377_1;
  wire                when_BusSlaveFactory_l379_1;
  reg                 reg_hcCommandStatus_BLF;
  reg                 when_BusSlaveFactory_l377_2;
  wire                when_BusSlaveFactory_l379_2;
  reg                 reg_hcCommandStatus_OCR;
  reg                 when_BusSlaveFactory_l377_3;
  wire                when_BusSlaveFactory_l379_3;
  reg        [1:0]    reg_hcCommandStatus_SOC;
  reg                 reg_hcInterrupt_unmaskedPending;
  reg                 reg_hcInterrupt_MIE;
  reg                 when_BusSlaveFactory_l377_4;
  wire                when_BusSlaveFactory_l379_4;
  reg                 when_BusSlaveFactory_l341;
  wire                when_BusSlaveFactory_l347;
  reg                 reg_hcInterrupt_SO_status;
  reg                 when_BusSlaveFactory_l341_1;
  wire                when_BusSlaveFactory_l347_1;
  reg                 reg_hcInterrupt_SO_enable;
  reg                 when_BusSlaveFactory_l377_5;
  wire                when_BusSlaveFactory_l379_5;
  reg                 when_BusSlaveFactory_l341_2;
  wire                when_BusSlaveFactory_l347_2;
  wire                when_UsbOhci_l290;
  reg                 reg_hcInterrupt_WDH_status;
  reg                 when_BusSlaveFactory_l341_3;
  wire                when_BusSlaveFactory_l347_3;
  reg                 reg_hcInterrupt_WDH_enable;
  reg                 when_BusSlaveFactory_l377_6;
  wire                when_BusSlaveFactory_l379_6;
  reg                 when_BusSlaveFactory_l341_4;
  wire                when_BusSlaveFactory_l347_4;
  wire                when_UsbOhci_l290_1;
  reg                 reg_hcInterrupt_SF_status;
  reg                 when_BusSlaveFactory_l341_5;
  wire                when_BusSlaveFactory_l347_5;
  reg                 reg_hcInterrupt_SF_enable;
  reg                 when_BusSlaveFactory_l377_7;
  wire                when_BusSlaveFactory_l379_7;
  reg                 when_BusSlaveFactory_l341_6;
  wire                when_BusSlaveFactory_l347_6;
  wire                when_UsbOhci_l290_2;
  reg                 reg_hcInterrupt_RD_status;
  reg                 when_BusSlaveFactory_l341_7;
  wire                when_BusSlaveFactory_l347_7;
  reg                 reg_hcInterrupt_RD_enable;
  reg                 when_BusSlaveFactory_l377_8;
  wire                when_BusSlaveFactory_l379_8;
  reg                 when_BusSlaveFactory_l341_8;
  wire                when_BusSlaveFactory_l347_8;
  wire                when_UsbOhci_l290_3;
  reg                 reg_hcInterrupt_UE_status;
  reg                 when_BusSlaveFactory_l341_9;
  wire                when_BusSlaveFactory_l347_9;
  reg                 reg_hcInterrupt_UE_enable;
  reg                 when_BusSlaveFactory_l377_9;
  wire                when_BusSlaveFactory_l379_9;
  reg                 when_BusSlaveFactory_l341_10;
  wire                when_BusSlaveFactory_l347_10;
  wire                when_UsbOhci_l290_4;
  reg                 reg_hcInterrupt_FNO_status;
  reg                 when_BusSlaveFactory_l341_11;
  wire                when_BusSlaveFactory_l347_11;
  reg                 reg_hcInterrupt_FNO_enable;
  reg                 when_BusSlaveFactory_l377_10;
  wire                when_BusSlaveFactory_l379_10;
  reg                 when_BusSlaveFactory_l341_12;
  wire                when_BusSlaveFactory_l347_12;
  wire                when_UsbOhci_l290_5;
  reg                 reg_hcInterrupt_RHSC_status;
  reg                 when_BusSlaveFactory_l341_13;
  wire                when_BusSlaveFactory_l347_13;
  reg                 reg_hcInterrupt_RHSC_enable;
  reg                 when_BusSlaveFactory_l377_11;
  wire                when_BusSlaveFactory_l379_11;
  reg                 when_BusSlaveFactory_l341_14;
  wire                when_BusSlaveFactory_l347_14;
  wire                when_UsbOhci_l290_6;
  reg                 reg_hcInterrupt_OC_status;
  reg                 when_BusSlaveFactory_l341_15;
  wire                when_BusSlaveFactory_l347_15;
  reg                 reg_hcInterrupt_OC_enable;
  reg                 when_BusSlaveFactory_l377_12;
  wire                when_BusSlaveFactory_l379_12;
  reg                 when_BusSlaveFactory_l341_16;
  wire                when_BusSlaveFactory_l347_16;
  wire                reg_hcInterrupt_doIrq;
  wire       [31:0]   reg_hcHCCA_HCCA_address;
  reg        [23:0]   reg_hcHCCA_HCCA_reg;
  wire       [31:0]   reg_hcPeriodCurrentED_PCED_address;
  reg        [27:0]   reg_hcPeriodCurrentED_PCED_reg;
  wire                reg_hcPeriodCurrentED_isZero;
  wire       [31:0]   reg_hcControlHeadED_CHED_address;
  reg        [27:0]   reg_hcControlHeadED_CHED_reg;
  wire       [31:0]   reg_hcControlCurrentED_CCED_address;
  reg        [27:0]   reg_hcControlCurrentED_CCED_reg;
  wire                reg_hcControlCurrentED_isZero;
  wire       [31:0]   reg_hcBulkHeadED_BHED_address;
  reg        [27:0]   reg_hcBulkHeadED_BHED_reg;
  wire       [31:0]   reg_hcBulkCurrentED_BCED_address;
  reg        [27:0]   reg_hcBulkCurrentED_BCED_reg;
  wire                reg_hcBulkCurrentED_isZero;
  wire       [31:0]   reg_hcDoneHead_DH_address;
  reg        [27:0]   reg_hcDoneHead_DH_reg;
  reg        [13:0]   reg_hcFmInterval_FI;
  reg        [14:0]   reg_hcFmInterval_FSMPS;
  reg                 reg_hcFmInterval_FIT;
  reg        [13:0]   reg_hcFmRemaining_FR;
  reg                 reg_hcFmRemaining_FRT;
  reg        [15:0]   reg_hcFmNumber_FN;
  reg                 reg_hcFmNumber_overflow;
  wire       [15:0]   reg_hcFmNumber_FNp1;
  reg        [13:0]   reg_hcPeriodicStart_PS;
  reg        [11:0]   reg_hcLSThreshold_LST;
  wire                reg_hcLSThreshold_hit;
  wire       [7:0]    reg_hcRhDescriptorA_NDP;
  reg                 reg_hcRhDescriptorA_PSM;
  reg                 reg_hcRhDescriptorA_NPS;
  reg                 reg_hcRhDescriptorA_OCPM;
  reg                 reg_hcRhDescriptorA_NOCP;
  reg        [7:0]    reg_hcRhDescriptorA_POTPGT;
  reg        [1:0]    reg_hcRhDescriptorB_DR;
  reg        [1:0]    reg_hcRhDescriptorB_PPCM;
  reg                 reg_hcRhStatus_DRWE;
  reg                 reg_hcRhStatus_CCIC;
  reg                 when_BusSlaveFactory_l341_17;
  wire                when_BusSlaveFactory_l347_17;
  reg                 io_phy_overcurrent_regNext;
  wire                when_UsbOhci_l397;
  reg                 reg_hcRhStatus_clearGlobalPower;
  reg                 when_BusSlaveFactory_l377_13;
  wire                when_BusSlaveFactory_l379_13;
  reg                 reg_hcRhStatus_setRemoteWakeupEnable;
  reg                 when_BusSlaveFactory_l377_14;
  wire                when_BusSlaveFactory_l379_14;
  reg                 reg_hcRhStatus_setGlobalPower;
  reg                 when_BusSlaveFactory_l377_15;
  wire                when_BusSlaveFactory_l379_15;
  reg                 reg_hcRhStatus_clearRemoteWakeupEnable;
  reg                 when_BusSlaveFactory_l377_16;
  wire                when_BusSlaveFactory_l379_16;
  reg                 reg_hcRhPortStatus_0_clearPortEnable;
  reg                 when_BusSlaveFactory_l377_17;
  wire                when_BusSlaveFactory_l379_17;
  reg                 reg_hcRhPortStatus_0_setPortEnable;
  reg                 when_BusSlaveFactory_l377_18;
  wire                when_BusSlaveFactory_l379_18;
  reg                 reg_hcRhPortStatus_0_setPortSuspend;
  reg                 when_BusSlaveFactory_l377_19;
  wire                when_BusSlaveFactory_l379_19;
  reg                 reg_hcRhPortStatus_0_clearSuspendStatus;
  reg                 when_BusSlaveFactory_l377_20;
  wire                when_BusSlaveFactory_l379_20;
  reg                 reg_hcRhPortStatus_0_setPortReset;
  reg                 when_BusSlaveFactory_l377_21;
  wire                when_BusSlaveFactory_l379_21;
  reg                 reg_hcRhPortStatus_0_setPortPower;
  reg                 when_BusSlaveFactory_l377_22;
  wire                when_BusSlaveFactory_l379_22;
  reg                 reg_hcRhPortStatus_0_clearPortPower;
  reg                 when_BusSlaveFactory_l377_23;
  wire                when_BusSlaveFactory_l379_23;
  reg                 reg_hcRhPortStatus_0_resume;
  reg                 reg_hcRhPortStatus_0_reset;
  reg                 reg_hcRhPortStatus_0_suspend;
  reg                 reg_hcRhPortStatus_0_connected;
  reg                 reg_hcRhPortStatus_0_PSS;
  reg                 reg_hcRhPortStatus_0_PPS;
  wire                reg_hcRhPortStatus_0_CCS;
  reg                 reg_hcRhPortStatus_0_PES;
  wire                reg_hcRhPortStatus_0_CSC_set;
  reg                 reg_hcRhPortStatus_0_CSC_clear;
  reg                 reg_hcRhPortStatus_0_CSC_reg;
  reg                 when_BusSlaveFactory_l377_24;
  wire                when_BusSlaveFactory_l379_24;
  wire                reg_hcRhPortStatus_0_PESC_set;
  reg                 reg_hcRhPortStatus_0_PESC_clear;
  reg                 reg_hcRhPortStatus_0_PESC_reg;
  reg                 when_BusSlaveFactory_l377_25;
  wire                when_BusSlaveFactory_l379_25;
  wire                reg_hcRhPortStatus_0_PSSC_set;
  reg                 reg_hcRhPortStatus_0_PSSC_clear;
  reg                 reg_hcRhPortStatus_0_PSSC_reg;
  reg                 when_BusSlaveFactory_l377_26;
  wire                when_BusSlaveFactory_l379_26;
  wire                reg_hcRhPortStatus_0_OCIC_set;
  reg                 reg_hcRhPortStatus_0_OCIC_clear;
  reg                 reg_hcRhPortStatus_0_OCIC_reg;
  reg                 when_BusSlaveFactory_l377_27;
  wire                when_BusSlaveFactory_l379_27;
  wire                reg_hcRhPortStatus_0_PRSC_set;
  reg                 reg_hcRhPortStatus_0_PRSC_clear;
  reg                 reg_hcRhPortStatus_0_PRSC_reg;
  reg                 when_BusSlaveFactory_l377_28;
  wire                when_BusSlaveFactory_l379_28;
  wire                when_UsbOhci_l448;
  wire                when_UsbOhci_l448_1;
  wire                when_UsbOhci_l448_2;
  wire                when_UsbOhci_l449;
  wire                when_UsbOhci_l449_1;
  wire                when_UsbOhci_l450;
  wire                when_UsbOhci_l451;
  wire                when_UsbOhci_l452;
  wire                when_UsbOhci_l458;
  reg                 reg_hcRhPortStatus_0_CCS_regNext;
  wire                io_phy_ports_0_suspend_fire;
  wire                io_phy_ports_0_reset_fire;
  wire                io_phy_ports_0_resume_fire;
  reg                 reg_hcRhPortStatus_1_clearPortEnable;
  reg                 when_BusSlaveFactory_l377_29;
  wire                when_BusSlaveFactory_l379_29;
  reg                 reg_hcRhPortStatus_1_setPortEnable;
  reg                 when_BusSlaveFactory_l377_30;
  wire                when_BusSlaveFactory_l379_30;
  reg                 reg_hcRhPortStatus_1_setPortSuspend;
  reg                 when_BusSlaveFactory_l377_31;
  wire                when_BusSlaveFactory_l379_31;
  reg                 reg_hcRhPortStatus_1_clearSuspendStatus;
  reg                 when_BusSlaveFactory_l377_32;
  wire                when_BusSlaveFactory_l379_32;
  reg                 reg_hcRhPortStatus_1_setPortReset;
  reg                 when_BusSlaveFactory_l377_33;
  wire                when_BusSlaveFactory_l379_33;
  reg                 reg_hcRhPortStatus_1_setPortPower;
  reg                 when_BusSlaveFactory_l377_34;
  wire                when_BusSlaveFactory_l379_34;
  reg                 reg_hcRhPortStatus_1_clearPortPower;
  reg                 when_BusSlaveFactory_l377_35;
  wire                when_BusSlaveFactory_l379_35;
  reg                 reg_hcRhPortStatus_1_resume;
  reg                 reg_hcRhPortStatus_1_reset;
  reg                 reg_hcRhPortStatus_1_suspend;
  reg                 reg_hcRhPortStatus_1_connected;
  reg                 reg_hcRhPortStatus_1_PSS;
  reg                 reg_hcRhPortStatus_1_PPS;
  wire                reg_hcRhPortStatus_1_CCS;
  reg                 reg_hcRhPortStatus_1_PES;
  wire                reg_hcRhPortStatus_1_CSC_set;
  reg                 reg_hcRhPortStatus_1_CSC_clear;
  reg                 reg_hcRhPortStatus_1_CSC_reg;
  reg                 when_BusSlaveFactory_l377_36;
  wire                when_BusSlaveFactory_l379_36;
  wire                reg_hcRhPortStatus_1_PESC_set;
  reg                 reg_hcRhPortStatus_1_PESC_clear;
  reg                 reg_hcRhPortStatus_1_PESC_reg;
  reg                 when_BusSlaveFactory_l377_37;
  wire                when_BusSlaveFactory_l379_37;
  wire                reg_hcRhPortStatus_1_PSSC_set;
  reg                 reg_hcRhPortStatus_1_PSSC_clear;
  reg                 reg_hcRhPortStatus_1_PSSC_reg;
  reg                 when_BusSlaveFactory_l377_38;
  wire                when_BusSlaveFactory_l379_38;
  wire                reg_hcRhPortStatus_1_OCIC_set;
  reg                 reg_hcRhPortStatus_1_OCIC_clear;
  reg                 reg_hcRhPortStatus_1_OCIC_reg;
  reg                 when_BusSlaveFactory_l377_39;
  wire                when_BusSlaveFactory_l379_39;
  wire                reg_hcRhPortStatus_1_PRSC_set;
  reg                 reg_hcRhPortStatus_1_PRSC_clear;
  reg                 reg_hcRhPortStatus_1_PRSC_reg;
  reg                 when_BusSlaveFactory_l377_40;
  wire                when_BusSlaveFactory_l379_40;
  wire                when_UsbOhci_l448_3;
  wire                when_UsbOhci_l448_4;
  wire                when_UsbOhci_l448_5;
  wire                when_UsbOhci_l449_2;
  wire                when_UsbOhci_l449_3;
  wire                when_UsbOhci_l450_1;
  wire                when_UsbOhci_l451_1;
  wire                when_UsbOhci_l452_1;
  wire                when_UsbOhci_l458_1;
  reg                 reg_hcRhPortStatus_1_CCS_regNext;
  wire                io_phy_ports_1_suspend_fire;
  wire                io_phy_ports_1_reset_fire;
  wire                io_phy_ports_1_resume_fire;
  reg                 frame_run;
  reg                 frame_reload;
  wire                frame_overflow;
  reg                 frame_tick;
  wire                frame_section1;
  reg        [14:0]   frame_limitCounter;
  wire                frame_limitHit;
  reg        [2:0]    frame_decrementTimer;
  wire                frame_decrementTimerOverflow;
  wire                when_UsbOhci_l514;
  wire                when_UsbOhci_l516;
  wire                when_UsbOhci_l528;
  reg                 token_wantExit;
  reg                 token_wantStart;
  reg                 token_wantKill;
  reg        [3:0]    token_pid;
  reg        [10:0]   token_data;
  reg                 dataTx_wantExit;
  reg                 dataTx_wantStart;
  reg                 dataTx_wantKill;
  reg        [3:0]    dataTx_pid;
  reg                 dataTx_data_valid;
  reg                 dataTx_data_ready;
  reg                 dataTx_data_payload_last;
  reg        [7:0]    dataTx_data_payload_fragment;
  wire                dataTx_data_fire;
  wire                rxTimer_lowSpeed;
  reg        [7:0]    rxTimer_counter;
  reg                 rxTimer_clear;
  wire                rxTimer_rxTimeout;
  wire                rxTimer_ackTx;
  wire                rxPidOk;
  wire                _zz_2;
  wire       [7:0]    _zz_dataRx_pid;
  wire                when_Misc_l87;
  reg                 dataRx_wantExit;
  reg                 dataRx_wantStart;
  reg                 dataRx_wantKill;
  reg        [3:0]    dataRx_pid;
  reg                 dataRx_data_valid;
  wire       [7:0]    dataRx_data_payload;
  wire       [7:0]    dataRx_history_0;
  wire       [7:0]    dataRx_history_1;
  reg        [7:0]    _zz_dataRx_history_0;
  reg        [7:0]    _zz_dataRx_history_1;
  reg        [1:0]    dataRx_valids;
  reg                 dataRx_notResponding;
  reg                 dataRx_stuffingError;
  reg                 dataRx_pidError;
  reg                 dataRx_crcError;
  wire                dataRx_hasError;
  reg                 sof_wantExit;
  reg                 sof_wantStart;
  reg                 sof_wantKill;
  reg                 sof_doInterruptDelay;
  reg                 priority_bulk;
  reg        [1:0]    priority_counter;
  reg                 priority_tick;
  reg                 priority_skip;
  wire                when_UsbOhci_l651;
  reg        [2:0]    interruptDelay_counter;
  reg                 interruptDelay_tick;
  wire                interruptDelay_done;
  wire                interruptDelay_disabled;
  reg                 interruptDelay_disable;
  reg                 interruptDelay_load_valid;
  reg        [2:0]    interruptDelay_load_payload;
  wire                when_UsbOhci_l673;
  wire                when_UsbOhci_l677;
  reg                 endpoint_wantExit;
  reg                 endpoint_wantStart;
  reg                 endpoint_wantKill;
  reg        [1:0]    endpoint_flowType;
  reg        [0:0]    endpoint_status_1;
  reg                 endpoint_dataPhase;
  reg        [31:0]   endpoint_ED_address;
  reg        [31:0]   endpoint_ED_words_0;
  reg        [31:0]   endpoint_ED_words_1;
  reg        [31:0]   endpoint_ED_words_2;
  reg        [31:0]   endpoint_ED_words_3;
  wire       [6:0]    endpoint_ED_FA;
  wire       [3:0]    endpoint_ED_EN;
  wire       [1:0]    endpoint_ED_D;
  wire                endpoint_ED_S;
  wire                endpoint_ED_K;
  wire                endpoint_ED_F;
  wire       [10:0]   endpoint_ED_MPS;
  wire       [27:0]   endpoint_ED_tailP;
  wire                endpoint_ED_H;
  wire                endpoint_ED_C;
  wire       [27:0]   endpoint_ED_headP;
  wire       [27:0]   endpoint_ED_nextED;
  wire                endpoint_ED_tdEmpty;
  wire                endpoint_ED_isFs;
  wire                endpoint_ED_isoOut;
  wire                when_UsbOhci_l738;
  wire       [31:0]   endpoint_TD_address;
  reg        [31:0]   endpoint_TD_words_0;
  reg        [31:0]   endpoint_TD_words_1;
  reg        [31:0]   endpoint_TD_words_2;
  reg        [31:0]   endpoint_TD_words_3;
  wire       [3:0]    endpoint_TD_CC;
  wire       [1:0]    endpoint_TD_EC;
  wire       [1:0]    endpoint_TD_T;
  wire       [2:0]    endpoint_TD_DI;
  wire       [1:0]    endpoint_TD_DP;
  wire                endpoint_TD_R;
  wire       [31:0]   endpoint_TD_CBP;
  wire       [27:0]   endpoint_TD_nextTD;
  wire       [31:0]   endpoint_TD_BE;
  wire       [2:0]    endpoint_TD_FC;
  wire       [15:0]   endpoint_TD_SF;
  wire       [15:0]   endpoint_TD_isoRelativeFrameNumber;
  wire                endpoint_TD_tooEarly;
  wire       [2:0]    endpoint_TD_isoFrameNumber;
  wire                endpoint_TD_isoOverrun;
  reg                 endpoint_TD_isoOverrunReg;
  wire                endpoint_TD_isoLast;
  reg        [12:0]   endpoint_TD_isoBase;
  reg        [12:0]   endpoint_TD_isoBaseNext;
  reg                 endpoint_TD_isoZero;
  reg                 endpoint_TD_isoLastReg;
  reg                 endpoint_TD_tooEarlyReg;
  wire                endpoint_TD_isSinglePage;
  wire       [12:0]   endpoint_TD_firstOffset;
  reg        [12:0]   endpoint_TD_lastOffset;
  wire                endpoint_TD_allowRounding;
  reg                 endpoint_TD_retire;
  reg                 endpoint_TD_upateCBP;
  reg                 endpoint_TD_noUpdate;
  reg                 endpoint_TD_dataPhaseUpdate;
  wire       [1:0]    endpoint_TD_TNext;
  wire                endpoint_TD_dataPhaseNext;
  wire       [3:0]    endpoint_TD_dataPid;
  wire       [3:0]    endpoint_TD_dataPidWrong;
  reg                 endpoint_TD_clear;
  wire       [1:0]    endpoint_tockenType;
  wire                endpoint_isIn;
  reg                 endpoint_applyNextED;
  reg        [13:0]   endpoint_currentAddress;
  wire       [31:0]   endpoint_currentAddressFull;
  wire       [31:0]   endpoint_currentAddressBmb;
  reg        [12:0]   endpoint_lastAddress;
  wire       [13:0]   endpoint_transactionSizeMinusOne;
  wire       [13:0]   endpoint_transactionSize;
  reg                 endpoint_zeroLength;
  wire                endpoint_dataDone;
  reg                 endpoint_dmaLogic_wantExit;
  reg                 endpoint_dmaLogic_wantStart;
  reg                 endpoint_dmaLogic_wantKill;
  reg                 endpoint_dmaLogic_storage_readCmd_valid;
  wire                endpoint_dmaLogic_storage_readCmd_ready;
  reg        [5:0]    endpoint_dmaLogic_storage_readCmd_payload;
  wire                endpoint_dmaLogic_storage_readRsp_valid;
  reg                 endpoint_dmaLogic_storage_readRsp_ready;
  wire       [31:0]   endpoint_dmaLogic_storage_readRsp_payload;
  reg                 _zz_endpoint_dmaLogic_storage_readRsp_valid;
  wire                endpoint_dmaLogic_storage_readCmd_fire;
  wire                endpoint_dmaLogic_storage_readRsp_isFree;
  reg                 endpoint_dmaLogic_storage_write_valid;
  reg        [5:0]    endpoint_dmaLogic_storage_write_payload_address;
  reg        [31:0]   endpoint_dmaLogic_storage_write_payload_data;
  reg        [6:0]    endpoint_dmaLogic_storage_writePtr;
  reg        [6:0]    endpoint_dmaLogic_storage_readPtr;
  wire       [2:0]    _zz_endpoint_dmaLogic_storage_full;
  wire                endpoint_dmaLogic_storage_full;
  reg                 endpoint_dmaLogic_validated;
  reg        [5:0]    endpoint_dmaLogic_length;
  wire       [5:0]    endpoint_dmaLogic_lengthMax;
  wire       [5:0]    endpoint_dmaLogic_lengthCalc;
  wire       [4:0]    endpoint_dmaLogic_beatCount;
  reg        [10:0]   endpoint_dmaLogic_fromUsbCounter;
  reg                 endpoint_dmaLogic_overflow;
  reg                 endpoint_dmaLogic_underflow;
  wire                endpoint_dmaLogic_underflowError;
  wire                when_UsbOhci_l937;
  reg        [12:0]   endpoint_dmaLogic_byteCtx_counter;
  wire                endpoint_dmaLogic_byteCtx_last;
  wire       [1:0]    endpoint_dmaLogic_byteCtx_sel;
  reg                 endpoint_dmaLogic_byteCtx_increment;
  reg                 endpoint_dmaLogic_toUsb_dmaReady;
  reg                 endpoint_dmaLogic_toUsb_run;
  wire                when_UsbOhci_l958;
  reg        [31:0]   endpoint_dmaLogic_fromUsb_buffer;
  reg                 endpoint_dmaLogic_fromUsb_push;
  reg                 endpoint_dmaLogic_fromUsb_start;
  reg                 endpoint_dmaLogic_fromUsb_run;
  wire                when_UsbOhci_l997;
  wire                endpoint_dmaLogic_fromUsb_dmaReady;
  reg        [13:0]   endpoint_dmaLogic_fromUsb_transactionSizeMax;
  wire                when_UsbOhci_l1011;
  wire       [3:0]    _zz_5;
  wire                when_UsbOhci_l1020;
  wire       [3:0]    endpoint_dmaLogic_headMask;
  wire       [3:0]    endpoint_dmaLogic_lastMask;
  wire       [3:0]    endpoint_dmaLogic_fullMask;
  wire                endpoint_dmaLogic_beatLast;
  reg                 endpoint_dmaLogic_storageReadDone;
  wire                endpoint_dmaLogic_headHit;
  wire                endpoint_dmaLogic_lastHit;
  reg                 endpoint_dmaLogic_inBurst;
  wire                endpoint_dmaLogic_fsmStopped;
  wire       [13:0]   endpoint_byteCountCalc;
  wire                endpoint_fsTimeCheck;
  wire                endpoint_timeCheck;
  reg                 endpoint_ackRxFired;
  reg                 endpoint_ackRxActivated;
  reg                 endpoint_ackRxPidFailure;
  reg                 endpoint_ackRxStuffing;
  reg        [3:0]    endpoint_ackRxPid;
  wire       [31:0]   endpoint_tdUpdateAddress;
  reg                 operational_wantExit;
  reg                 operational_wantStart;
  reg                 operational_wantKill;
  reg                 operational_periodicHeadFetched;
  reg                 operational_periodicDone;
  reg                 operational_allowBulk;
  reg                 operational_allowControl;
  reg                 operational_allowPeriodic;
  reg                 operational_allowIsochronous;
  reg                 operational_askExit;
  wire                hc_wantExit;
  reg                 hc_wantStart;
  wire                hc_wantKill;
  reg                 hc_error;
  wire                hc_operationalIsDone;
  wire       [1:0]    _zz_reg_hcControl_HCFSWrite_payload;
  wire                when_BusSlaveFactory_l1041;
  wire                when_BusSlaveFactory_l1041_1;
  wire                when_BusSlaveFactory_l1041_2;
  wire                when_BusSlaveFactory_l1041_3;
  wire                when_BusSlaveFactory_l1041_4;
  wire                when_BusSlaveFactory_l1041_5;
  wire                when_BusSlaveFactory_l1041_6;
  wire                when_BusSlaveFactory_l1041_7;
  wire                when_BusSlaveFactory_l1041_8;
  wire                when_BusSlaveFactory_l1041_9;
  wire                when_BusSlaveFactory_l1041_10;
  wire                when_BusSlaveFactory_l1041_11;
  wire                when_BusSlaveFactory_l1041_12;
  wire                when_BusSlaveFactory_l1041_13;
  wire                when_BusSlaveFactory_l1041_14;
  wire                when_BusSlaveFactory_l1041_15;
  wire                when_BusSlaveFactory_l1041_16;
  wire                when_BusSlaveFactory_l1041_17;
  wire                when_BusSlaveFactory_l1041_18;
  wire                when_BusSlaveFactory_l1041_19;
  wire                when_BusSlaveFactory_l1041_20;
  wire                when_BusSlaveFactory_l1041_21;
  wire                when_BusSlaveFactory_l1041_22;
  wire                when_BusSlaveFactory_l1041_23;
  wire                when_BusSlaveFactory_l1041_24;
  wire                when_BusSlaveFactory_l1041_25;
  wire                when_BusSlaveFactory_l1041_26;
  wire                when_BusSlaveFactory_l1041_27;
  wire                when_BusSlaveFactory_l1041_28;
  wire                when_BusSlaveFactory_l1041_29;
  wire                when_BusSlaveFactory_l1041_30;
  wire                when_BusSlaveFactory_l1041_31;
  wire                when_BusSlaveFactory_l1041_32;
  wire                when_BusSlaveFactory_l1041_33;
  wire                when_BusSlaveFactory_l1041_34;
  wire                when_BusSlaveFactory_l1041_35;
  wire                when_BusSlaveFactory_l1041_36;
  wire                when_BusSlaveFactory_l1041_37;
  wire                when_BusSlaveFactory_l1041_38;
  wire                when_BusSlaveFactory_l1041_39;
  wire                when_BusSlaveFactory_l1041_40;
  wire                when_BusSlaveFactory_l1041_41;
  wire                when_BusSlaveFactory_l1041_42;
  wire                when_BusSlaveFactory_l1041_43;
  wire                when_BusSlaveFactory_l1041_44;
  wire                when_BusSlaveFactory_l1041_45;
  wire                when_BusSlaveFactory_l1041_46;
  reg                 _zz_when_UsbOhci_l241;
  wire                when_UsbOhci_l241;
  reg        [2:0]    token_stateReg;
  reg        [2:0]    token_stateNext;
  wire                when_StateMachine_l237;
  wire                unscheduleAll_fire;
  reg        [2:0]    dataTx_stateReg;
  reg        [2:0]    dataTx_stateNext;
  reg        [1:0]    dataRx_stateReg;
  reg        [1:0]    dataRx_stateNext;
  wire                when_Misc_l64;
  wire                when_Misc_l70;
  wire                when_Misc_l71;
  wire                when_Misc_l78;
  wire                when_StateMachine_l253;
  wire                when_Misc_l85;
  reg        [1:0]    sof_stateReg;
  reg        [1:0]    sof_stateNext;
  wire                when_UsbOhci_l207;
  wire                when_UsbOhci_l207_1;
  wire                when_UsbOhci_l614;
  wire                when_StateMachine_l237_1;
  reg        [4:0]    endpoint_stateReg;
  reg        [4:0]    endpoint_stateNext;
  wire                when_UsbOhci_l1366;
  wire                when_UsbOhci_l189;
  wire                when_UsbOhci_l189_1;
  wire                when_UsbOhci_l189_2;
  wire                when_UsbOhci_l189_3;
  wire                when_UsbOhci_l843;
  wire                when_UsbOhci_l849;
  wire                when_UsbOhci_l189_4;
  wire                when_UsbOhci_l189_5;
  wire                when_UsbOhci_l189_6;
  wire                when_UsbOhci_l189_7;
  wire                when_UsbOhci_l879;
  wire                when_UsbOhci_l189_8;
  wire                when_UsbOhci_l189_9;
  wire                when_UsbOhci_l879_1;
  wire                when_UsbOhci_l189_10;
  wire                when_UsbOhci_l189_11;
  wire                when_UsbOhci_l879_2;
  wire                when_UsbOhci_l189_12;
  wire                when_UsbOhci_l189_13;
  wire                when_UsbOhci_l879_3;
  wire                when_UsbOhci_l189_14;
  wire                when_UsbOhci_l189_15;
  wire                when_UsbOhci_l879_4;
  wire                when_UsbOhci_l189_16;
  wire                when_UsbOhci_l189_17;
  wire                when_UsbOhci_l879_5;
  wire                when_UsbOhci_l189_18;
  wire                when_UsbOhci_l189_19;
  wire                when_UsbOhci_l879_6;
  wire                when_UsbOhci_l189_20;
  wire                when_UsbOhci_l189_21;
  wire                when_UsbOhci_l879_7;
  wire                when_UsbOhci_l189_22;
  wire                when_UsbOhci_l886;
  wire       [13:0]   _zz_endpoint_lastAddress;
  wire                when_UsbOhci_l1173;
  reg                 when_UsbOhci_l1329;
  wire                when_UsbOhci_l1318;
  wire                when_UsbOhci_l1338;
  wire                when_UsbOhci_l1255;
  wire                when_UsbOhci_l1260;
  wire                when_UsbOhci_l1262;
  wire                when_UsbOhci_l1386;
  wire                when_UsbOhci_l1401;
  wire                when_UsbOhci_l207_2;
  wire                when_UsbOhci_l207_3;
  wire       [15:0]   _zz_ioDma_cmd_payload_fragment_data;
  wire                when_UsbOhci_l1433;
  wire                when_UsbOhci_l207_4;
  wire                when_UsbOhci_l1433_1;
  wire                when_UsbOhci_l207_5;
  wire                when_UsbOhci_l1433_2;
  wire                when_UsbOhci_l207_6;
  wire                when_UsbOhci_l1433_3;
  wire                when_UsbOhci_l207_7;
  wire                when_UsbOhci_l1433_4;
  wire                when_UsbOhci_l207_8;
  wire                when_UsbOhci_l1433_5;
  wire                when_UsbOhci_l207_9;
  wire                when_UsbOhci_l1433_6;
  wire                when_UsbOhci_l207_10;
  wire                when_UsbOhci_l1433_7;
  wire                when_UsbOhci_l207_11;
  wire                when_UsbOhci_l207_12;
  wire                when_UsbOhci_l207_13;
  wire                when_UsbOhci_l207_14;
  wire                when_UsbOhci_l1448;
  wire                when_UsbOhci_l207_15;
  wire                when_UsbOhci_l1463;
  wire                when_UsbOhci_l1470;
  wire                when_UsbOhci_l1473;
  wire                when_StateMachine_l237_2;
  wire                when_StateMachine_l253_1;
  wire                when_StateMachine_l253_2;
  wire                when_StateMachine_l253_3;
  wire                when_StateMachine_l253_4;
  reg        [2:0]    endpoint_dmaLogic_stateReg;
  reg        [2:0]    endpoint_dmaLogic_stateNext;
  wire                when_UsbOhci_l1047;
  wire                when_UsbOhci_l1057;
  wire                when_UsbOhci_l1093;
  wire                when_UsbOhci_l1098;
  wire                when_StateMachine_l253_5;
  wire                when_UsbOhci_l973;
  reg        [2:0]    operational_stateReg;
  reg        [2:0]    operational_stateNext;
  wire                when_UsbOhci_l1516;
  wire                when_UsbOhci_l1543;
  wire                when_UsbOhci_l1542;
  wire                when_StateMachine_l237_3;
  wire                when_StateMachine_l253_6;
  reg        [2:0]    hc_stateReg;
  reg        [2:0]    hc_stateNext;
  wire                when_UsbOhci_l1671;
  wire                when_UsbOhci_l1680;
  wire                when_UsbOhci_l1683;
  wire                when_UsbOhci_l1694;
  wire                when_UsbOhci_l1707;
  wire                when_StateMachine_l253_7;
  wire                when_StateMachine_l253_8;
  wire                when_StateMachine_l253_9;
  wire                when_UsbOhci_l1714;
  `ifndef SYNTHESIS
  reg [87:0] reg_hcControl_HCFS_string;
  reg [87:0] reg_hcControl_HCFSWrite_payload_string;
  reg [63:0] endpoint_flowType_string;
  reg [79:0] endpoint_status_1_string;
  reg [87:0] _zz_reg_hcControl_HCFSWrite_payload_string;
  reg [31:0] token_stateReg_string;
  reg [31:0] token_stateNext_string;
  reg [39:0] dataTx_stateReg_string;
  reg [39:0] dataTx_stateNext_string;
  reg [31:0] dataRx_stateReg_string;
  reg [31:0] dataRx_stateNext_string;
  reg [127:0] sof_stateReg_string;
  reg [127:0] sof_stateNext_string;
  reg [135:0] endpoint_stateReg_string;
  reg [135:0] endpoint_stateNext_string;
  reg [79:0] endpoint_dmaLogic_stateReg_string;
  reg [79:0] endpoint_dmaLogic_stateNext_string;
  reg [135:0] operational_stateReg_string;
  reg [135:0] operational_stateNext_string;
  reg [111:0] hc_stateReg_string;
  reg [111:0] hc_stateNext_string;
  `endif

  reg [31:0] endpoint_dmaLogic_storage_ram [0:63];

  assign _zz_dmaCtx_pendingCounter = (dmaCtx_pendingCounter + _zz_dmaCtx_pendingCounter_1);
  assign _zz_dmaCtx_pendingCounter_2 = (ioDma_cmd_fire && ioDma_cmd_payload_last);
  assign _zz_dmaCtx_pendingCounter_1 = {3'd0, _zz_dmaCtx_pendingCounter_2};
  assign _zz_dmaCtx_pendingCounter_4 = (ioDma_rsp_fire && ioDma_rsp_payload_last);
  assign _zz_dmaCtx_pendingCounter_3 = {3'd0, _zz_dmaCtx_pendingCounter_4};
  assign _zz_reg_hcCommandStatus_startSoftReset = 1'b1;
  assign _zz_reg_hcCommandStatus_CLF = 1'b1;
  assign _zz_reg_hcCommandStatus_BLF = 1'b1;
  assign _zz_reg_hcCommandStatus_OCR = 1'b1;
  assign _zz_reg_hcInterrupt_MIE = 1'b1;
  assign _zz_reg_hcInterrupt_MIE_1 = 1'b0;
  assign _zz_reg_hcInterrupt_SO_status = 1'b0;
  assign _zz_reg_hcInterrupt_SO_enable = 1'b1;
  assign _zz_reg_hcInterrupt_SO_enable_1 = 1'b0;
  assign _zz_reg_hcInterrupt_WDH_status = 1'b0;
  assign _zz_reg_hcInterrupt_WDH_enable = 1'b1;
  assign _zz_reg_hcInterrupt_WDH_enable_1 = 1'b0;
  assign _zz_reg_hcInterrupt_SF_status = 1'b0;
  assign _zz_reg_hcInterrupt_SF_enable = 1'b1;
  assign _zz_reg_hcInterrupt_SF_enable_1 = 1'b0;
  assign _zz_reg_hcInterrupt_RD_status = 1'b0;
  assign _zz_reg_hcInterrupt_RD_enable = 1'b1;
  assign _zz_reg_hcInterrupt_RD_enable_1 = 1'b0;
  assign _zz_reg_hcInterrupt_UE_status = 1'b0;
  assign _zz_reg_hcInterrupt_UE_enable = 1'b1;
  assign _zz_reg_hcInterrupt_UE_enable_1 = 1'b0;
  assign _zz_reg_hcInterrupt_FNO_status = 1'b0;
  assign _zz_reg_hcInterrupt_FNO_enable = 1'b1;
  assign _zz_reg_hcInterrupt_FNO_enable_1 = 1'b0;
  assign _zz_reg_hcInterrupt_RHSC_status = 1'b0;
  assign _zz_reg_hcInterrupt_RHSC_enable = 1'b1;
  assign _zz_reg_hcInterrupt_RHSC_enable_1 = 1'b0;
  assign _zz_reg_hcInterrupt_OC_status = 1'b0;
  assign _zz_reg_hcInterrupt_OC_enable = 1'b1;
  assign _zz_reg_hcInterrupt_OC_enable_1 = 1'b0;
  assign _zz_reg_hcLSThreshold_hit = {2'd0, reg_hcLSThreshold_LST};
  assign _zz_reg_hcRhStatus_CCIC = 1'b0;
  assign _zz_reg_hcRhStatus_clearGlobalPower = 1'b1;
  assign _zz_reg_hcRhStatus_setRemoteWakeupEnable = 1'b1;
  assign _zz_reg_hcRhStatus_setGlobalPower = 1'b1;
  assign _zz_reg_hcRhStatus_clearRemoteWakeupEnable = 1'b1;
  assign _zz_reg_hcRhPortStatus_0_clearPortEnable = 1'b1;
  assign _zz_reg_hcRhPortStatus_0_setPortEnable = 1'b1;
  assign _zz_reg_hcRhPortStatus_0_setPortSuspend = 1'b1;
  assign _zz_reg_hcRhPortStatus_0_clearSuspendStatus = 1'b1;
  assign _zz_reg_hcRhPortStatus_0_setPortReset = 1'b1;
  assign _zz_reg_hcRhPortStatus_0_setPortPower = 1'b1;
  assign _zz_reg_hcRhPortStatus_0_clearPortPower = 1'b1;
  assign _zz_reg_hcRhPortStatus_0_CSC_clear = 1'b1;
  assign _zz_reg_hcRhPortStatus_0_PESC_clear = 1'b1;
  assign _zz_reg_hcRhPortStatus_0_PSSC_clear = 1'b1;
  assign _zz_reg_hcRhPortStatus_0_OCIC_clear = 1'b1;
  assign _zz_reg_hcRhPortStatus_0_PRSC_clear = 1'b1;
  assign _zz_reg_hcRhPortStatus_1_clearPortEnable = 1'b1;
  assign _zz_reg_hcRhPortStatus_1_setPortEnable = 1'b1;
  assign _zz_reg_hcRhPortStatus_1_setPortSuspend = 1'b1;
  assign _zz_reg_hcRhPortStatus_1_clearSuspendStatus = 1'b1;
  assign _zz_reg_hcRhPortStatus_1_setPortReset = 1'b1;
  assign _zz_reg_hcRhPortStatus_1_setPortPower = 1'b1;
  assign _zz_reg_hcRhPortStatus_1_clearPortPower = 1'b1;
  assign _zz_reg_hcRhPortStatus_1_CSC_clear = 1'b1;
  assign _zz_reg_hcRhPortStatus_1_PESC_clear = 1'b1;
  assign _zz_reg_hcRhPortStatus_1_PSSC_clear = 1'b1;
  assign _zz_reg_hcRhPortStatus_1_OCIC_clear = 1'b1;
  assign _zz_reg_hcRhPortStatus_1_PRSC_clear = 1'b1;
  assign _zz_rxTimer_ackTx_1 = (rxTimer_lowSpeed ? 4'b1111 : 4'b0001);
  assign _zz_rxTimer_ackTx = {4'd0, _zz_rxTimer_ackTx_1};
  assign _zz_endpoint_TD_isoOverrun = {13'd0, endpoint_TD_FC};
  assign _zz_endpoint_TD_firstOffset_1 = endpoint_TD_CBP[11 : 0];
  assign _zz_endpoint_TD_firstOffset = {1'd0, _zz_endpoint_TD_firstOffset_1};
  assign _zz_endpoint_TD_lastOffset = (endpoint_TD_isoBaseNext - _zz_endpoint_TD_lastOffset_1);
  assign _zz_endpoint_TD_lastOffset_2 = (! endpoint_TD_isoLast);
  assign _zz_endpoint_TD_lastOffset_1 = {12'd0, _zz_endpoint_TD_lastOffset_2};
  assign _zz_endpoint_currentAddressBmb = (endpoint_currentAddressFull >>> 3'd6);
  assign _zz_endpoint_transactionSizeMinusOne = {1'd0, endpoint_lastAddress};
  assign _zz_endpoint_dataDone = {1'd0, endpoint_lastAddress};
  assign _zz_endpoint_dmaLogic_storage_full_2 = endpoint_currentAddress[13 : 6];
  assign _zz_endpoint_dmaLogic_storage_full_1 = _zz_endpoint_dmaLogic_storage_full_2[2:0];
  assign _zz_endpoint_dmaLogic_lengthMax = endpoint_currentAddress[5:0];
  assign _zz_endpoint_dmaLogic_lengthCalc = ((endpoint_transactionSizeMinusOne < _zz_endpoint_dmaLogic_lengthCalc_1) ? endpoint_transactionSizeMinusOne : _zz_endpoint_dmaLogic_lengthCalc_2);
  assign _zz_endpoint_dmaLogic_lengthCalc_1 = {8'd0, endpoint_dmaLogic_lengthMax};
  assign _zz_endpoint_dmaLogic_lengthCalc_2 = {8'd0, endpoint_dmaLogic_lengthMax};
  assign _zz_endpoint_dmaLogic_beatCount = ({1'b0,endpoint_dmaLogic_length} + _zz_endpoint_dmaLogic_beatCount_1);
  assign _zz_endpoint_dmaLogic_beatCount_2 = endpoint_currentAddressFull[1 : 0];
  assign _zz_endpoint_dmaLogic_beatCount_1 = {5'd0, _zz_endpoint_dmaLogic_beatCount_2};
  assign _zz_endpoint_dmaLogic_fromUsb_dmaReady = (endpoint_dmaLogic_storage_writePtr ^ endpoint_dmaLogic_storage_readPtr);
  assign _zz_when_UsbOhci_l1011 = {3'd0, endpoint_dmaLogic_fromUsbCounter};
  assign _zz_endpoint_dmaLogic_overflow = {3'd0, endpoint_dmaLogic_fromUsbCounter};
  assign _zz_endpoint_lastAddress_1 = (endpoint_TD_firstOffset + _zz_endpoint_lastAddress_2);
  assign _zz_endpoint_lastAddress_2 = {2'd0, endpoint_dmaLogic_fromUsbCounter};
  assign _zz_endpoint_dmaLogic_fromUsbCounter_1 = (! endpoint_dmaLogic_fromUsbCounter[10]);
  assign _zz_endpoint_dmaLogic_fromUsbCounter = {10'd0, _zz_endpoint_dmaLogic_fromUsbCounter_1};
  assign _zz_endpoint_dmaLogic_lastMask = (endpoint_currentAddress + _zz_endpoint_dmaLogic_lastMask_1);
  assign _zz_endpoint_dmaLogic_lastMask_1 = {8'd0, endpoint_dmaLogic_length};
  assign _zz_endpoint_dmaLogic_lastMask_2 = (endpoint_currentAddress + _zz_endpoint_dmaLogic_lastMask_3);
  assign _zz_endpoint_dmaLogic_lastMask_3 = {8'd0, endpoint_dmaLogic_length};
  assign _zz_endpoint_dmaLogic_lastMask_4 = (endpoint_currentAddress + _zz_endpoint_dmaLogic_lastMask_5);
  assign _zz_endpoint_dmaLogic_lastMask_5 = {8'd0, endpoint_dmaLogic_length};
  assign _zz_endpoint_dmaLogic_lastMask_6 = (endpoint_currentAddress + _zz_endpoint_dmaLogic_lastMask_7);
  assign _zz_endpoint_dmaLogic_lastMask_7 = {8'd0, endpoint_dmaLogic_length};
  assign _zz_endpoint_dmaLogic_headHit_1 = endpoint_currentAddress[13 : 2];
  assign _zz_endpoint_dmaLogic_headHit = _zz_endpoint_dmaLogic_headHit_1[3:0];
  assign _zz_endpoint_dmaLogic_lastHit_1 = _zz_endpoint_dmaLogic_lastHit_2[13 : 2];
  assign _zz_endpoint_dmaLogic_lastHit = _zz_endpoint_dmaLogic_lastHit_1[3:0];
  assign _zz_endpoint_dmaLogic_lastHit_2 = (endpoint_currentAddress + _zz_endpoint_dmaLogic_lastHit_3);
  assign _zz_endpoint_dmaLogic_lastHit_3 = {8'd0, endpoint_dmaLogic_length};
  assign _zz_endpoint_byteCountCalc = (_zz_endpoint_byteCountCalc_1 - endpoint_currentAddress);
  assign _zz_endpoint_byteCountCalc_1 = {1'd0, endpoint_lastAddress};
  assign _zz_endpoint_fsTimeCheck = {2'd0, frame_limitCounter};
  assign _zz_endpoint_fsTimeCheck_1 = ({3'd0,endpoint_byteCountCalc} <<< 2'd3);
  assign _zz_token_data = reg_hcFmNumber_FN;
  assign _zz_ioDma_cmd_payload_fragment_length = (endpoint_ED_F ? 5'h1f : 5'h0f);
  assign _zz__zz_endpoint_lastAddress = ({1'b0,endpoint_TD_firstOffset} + _zz__zz_endpoint_lastAddress_1);
  assign _zz__zz_endpoint_lastAddress_2 = {1'b0,endpoint_ED_MPS};
  assign _zz__zz_endpoint_lastAddress_1 = {2'd0, _zz__zz_endpoint_lastAddress_2};
  assign _zz_endpoint_lastAddress_3 = (endpoint_ED_F ? _zz_endpoint_lastAddress_4 : ((_zz_endpoint_lastAddress_5 < _zz_endpoint_lastAddress) ? _zz_endpoint_lastAddress_6 : _zz_endpoint_lastAddress));
  assign _zz_endpoint_lastAddress_4 = {1'd0, endpoint_TD_lastOffset};
  assign _zz_endpoint_lastAddress_5 = {1'd0, endpoint_TD_lastOffset};
  assign _zz_endpoint_lastAddress_6 = {1'd0, endpoint_TD_lastOffset};
  assign _zz_when_UsbOhci_l1386 = {1'd0, endpoint_TD_lastOffset};
  assign _zz_endpoint_TD_words_0 = (endpoint_TD_EC + 2'b01);
  assign _zz_ioDma_cmd_payload_fragment_length_1 = (endpoint_ED_F ? 5'h1f : 5'h0f);
  assign _zz_ioDma_cmd_payload_last_1 = (endpoint_ED_F ? 3'b111 : 3'b011);
  assign _zz_ioDma_cmd_payload_last = {1'd0, _zz_ioDma_cmd_payload_last_1};
  assign _zz__zz_ioDma_cmd_payload_fragment_data_1 = (endpoint_ED_isoOut ? 14'h0 : _zz__zz_ioDma_cmd_payload_fragment_data_2);
  assign _zz__zz_ioDma_cmd_payload_fragment_data = _zz__zz_ioDma_cmd_payload_fragment_data_1[11:0];
  assign _zz__zz_ioDma_cmd_payload_fragment_data_2 = (endpoint_currentAddress - _zz__zz_ioDma_cmd_payload_fragment_data_3);
  assign _zz__zz_ioDma_cmd_payload_fragment_data_3 = {1'd0, endpoint_TD_isoBase};
  assign _zz_endpoint_dmaLogic_storage_writePtr = endpoint_currentAddress[13 : 2];
  assign _zz_endpoint_dmaLogic_storage_readPtr = _zz_endpoint_dmaLogic_storage_readPtr_1[13 : 2];
  assign _zz_endpoint_dmaLogic_storage_readPtr_1 = ({6'd0,_zz_endpoint_dmaLogic_storage_readPtr_2} <<< 3'd6);
  assign _zz_endpoint_dmaLogic_storage_readPtr_2 = (endpoint_currentAddress >>> 3'd6);
  assign _zz_endpoint_dmaLogic_storage_writePtr_1 = _zz_endpoint_dmaLogic_storage_writePtr_2[13 : 2];
  assign _zz_endpoint_dmaLogic_storage_writePtr_2 = ({6'd0,_zz_endpoint_dmaLogic_storage_writePtr_3} <<< 3'd6);
  assign _zz_endpoint_dmaLogic_storage_writePtr_3 = (endpoint_currentAddress >>> 3'd6);
  assign _zz_endpoint_dmaLogic_storage_readPtr_3 = endpoint_currentAddress[13 : 2];
  assign _zz_endpoint_dmaLogic_fromUsb_transactionSizeMax = (_zz_endpoint_dmaLogic_fromUsb_transactionSizeMax_1 - endpoint_currentAddress);
  assign _zz_endpoint_dmaLogic_fromUsb_transactionSizeMax_1 = {1'd0, endpoint_lastAddress};
  assign _zz_endpoint_currentAddress = (endpoint_currentAddress + _zz_endpoint_currentAddress_1);
  assign _zz_endpoint_currentAddress_1 = {8'd0, endpoint_dmaLogic_length};
  assign _zz_endpoint_currentAddress_2 = (endpoint_currentAddress + _zz_endpoint_currentAddress_3);
  assign _zz_endpoint_currentAddress_3 = {8'd0, endpoint_dmaLogic_length};
  assign _zz_ioDma_cmd_payload_fragment_address_1 = ({2'd0,reg_hcFmNumber_FN[4 : 0]} <<< 2'd2);
  assign _zz_ioDma_cmd_payload_fragment_address = {25'd0, _zz_ioDma_cmd_payload_fragment_address_1};
  always @(posedge clk_peripheral) begin
    if(endpoint_dmaLogic_storage_readCmd_fire) begin
      endpoint_dmaLogic_storage_ram_spinal_port0 <= endpoint_dmaLogic_storage_ram[endpoint_dmaLogic_storage_readCmd_payload];
    end
  end

  always @(posedge clk_peripheral) begin
    if(_zz_1) begin
      endpoint_dmaLogic_storage_ram[endpoint_dmaLogic_storage_write_payload_address] <= endpoint_dmaLogic_storage_write_payload_data;
    end
  end

  Crc token_crc5 (
    .io_flush         (token_crc5_io_flush          ), //i
    .io_input_valid   (token_crc5_io_input_valid    ), //i
    .io_input_payload (token_data[10:0]             ), //i
    .io_result        (token_crc5_io_result[4:0]    ), //o
    .io_resultNext    (token_crc5_io_resultNext[4:0]), //o
    .clk_peripheral   (clk_peripheral               ), //i
    .reset_peripheral (reset_peripheral             )  //i
  );
  Crc_1 dataTx_crc16 (
    .io_flush         (dataTx_crc16_io_flush            ), //i
    .io_input_valid   (dataTx_data_fire                 ), //i
    .io_input_payload (dataTx_data_payload_fragment[7:0]), //i
    .io_result        (dataTx_crc16_io_result[15:0]     ), //o
    .io_resultNext    (dataTx_crc16_io_resultNext[15:0] ), //o
    .clk_peripheral   (clk_peripheral                   ), //i
    .reset_peripheral (reset_peripheral                 )  //i
  );
  Crc_2 dataRx_crc16 (
    .io_flush         (dataRx_crc16_io_flush           ), //i
    .io_input_valid   (dataRx_crc16_io_input_valid     ), //i
    .io_input_payload (_zz_dataRx_pid[7:0]             ), //i
    .io_result        (dataRx_crc16_io_result[15:0]    ), //o
    .io_resultNext    (dataRx_crc16_io_resultNext[15:0]), //o
    .clk_peripheral   (clk_peripheral                  ), //i
    .reset_peripheral (reset_peripheral                )  //i
  );
  always @(*) begin
    case(endpoint_dmaLogic_byteCtx_sel)
      2'b00 : _zz_dataTx_data_payload_fragment = endpoint_dmaLogic_storage_readRsp_payload[7 : 0];
      2'b01 : _zz_dataTx_data_payload_fragment = endpoint_dmaLogic_storage_readRsp_payload[15 : 8];
      2'b10 : _zz_dataTx_data_payload_fragment = endpoint_dmaLogic_storage_readRsp_payload[23 : 16];
      default : _zz_dataTx_data_payload_fragment = endpoint_dmaLogic_storage_readRsp_payload[31 : 24];
    endcase
  end

  `ifndef SYNTHESIS
  always @(*) begin
    case(reg_hcControl_HCFS)
      MainState_RESET : reg_hcControl_HCFS_string = "RESET      ";
      MainState_RESUME : reg_hcControl_HCFS_string = "RESUME     ";
      MainState_OPERATIONAL : reg_hcControl_HCFS_string = "OPERATIONAL";
      MainState_SUSPEND : reg_hcControl_HCFS_string = "SUSPEND    ";
      default : reg_hcControl_HCFS_string = "???????????";
    endcase
  end
  always @(*) begin
    case(reg_hcControl_HCFSWrite_payload)
      MainState_RESET : reg_hcControl_HCFSWrite_payload_string = "RESET      ";
      MainState_RESUME : reg_hcControl_HCFSWrite_payload_string = "RESUME     ";
      MainState_OPERATIONAL : reg_hcControl_HCFSWrite_payload_string = "OPERATIONAL";
      MainState_SUSPEND : reg_hcControl_HCFSWrite_payload_string = "SUSPEND    ";
      default : reg_hcControl_HCFSWrite_payload_string = "???????????";
    endcase
  end
  always @(*) begin
    case(endpoint_flowType)
      FlowType_BULK : endpoint_flowType_string = "BULK    ";
      FlowType_CONTROL : endpoint_flowType_string = "CONTROL ";
      FlowType_PERIODIC : endpoint_flowType_string = "PERIODIC";
      default : endpoint_flowType_string = "????????";
    endcase
  end
  always @(*) begin
    case(endpoint_status_1)
      endpoint_Status_OK : endpoint_status_1_string = "OK        ";
      endpoint_Status_FRAME_TIME : endpoint_status_1_string = "FRAME_TIME";
      default : endpoint_status_1_string = "??????????";
    endcase
  end
  always @(*) begin
    case(_zz_reg_hcControl_HCFSWrite_payload)
      MainState_RESET : _zz_reg_hcControl_HCFSWrite_payload_string = "RESET      ";
      MainState_RESUME : _zz_reg_hcControl_HCFSWrite_payload_string = "RESUME     ";
      MainState_OPERATIONAL : _zz_reg_hcControl_HCFSWrite_payload_string = "OPERATIONAL";
      MainState_SUSPEND : _zz_reg_hcControl_HCFSWrite_payload_string = "SUSPEND    ";
      default : _zz_reg_hcControl_HCFSWrite_payload_string = "???????????";
    endcase
  end
  always @(*) begin
    case(token_stateReg)
      token_enumDef_BOOT : token_stateReg_string = "BOOT";
      token_enumDef_INIT : token_stateReg_string = "INIT";
      token_enumDef_PID : token_stateReg_string = "PID ";
      token_enumDef_B1 : token_stateReg_string = "B1  ";
      token_enumDef_B2 : token_stateReg_string = "B2  ";
      token_enumDef_EOP : token_stateReg_string = "EOP ";
      default : token_stateReg_string = "????";
    endcase
  end
  always @(*) begin
    case(token_stateNext)
      token_enumDef_BOOT : token_stateNext_string = "BOOT";
      token_enumDef_INIT : token_stateNext_string = "INIT";
      token_enumDef_PID : token_stateNext_string = "PID ";
      token_enumDef_B1 : token_stateNext_string = "B1  ";
      token_enumDef_B2 : token_stateNext_string = "B2  ";
      token_enumDef_EOP : token_stateNext_string = "EOP ";
      default : token_stateNext_string = "????";
    endcase
  end
  always @(*) begin
    case(dataTx_stateReg)
      dataTx_enumDef_BOOT : dataTx_stateReg_string = "BOOT ";
      dataTx_enumDef_PID : dataTx_stateReg_string = "PID  ";
      dataTx_enumDef_DATA : dataTx_stateReg_string = "DATA ";
      dataTx_enumDef_CRC_0 : dataTx_stateReg_string = "CRC_0";
      dataTx_enumDef_CRC_1 : dataTx_stateReg_string = "CRC_1";
      dataTx_enumDef_EOP : dataTx_stateReg_string = "EOP  ";
      default : dataTx_stateReg_string = "?????";
    endcase
  end
  always @(*) begin
    case(dataTx_stateNext)
      dataTx_enumDef_BOOT : dataTx_stateNext_string = "BOOT ";
      dataTx_enumDef_PID : dataTx_stateNext_string = "PID  ";
      dataTx_enumDef_DATA : dataTx_stateNext_string = "DATA ";
      dataTx_enumDef_CRC_0 : dataTx_stateNext_string = "CRC_0";
      dataTx_enumDef_CRC_1 : dataTx_stateNext_string = "CRC_1";
      dataTx_enumDef_EOP : dataTx_stateNext_string = "EOP  ";
      default : dataTx_stateNext_string = "?????";
    endcase
  end
  always @(*) begin
    case(dataRx_stateReg)
      dataRx_enumDef_BOOT : dataRx_stateReg_string = "BOOT";
      dataRx_enumDef_IDLE : dataRx_stateReg_string = "IDLE";
      dataRx_enumDef_PID : dataRx_stateReg_string = "PID ";
      dataRx_enumDef_DATA : dataRx_stateReg_string = "DATA";
      default : dataRx_stateReg_string = "????";
    endcase
  end
  always @(*) begin
    case(dataRx_stateNext)
      dataRx_enumDef_BOOT : dataRx_stateNext_string = "BOOT";
      dataRx_enumDef_IDLE : dataRx_stateNext_string = "IDLE";
      dataRx_enumDef_PID : dataRx_stateNext_string = "PID ";
      dataRx_enumDef_DATA : dataRx_stateNext_string = "DATA";
      default : dataRx_stateNext_string = "????";
    endcase
  end
  always @(*) begin
    case(sof_stateReg)
      sof_enumDef_BOOT : sof_stateReg_string = "BOOT            ";
      sof_enumDef_FRAME_TX : sof_stateReg_string = "FRAME_TX        ";
      sof_enumDef_FRAME_NUMBER_CMD : sof_stateReg_string = "FRAME_NUMBER_CMD";
      sof_enumDef_FRAME_NUMBER_RSP : sof_stateReg_string = "FRAME_NUMBER_RSP";
      default : sof_stateReg_string = "????????????????";
    endcase
  end
  always @(*) begin
    case(sof_stateNext)
      sof_enumDef_BOOT : sof_stateNext_string = "BOOT            ";
      sof_enumDef_FRAME_TX : sof_stateNext_string = "FRAME_TX        ";
      sof_enumDef_FRAME_NUMBER_CMD : sof_stateNext_string = "FRAME_NUMBER_CMD";
      sof_enumDef_FRAME_NUMBER_RSP : sof_stateNext_string = "FRAME_NUMBER_RSP";
      default : sof_stateNext_string = "????????????????";
    endcase
  end
  always @(*) begin
    case(endpoint_stateReg)
      endpoint_enumDef_BOOT : endpoint_stateReg_string = "BOOT             ";
      endpoint_enumDef_ED_READ_CMD : endpoint_stateReg_string = "ED_READ_CMD      ";
      endpoint_enumDef_ED_READ_RSP : endpoint_stateReg_string = "ED_READ_RSP      ";
      endpoint_enumDef_ED_ANALYSE : endpoint_stateReg_string = "ED_ANALYSE       ";
      endpoint_enumDef_TD_READ_CMD : endpoint_stateReg_string = "TD_READ_CMD      ";
      endpoint_enumDef_TD_READ_RSP : endpoint_stateReg_string = "TD_READ_RSP      ";
      endpoint_enumDef_TD_READ_DELAY : endpoint_stateReg_string = "TD_READ_DELAY    ";
      endpoint_enumDef_TD_ANALYSE : endpoint_stateReg_string = "TD_ANALYSE       ";
      endpoint_enumDef_TD_CHECK_TIME : endpoint_stateReg_string = "TD_CHECK_TIME    ";
      endpoint_enumDef_BUFFER_READ : endpoint_stateReg_string = "BUFFER_READ      ";
      endpoint_enumDef_TOKEN : endpoint_stateReg_string = "TOKEN            ";
      endpoint_enumDef_DATA_TX : endpoint_stateReg_string = "DATA_TX          ";
      endpoint_enumDef_DATA_RX : endpoint_stateReg_string = "DATA_RX          ";
      endpoint_enumDef_DATA_RX_VALIDATE : endpoint_stateReg_string = "DATA_RX_VALIDATE ";
      endpoint_enumDef_ACK_RX : endpoint_stateReg_string = "ACK_RX           ";
      endpoint_enumDef_ACK_TX_0 : endpoint_stateReg_string = "ACK_TX_0         ";
      endpoint_enumDef_ACK_TX_1 : endpoint_stateReg_string = "ACK_TX_1         ";
      endpoint_enumDef_ACK_TX_EOP : endpoint_stateReg_string = "ACK_TX_EOP       ";
      endpoint_enumDef_DATA_RX_WAIT_DMA : endpoint_stateReg_string = "DATA_RX_WAIT_DMA ";
      endpoint_enumDef_UPDATE_TD_PROCESS : endpoint_stateReg_string = "UPDATE_TD_PROCESS";
      endpoint_enumDef_UPDATE_TD_CMD : endpoint_stateReg_string = "UPDATE_TD_CMD    ";
      endpoint_enumDef_UPDATE_ED_CMD : endpoint_stateReg_string = "UPDATE_ED_CMD    ";
      endpoint_enumDef_UPDATE_SYNC : endpoint_stateReg_string = "UPDATE_SYNC      ";
      endpoint_enumDef_ABORD : endpoint_stateReg_string = "ABORD            ";
      default : endpoint_stateReg_string = "?????????????????";
    endcase
  end
  always @(*) begin
    case(endpoint_stateNext)
      endpoint_enumDef_BOOT : endpoint_stateNext_string = "BOOT             ";
      endpoint_enumDef_ED_READ_CMD : endpoint_stateNext_string = "ED_READ_CMD      ";
      endpoint_enumDef_ED_READ_RSP : endpoint_stateNext_string = "ED_READ_RSP      ";
      endpoint_enumDef_ED_ANALYSE : endpoint_stateNext_string = "ED_ANALYSE       ";
      endpoint_enumDef_TD_READ_CMD : endpoint_stateNext_string = "TD_READ_CMD      ";
      endpoint_enumDef_TD_READ_RSP : endpoint_stateNext_string = "TD_READ_RSP      ";
      endpoint_enumDef_TD_READ_DELAY : endpoint_stateNext_string = "TD_READ_DELAY    ";
      endpoint_enumDef_TD_ANALYSE : endpoint_stateNext_string = "TD_ANALYSE       ";
      endpoint_enumDef_TD_CHECK_TIME : endpoint_stateNext_string = "TD_CHECK_TIME    ";
      endpoint_enumDef_BUFFER_READ : endpoint_stateNext_string = "BUFFER_READ      ";
      endpoint_enumDef_TOKEN : endpoint_stateNext_string = "TOKEN            ";
      endpoint_enumDef_DATA_TX : endpoint_stateNext_string = "DATA_TX          ";
      endpoint_enumDef_DATA_RX : endpoint_stateNext_string = "DATA_RX          ";
      endpoint_enumDef_DATA_RX_VALIDATE : endpoint_stateNext_string = "DATA_RX_VALIDATE ";
      endpoint_enumDef_ACK_RX : endpoint_stateNext_string = "ACK_RX           ";
      endpoint_enumDef_ACK_TX_0 : endpoint_stateNext_string = "ACK_TX_0         ";
      endpoint_enumDef_ACK_TX_1 : endpoint_stateNext_string = "ACK_TX_1         ";
      endpoint_enumDef_ACK_TX_EOP : endpoint_stateNext_string = "ACK_TX_EOP       ";
      endpoint_enumDef_DATA_RX_WAIT_DMA : endpoint_stateNext_string = "DATA_RX_WAIT_DMA ";
      endpoint_enumDef_UPDATE_TD_PROCESS : endpoint_stateNext_string = "UPDATE_TD_PROCESS";
      endpoint_enumDef_UPDATE_TD_CMD : endpoint_stateNext_string = "UPDATE_TD_CMD    ";
      endpoint_enumDef_UPDATE_ED_CMD : endpoint_stateNext_string = "UPDATE_ED_CMD    ";
      endpoint_enumDef_UPDATE_SYNC : endpoint_stateNext_string = "UPDATE_SYNC      ";
      endpoint_enumDef_ABORD : endpoint_stateNext_string = "ABORD            ";
      default : endpoint_stateNext_string = "?????????????????";
    endcase
  end
  always @(*) begin
    case(endpoint_dmaLogic_stateReg)
      endpoint_dmaLogic_enumDef_BOOT : endpoint_dmaLogic_stateReg_string = "BOOT      ";
      endpoint_dmaLogic_enumDef_INIT : endpoint_dmaLogic_stateReg_string = "INIT      ";
      endpoint_dmaLogic_enumDef_TO_USB : endpoint_dmaLogic_stateReg_string = "TO_USB    ";
      endpoint_dmaLogic_enumDef_FROM_USB : endpoint_dmaLogic_stateReg_string = "FROM_USB  ";
      endpoint_dmaLogic_enumDef_VALIDATION : endpoint_dmaLogic_stateReg_string = "VALIDATION";
      endpoint_dmaLogic_enumDef_CALC_CMD : endpoint_dmaLogic_stateReg_string = "CALC_CMD  ";
      endpoint_dmaLogic_enumDef_READ_CMD : endpoint_dmaLogic_stateReg_string = "READ_CMD  ";
      endpoint_dmaLogic_enumDef_WRITE_CMD : endpoint_dmaLogic_stateReg_string = "WRITE_CMD ";
      default : endpoint_dmaLogic_stateReg_string = "??????????";
    endcase
  end
  always @(*) begin
    case(endpoint_dmaLogic_stateNext)
      endpoint_dmaLogic_enumDef_BOOT : endpoint_dmaLogic_stateNext_string = "BOOT      ";
      endpoint_dmaLogic_enumDef_INIT : endpoint_dmaLogic_stateNext_string = "INIT      ";
      endpoint_dmaLogic_enumDef_TO_USB : endpoint_dmaLogic_stateNext_string = "TO_USB    ";
      endpoint_dmaLogic_enumDef_FROM_USB : endpoint_dmaLogic_stateNext_string = "FROM_USB  ";
      endpoint_dmaLogic_enumDef_VALIDATION : endpoint_dmaLogic_stateNext_string = "VALIDATION";
      endpoint_dmaLogic_enumDef_CALC_CMD : endpoint_dmaLogic_stateNext_string = "CALC_CMD  ";
      endpoint_dmaLogic_enumDef_READ_CMD : endpoint_dmaLogic_stateNext_string = "READ_CMD  ";
      endpoint_dmaLogic_enumDef_WRITE_CMD : endpoint_dmaLogic_stateNext_string = "WRITE_CMD ";
      default : endpoint_dmaLogic_stateNext_string = "??????????";
    endcase
  end
  always @(*) begin
    case(operational_stateReg)
      operational_enumDef_BOOT : operational_stateReg_string = "BOOT             ";
      operational_enumDef_SOF : operational_stateReg_string = "SOF              ";
      operational_enumDef_ARBITER : operational_stateReg_string = "ARBITER          ";
      operational_enumDef_END_POINT : operational_stateReg_string = "END_POINT        ";
      operational_enumDef_PERIODIC_HEAD_CMD : operational_stateReg_string = "PERIODIC_HEAD_CMD";
      operational_enumDef_PERIODIC_HEAD_RSP : operational_stateReg_string = "PERIODIC_HEAD_RSP";
      operational_enumDef_WAIT_SOF : operational_stateReg_string = "WAIT_SOF         ";
      default : operational_stateReg_string = "?????????????????";
    endcase
  end
  always @(*) begin
    case(operational_stateNext)
      operational_enumDef_BOOT : operational_stateNext_string = "BOOT             ";
      operational_enumDef_SOF : operational_stateNext_string = "SOF              ";
      operational_enumDef_ARBITER : operational_stateNext_string = "ARBITER          ";
      operational_enumDef_END_POINT : operational_stateNext_string = "END_POINT        ";
      operational_enumDef_PERIODIC_HEAD_CMD : operational_stateNext_string = "PERIODIC_HEAD_CMD";
      operational_enumDef_PERIODIC_HEAD_RSP : operational_stateNext_string = "PERIODIC_HEAD_RSP";
      operational_enumDef_WAIT_SOF : operational_stateNext_string = "WAIT_SOF         ";
      default : operational_stateNext_string = "?????????????????";
    endcase
  end
  always @(*) begin
    case(hc_stateReg)
      hc_enumDef_BOOT : hc_stateReg_string = "BOOT          ";
      hc_enumDef_RESET : hc_stateReg_string = "RESET         ";
      hc_enumDef_RESUME : hc_stateReg_string = "RESUME        ";
      hc_enumDef_OPERATIONAL : hc_stateReg_string = "OPERATIONAL   ";
      hc_enumDef_SUSPEND : hc_stateReg_string = "SUSPEND       ";
      hc_enumDef_ANY_TO_RESET : hc_stateReg_string = "ANY_TO_RESET  ";
      hc_enumDef_ANY_TO_SUSPEND : hc_stateReg_string = "ANY_TO_SUSPEND";
      default : hc_stateReg_string = "??????????????";
    endcase
  end
  always @(*) begin
    case(hc_stateNext)
      hc_enumDef_BOOT : hc_stateNext_string = "BOOT          ";
      hc_enumDef_RESET : hc_stateNext_string = "RESET         ";
      hc_enumDef_RESUME : hc_stateNext_string = "RESUME        ";
      hc_enumDef_OPERATIONAL : hc_stateNext_string = "OPERATIONAL   ";
      hc_enumDef_SUSPEND : hc_stateNext_string = "SUSPEND       ";
      hc_enumDef_ANY_TO_RESET : hc_stateNext_string = "ANY_TO_RESET  ";
      hc_enumDef_ANY_TO_SUSPEND : hc_stateNext_string = "ANY_TO_SUSPEND";
      default : hc_stateNext_string = "??????????????";
    endcase
  end
  `endif

  always @(*) begin
    _zz_1 = 1'b0;
    if(endpoint_dmaLogic_storage_write_valid) begin
      _zz_1 = 1'b1;
    end
  end

  always @(*) begin
    io_phy_lowSpeed = 1'b0;
    if(when_UsbOhci_l738) begin
      io_phy_lowSpeed = endpoint_ED_S;
    end
  end

  always @(*) begin
    unscheduleAll_valid = 1'b0;
    if(doUnschedule) begin
      unscheduleAll_valid = 1'b1;
    end
  end

  always @(*) begin
    unscheduleAll_ready = 1'b1;
    if(when_UsbOhci_l158) begin
      unscheduleAll_ready = 1'b0;
    end
  end

  assign ioDma_cmd_fire = (ioDma_cmd_valid && ioDma_cmd_ready);
  assign ioDma_rsp_fire = (ioDma_rsp_valid && ioDma_rsp_ready);
  assign dmaCtx_pendingFull = dmaCtx_pendingCounter[3];
  assign dmaCtx_pendingEmpty = (dmaCtx_pendingCounter == 4'b0000);
  assign when_UsbOhci_l158 = (! dmaCtx_pendingEmpty);
  assign io_dma_cmd_fire = (io_dma_cmd_valid && io_dma_cmd_ready);
  assign _zz_io_dma_cmd_valid = (! (dmaCtx_pendingFull || (unscheduleAll_valid && io_dma_cmd_payload_first)));
  assign ioDma_cmd_ready = (io_dma_cmd_ready && _zz_io_dma_cmd_valid);
  assign io_dma_cmd_valid = (ioDma_cmd_valid && _zz_io_dma_cmd_valid);
  assign io_dma_cmd_payload_last = ioDma_cmd_payload_last;
  assign io_dma_cmd_payload_fragment_opcode = ioDma_cmd_payload_fragment_opcode;
  assign io_dma_cmd_payload_fragment_address = ioDma_cmd_payload_fragment_address;
  assign io_dma_cmd_payload_fragment_length = ioDma_cmd_payload_fragment_length;
  assign io_dma_cmd_payload_fragment_data = ioDma_cmd_payload_fragment_data;
  assign io_dma_cmd_payload_fragment_mask = ioDma_cmd_payload_fragment_mask;
  assign ioDma_rsp_valid = io_dma_rsp_valid;
  assign io_dma_rsp_ready = ioDma_rsp_ready;
  assign ioDma_rsp_payload_last = io_dma_rsp_payload_last;
  assign ioDma_rsp_payload_fragment_opcode = io_dma_rsp_payload_fragment_opcode;
  assign ioDma_rsp_payload_fragment_data = io_dma_rsp_payload_fragment_data;
  always @(*) begin
    ioDma_cmd_valid = 1'b0;
    case(sof_stateReg)
      sof_enumDef_FRAME_TX : begin
      end
      sof_enumDef_FRAME_NUMBER_CMD : begin
        ioDma_cmd_valid = 1'b1;
      end
      sof_enumDef_FRAME_NUMBER_RSP : begin
      end
      default : begin
      end
    endcase
    case(endpoint_stateReg)
      endpoint_enumDef_ED_READ_CMD : begin
        ioDma_cmd_valid = 1'b1;
      end
      endpoint_enumDef_ED_READ_RSP : begin
      end
      endpoint_enumDef_ED_ANALYSE : begin
      end
      endpoint_enumDef_TD_READ_CMD : begin
        ioDma_cmd_valid = 1'b1;
      end
      endpoint_enumDef_TD_READ_RSP : begin
      end
      endpoint_enumDef_TD_READ_DELAY : begin
      end
      endpoint_enumDef_TD_ANALYSE : begin
      end
      endpoint_enumDef_TD_CHECK_TIME : begin
      end
      endpoint_enumDef_BUFFER_READ : begin
      end
      endpoint_enumDef_TOKEN : begin
      end
      endpoint_enumDef_DATA_TX : begin
      end
      endpoint_enumDef_DATA_RX : begin
      end
      endpoint_enumDef_DATA_RX_VALIDATE : begin
      end
      endpoint_enumDef_ACK_RX : begin
      end
      endpoint_enumDef_ACK_TX_0 : begin
      end
      endpoint_enumDef_ACK_TX_1 : begin
      end
      endpoint_enumDef_ACK_TX_EOP : begin
      end
      endpoint_enumDef_DATA_RX_WAIT_DMA : begin
      end
      endpoint_enumDef_UPDATE_TD_PROCESS : begin
      end
      endpoint_enumDef_UPDATE_TD_CMD : begin
        ioDma_cmd_valid = 1'b1;
      end
      endpoint_enumDef_UPDATE_ED_CMD : begin
        ioDma_cmd_valid = 1'b1;
      end
      endpoint_enumDef_UPDATE_SYNC : begin
      end
      endpoint_enumDef_ABORD : begin
      end
      default : begin
      end
    endcase
    case(endpoint_dmaLogic_stateReg)
      endpoint_dmaLogic_enumDef_INIT : begin
      end
      endpoint_dmaLogic_enumDef_TO_USB : begin
      end
      endpoint_dmaLogic_enumDef_FROM_USB : begin
      end
      endpoint_dmaLogic_enumDef_VALIDATION : begin
      end
      endpoint_dmaLogic_enumDef_CALC_CMD : begin
      end
      endpoint_dmaLogic_enumDef_READ_CMD : begin
        ioDma_cmd_valid = 1'b1;
      end
      endpoint_dmaLogic_enumDef_WRITE_CMD : begin
        ioDma_cmd_valid = endpoint_dmaLogic_storage_readRsp_valid;
      end
      default : begin
      end
    endcase
    case(operational_stateReg)
      operational_enumDef_SOF : begin
      end
      operational_enumDef_ARBITER : begin
      end
      operational_enumDef_END_POINT : begin
      end
      operational_enumDef_PERIODIC_HEAD_CMD : begin
        ioDma_cmd_valid = 1'b1;
      end
      operational_enumDef_PERIODIC_HEAD_RSP : begin
      end
      operational_enumDef_WAIT_SOF : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    ioDma_cmd_payload_last = 1'bx;
    case(sof_stateReg)
      sof_enumDef_FRAME_TX : begin
      end
      sof_enumDef_FRAME_NUMBER_CMD : begin
        ioDma_cmd_payload_last = (dmaWriteCtx_counter == 4'b0001);
      end
      sof_enumDef_FRAME_NUMBER_RSP : begin
      end
      default : begin
      end
    endcase
    case(endpoint_stateReg)
      endpoint_enumDef_ED_READ_CMD : begin
        ioDma_cmd_payload_last = 1'b1;
      end
      endpoint_enumDef_ED_READ_RSP : begin
      end
      endpoint_enumDef_ED_ANALYSE : begin
      end
      endpoint_enumDef_TD_READ_CMD : begin
        ioDma_cmd_payload_last = 1'b1;
      end
      endpoint_enumDef_TD_READ_RSP : begin
      end
      endpoint_enumDef_TD_READ_DELAY : begin
      end
      endpoint_enumDef_TD_ANALYSE : begin
      end
      endpoint_enumDef_TD_CHECK_TIME : begin
      end
      endpoint_enumDef_BUFFER_READ : begin
      end
      endpoint_enumDef_TOKEN : begin
      end
      endpoint_enumDef_DATA_TX : begin
      end
      endpoint_enumDef_DATA_RX : begin
      end
      endpoint_enumDef_DATA_RX_VALIDATE : begin
      end
      endpoint_enumDef_ACK_RX : begin
      end
      endpoint_enumDef_ACK_TX_0 : begin
      end
      endpoint_enumDef_ACK_TX_1 : begin
      end
      endpoint_enumDef_ACK_TX_EOP : begin
      end
      endpoint_enumDef_DATA_RX_WAIT_DMA : begin
      end
      endpoint_enumDef_UPDATE_TD_PROCESS : begin
      end
      endpoint_enumDef_UPDATE_TD_CMD : begin
        ioDma_cmd_payload_last = (dmaWriteCtx_counter == _zz_ioDma_cmd_payload_last);
      end
      endpoint_enumDef_UPDATE_ED_CMD : begin
        ioDma_cmd_payload_last = (dmaWriteCtx_counter == 4'b0011);
      end
      endpoint_enumDef_UPDATE_SYNC : begin
      end
      endpoint_enumDef_ABORD : begin
      end
      default : begin
      end
    endcase
    case(endpoint_dmaLogic_stateReg)
      endpoint_dmaLogic_enumDef_INIT : begin
      end
      endpoint_dmaLogic_enumDef_TO_USB : begin
      end
      endpoint_dmaLogic_enumDef_FROM_USB : begin
      end
      endpoint_dmaLogic_enumDef_VALIDATION : begin
      end
      endpoint_dmaLogic_enumDef_CALC_CMD : begin
      end
      endpoint_dmaLogic_enumDef_READ_CMD : begin
        ioDma_cmd_payload_last = 1'b1;
      end
      endpoint_dmaLogic_enumDef_WRITE_CMD : begin
        ioDma_cmd_payload_last = endpoint_dmaLogic_beatLast;
      end
      default : begin
      end
    endcase
    case(operational_stateReg)
      operational_enumDef_SOF : begin
      end
      operational_enumDef_ARBITER : begin
      end
      operational_enumDef_END_POINT : begin
      end
      operational_enumDef_PERIODIC_HEAD_CMD : begin
        ioDma_cmd_payload_last = 1'b1;
      end
      operational_enumDef_PERIODIC_HEAD_RSP : begin
      end
      operational_enumDef_WAIT_SOF : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    ioDma_cmd_payload_fragment_opcode = 1'bx;
    case(sof_stateReg)
      sof_enumDef_FRAME_TX : begin
      end
      sof_enumDef_FRAME_NUMBER_CMD : begin
        ioDma_cmd_payload_fragment_opcode = 1'b1;
      end
      sof_enumDef_FRAME_NUMBER_RSP : begin
      end
      default : begin
      end
    endcase
    case(endpoint_stateReg)
      endpoint_enumDef_ED_READ_CMD : begin
        ioDma_cmd_payload_fragment_opcode = 1'b0;
      end
      endpoint_enumDef_ED_READ_RSP : begin
      end
      endpoint_enumDef_ED_ANALYSE : begin
      end
      endpoint_enumDef_TD_READ_CMD : begin
        ioDma_cmd_payload_fragment_opcode = 1'b0;
      end
      endpoint_enumDef_TD_READ_RSP : begin
      end
      endpoint_enumDef_TD_READ_DELAY : begin
      end
      endpoint_enumDef_TD_ANALYSE : begin
      end
      endpoint_enumDef_TD_CHECK_TIME : begin
      end
      endpoint_enumDef_BUFFER_READ : begin
      end
      endpoint_enumDef_TOKEN : begin
      end
      endpoint_enumDef_DATA_TX : begin
      end
      endpoint_enumDef_DATA_RX : begin
      end
      endpoint_enumDef_DATA_RX_VALIDATE : begin
      end
      endpoint_enumDef_ACK_RX : begin
      end
      endpoint_enumDef_ACK_TX_0 : begin
      end
      endpoint_enumDef_ACK_TX_1 : begin
      end
      endpoint_enumDef_ACK_TX_EOP : begin
      end
      endpoint_enumDef_DATA_RX_WAIT_DMA : begin
      end
      endpoint_enumDef_UPDATE_TD_PROCESS : begin
      end
      endpoint_enumDef_UPDATE_TD_CMD : begin
        ioDma_cmd_payload_fragment_opcode = 1'b1;
      end
      endpoint_enumDef_UPDATE_ED_CMD : begin
        ioDma_cmd_payload_fragment_opcode = 1'b1;
      end
      endpoint_enumDef_UPDATE_SYNC : begin
      end
      endpoint_enumDef_ABORD : begin
      end
      default : begin
      end
    endcase
    case(endpoint_dmaLogic_stateReg)
      endpoint_dmaLogic_enumDef_INIT : begin
      end
      endpoint_dmaLogic_enumDef_TO_USB : begin
      end
      endpoint_dmaLogic_enumDef_FROM_USB : begin
      end
      endpoint_dmaLogic_enumDef_VALIDATION : begin
      end
      endpoint_dmaLogic_enumDef_CALC_CMD : begin
      end
      endpoint_dmaLogic_enumDef_READ_CMD : begin
        ioDma_cmd_payload_fragment_opcode = 1'b0;
      end
      endpoint_dmaLogic_enumDef_WRITE_CMD : begin
        ioDma_cmd_payload_fragment_opcode = 1'b1;
      end
      default : begin
      end
    endcase
    case(operational_stateReg)
      operational_enumDef_SOF : begin
      end
      operational_enumDef_ARBITER : begin
      end
      operational_enumDef_END_POINT : begin
      end
      operational_enumDef_PERIODIC_HEAD_CMD : begin
        ioDma_cmd_payload_fragment_opcode = 1'b0;
      end
      operational_enumDef_PERIODIC_HEAD_RSP : begin
      end
      operational_enumDef_WAIT_SOF : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    ioDma_cmd_payload_fragment_address = 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
    case(sof_stateReg)
      sof_enumDef_FRAME_TX : begin
      end
      sof_enumDef_FRAME_NUMBER_CMD : begin
        ioDma_cmd_payload_fragment_address = (reg_hcHCCA_HCCA_address | 32'h00000080);
      end
      sof_enumDef_FRAME_NUMBER_RSP : begin
      end
      default : begin
      end
    endcase
    case(endpoint_stateReg)
      endpoint_enumDef_ED_READ_CMD : begin
        ioDma_cmd_payload_fragment_address = endpoint_ED_address;
      end
      endpoint_enumDef_ED_READ_RSP : begin
      end
      endpoint_enumDef_ED_ANALYSE : begin
      end
      endpoint_enumDef_TD_READ_CMD : begin
        ioDma_cmd_payload_fragment_address = endpoint_TD_address;
      end
      endpoint_enumDef_TD_READ_RSP : begin
      end
      endpoint_enumDef_TD_READ_DELAY : begin
      end
      endpoint_enumDef_TD_ANALYSE : begin
      end
      endpoint_enumDef_TD_CHECK_TIME : begin
      end
      endpoint_enumDef_BUFFER_READ : begin
      end
      endpoint_enumDef_TOKEN : begin
      end
      endpoint_enumDef_DATA_TX : begin
      end
      endpoint_enumDef_DATA_RX : begin
      end
      endpoint_enumDef_DATA_RX_VALIDATE : begin
      end
      endpoint_enumDef_ACK_RX : begin
      end
      endpoint_enumDef_ACK_TX_0 : begin
      end
      endpoint_enumDef_ACK_TX_1 : begin
      end
      endpoint_enumDef_ACK_TX_EOP : begin
      end
      endpoint_enumDef_DATA_RX_WAIT_DMA : begin
      end
      endpoint_enumDef_UPDATE_TD_PROCESS : begin
      end
      endpoint_enumDef_UPDATE_TD_CMD : begin
        ioDma_cmd_payload_fragment_address = endpoint_TD_address;
      end
      endpoint_enumDef_UPDATE_ED_CMD : begin
        ioDma_cmd_payload_fragment_address = endpoint_ED_address;
      end
      endpoint_enumDef_UPDATE_SYNC : begin
      end
      endpoint_enumDef_ABORD : begin
      end
      default : begin
      end
    endcase
    case(endpoint_dmaLogic_stateReg)
      endpoint_dmaLogic_enumDef_INIT : begin
      end
      endpoint_dmaLogic_enumDef_TO_USB : begin
      end
      endpoint_dmaLogic_enumDef_FROM_USB : begin
      end
      endpoint_dmaLogic_enumDef_VALIDATION : begin
      end
      endpoint_dmaLogic_enumDef_CALC_CMD : begin
      end
      endpoint_dmaLogic_enumDef_READ_CMD : begin
        ioDma_cmd_payload_fragment_address = endpoint_currentAddressBmb;
      end
      endpoint_dmaLogic_enumDef_WRITE_CMD : begin
        ioDma_cmd_payload_fragment_address = endpoint_currentAddressBmb;
      end
      default : begin
      end
    endcase
    case(operational_stateReg)
      operational_enumDef_SOF : begin
      end
      operational_enumDef_ARBITER : begin
      end
      operational_enumDef_END_POINT : begin
      end
      operational_enumDef_PERIODIC_HEAD_CMD : begin
        ioDma_cmd_payload_fragment_address = (reg_hcHCCA_HCCA_address | _zz_ioDma_cmd_payload_fragment_address);
      end
      operational_enumDef_PERIODIC_HEAD_RSP : begin
      end
      operational_enumDef_WAIT_SOF : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    ioDma_cmd_payload_fragment_length = 6'bxxxxxx;
    case(sof_stateReg)
      sof_enumDef_FRAME_TX : begin
      end
      sof_enumDef_FRAME_NUMBER_CMD : begin
        ioDma_cmd_payload_fragment_length = 6'h07;
      end
      sof_enumDef_FRAME_NUMBER_RSP : begin
      end
      default : begin
      end
    endcase
    case(endpoint_stateReg)
      endpoint_enumDef_ED_READ_CMD : begin
        ioDma_cmd_payload_fragment_length = 6'h0f;
      end
      endpoint_enumDef_ED_READ_RSP : begin
      end
      endpoint_enumDef_ED_ANALYSE : begin
      end
      endpoint_enumDef_TD_READ_CMD : begin
        ioDma_cmd_payload_fragment_length = {1'd0, _zz_ioDma_cmd_payload_fragment_length};
      end
      endpoint_enumDef_TD_READ_RSP : begin
      end
      endpoint_enumDef_TD_READ_DELAY : begin
      end
      endpoint_enumDef_TD_ANALYSE : begin
      end
      endpoint_enumDef_TD_CHECK_TIME : begin
      end
      endpoint_enumDef_BUFFER_READ : begin
      end
      endpoint_enumDef_TOKEN : begin
      end
      endpoint_enumDef_DATA_TX : begin
      end
      endpoint_enumDef_DATA_RX : begin
      end
      endpoint_enumDef_DATA_RX_VALIDATE : begin
      end
      endpoint_enumDef_ACK_RX : begin
      end
      endpoint_enumDef_ACK_TX_0 : begin
      end
      endpoint_enumDef_ACK_TX_1 : begin
      end
      endpoint_enumDef_ACK_TX_EOP : begin
      end
      endpoint_enumDef_DATA_RX_WAIT_DMA : begin
      end
      endpoint_enumDef_UPDATE_TD_PROCESS : begin
      end
      endpoint_enumDef_UPDATE_TD_CMD : begin
        ioDma_cmd_payload_fragment_length = {1'd0, _zz_ioDma_cmd_payload_fragment_length_1};
      end
      endpoint_enumDef_UPDATE_ED_CMD : begin
        ioDma_cmd_payload_fragment_length = 6'h0f;
      end
      endpoint_enumDef_UPDATE_SYNC : begin
      end
      endpoint_enumDef_ABORD : begin
      end
      default : begin
      end
    endcase
    case(endpoint_dmaLogic_stateReg)
      endpoint_dmaLogic_enumDef_INIT : begin
      end
      endpoint_dmaLogic_enumDef_TO_USB : begin
      end
      endpoint_dmaLogic_enumDef_FROM_USB : begin
      end
      endpoint_dmaLogic_enumDef_VALIDATION : begin
      end
      endpoint_dmaLogic_enumDef_CALC_CMD : begin
      end
      endpoint_dmaLogic_enumDef_READ_CMD : begin
        ioDma_cmd_payload_fragment_length = 6'h3f;
      end
      endpoint_dmaLogic_enumDef_WRITE_CMD : begin
        ioDma_cmd_payload_fragment_length = 6'h3f;
      end
      default : begin
      end
    endcase
    case(operational_stateReg)
      operational_enumDef_SOF : begin
      end
      operational_enumDef_ARBITER : begin
      end
      operational_enumDef_END_POINT : begin
      end
      operational_enumDef_PERIODIC_HEAD_CMD : begin
        ioDma_cmd_payload_fragment_length = 6'h03;
      end
      operational_enumDef_PERIODIC_HEAD_RSP : begin
      end
      operational_enumDef_WAIT_SOF : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    ioDma_cmd_payload_fragment_data = 32'h0;
    case(sof_stateReg)
      sof_enumDef_FRAME_TX : begin
      end
      sof_enumDef_FRAME_NUMBER_CMD : begin
        if(when_UsbOhci_l207) begin
          ioDma_cmd_payload_fragment_data[31 : 0] = {16'h0,reg_hcFmNumber_FN};
        end
        if(sof_doInterruptDelay) begin
          if(when_UsbOhci_l207_1) begin
            ioDma_cmd_payload_fragment_data[31 : 0] = {reg_hcDoneHead_DH_address[31 : 1],reg_hcInterrupt_unmaskedPending};
          end
        end
      end
      sof_enumDef_FRAME_NUMBER_RSP : begin
      end
      default : begin
      end
    endcase
    case(endpoint_stateReg)
      endpoint_enumDef_ED_READ_CMD : begin
      end
      endpoint_enumDef_ED_READ_RSP : begin
      end
      endpoint_enumDef_ED_ANALYSE : begin
      end
      endpoint_enumDef_TD_READ_CMD : begin
      end
      endpoint_enumDef_TD_READ_RSP : begin
      end
      endpoint_enumDef_TD_READ_DELAY : begin
      end
      endpoint_enumDef_TD_ANALYSE : begin
      end
      endpoint_enumDef_TD_CHECK_TIME : begin
      end
      endpoint_enumDef_BUFFER_READ : begin
      end
      endpoint_enumDef_TOKEN : begin
      end
      endpoint_enumDef_DATA_TX : begin
      end
      endpoint_enumDef_DATA_RX : begin
      end
      endpoint_enumDef_DATA_RX_VALIDATE : begin
      end
      endpoint_enumDef_ACK_RX : begin
      end
      endpoint_enumDef_ACK_TX_0 : begin
      end
      endpoint_enumDef_ACK_TX_1 : begin
      end
      endpoint_enumDef_ACK_TX_EOP : begin
      end
      endpoint_enumDef_DATA_RX_WAIT_DMA : begin
      end
      endpoint_enumDef_UPDATE_TD_PROCESS : begin
      end
      endpoint_enumDef_UPDATE_TD_CMD : begin
        if(endpoint_ED_F) begin
          if(endpoint_TD_isoOverrunReg) begin
            if(when_UsbOhci_l207_2) begin
              ioDma_cmd_payload_fragment_data[31 : 24] = {{4'b1000,endpoint_TD_words_0[27]},endpoint_TD_FC};
            end
          end else begin
            if(endpoint_TD_isoLastReg) begin
              if(when_UsbOhci_l207_3) begin
                ioDma_cmd_payload_fragment_data[31 : 24] = {{4'b0000,endpoint_TD_words_0[27]},endpoint_TD_FC};
              end
            end
            if(when_UsbOhci_l1433) begin
              if(when_UsbOhci_l207_4) begin
                ioDma_cmd_payload_fragment_data[15 : 0] = _zz_ioDma_cmd_payload_fragment_data;
              end
            end
            if(when_UsbOhci_l1433_1) begin
              if(when_UsbOhci_l207_5) begin
                ioDma_cmd_payload_fragment_data[31 : 16] = _zz_ioDma_cmd_payload_fragment_data;
              end
            end
            if(when_UsbOhci_l1433_2) begin
              if(when_UsbOhci_l207_6) begin
                ioDma_cmd_payload_fragment_data[15 : 0] = _zz_ioDma_cmd_payload_fragment_data;
              end
            end
            if(when_UsbOhci_l1433_3) begin
              if(when_UsbOhci_l207_7) begin
                ioDma_cmd_payload_fragment_data[31 : 16] = _zz_ioDma_cmd_payload_fragment_data;
              end
            end
            if(when_UsbOhci_l1433_4) begin
              if(when_UsbOhci_l207_8) begin
                ioDma_cmd_payload_fragment_data[15 : 0] = _zz_ioDma_cmd_payload_fragment_data;
              end
            end
            if(when_UsbOhci_l1433_5) begin
              if(when_UsbOhci_l207_9) begin
                ioDma_cmd_payload_fragment_data[31 : 16] = _zz_ioDma_cmd_payload_fragment_data;
              end
            end
            if(when_UsbOhci_l1433_6) begin
              if(when_UsbOhci_l207_10) begin
                ioDma_cmd_payload_fragment_data[15 : 0] = _zz_ioDma_cmd_payload_fragment_data;
              end
            end
            if(when_UsbOhci_l1433_7) begin
              if(when_UsbOhci_l207_11) begin
                ioDma_cmd_payload_fragment_data[31 : 16] = _zz_ioDma_cmd_payload_fragment_data;
              end
            end
          end
        end else begin
          if(when_UsbOhci_l207_12) begin
            ioDma_cmd_payload_fragment_data[31 : 24] = {{endpoint_TD_CC,endpoint_TD_EC},endpoint_TD_TNext};
          end
          if(endpoint_TD_upateCBP) begin
            if(when_UsbOhci_l207_13) begin
              ioDma_cmd_payload_fragment_data[31 : 0] = endpoint_tdUpdateAddress;
            end
          end
        end
        if(endpoint_TD_retire) begin
          if(when_UsbOhci_l207_14) begin
            ioDma_cmd_payload_fragment_data[31 : 0] = reg_hcDoneHead_DH_address;
          end
        end
      end
      endpoint_enumDef_UPDATE_ED_CMD : begin
        if(endpoint_TD_retire) begin
          if(when_UsbOhci_l207_15) begin
            ioDma_cmd_payload_fragment_data[31 : 0] = {{{endpoint_TD_nextTD,2'b00},endpoint_TD_dataPhaseNext},endpoint_ED_H};
          end
        end
      end
      endpoint_enumDef_UPDATE_SYNC : begin
      end
      endpoint_enumDef_ABORD : begin
      end
      default : begin
      end
    endcase
    case(endpoint_dmaLogic_stateReg)
      endpoint_dmaLogic_enumDef_INIT : begin
      end
      endpoint_dmaLogic_enumDef_TO_USB : begin
      end
      endpoint_dmaLogic_enumDef_FROM_USB : begin
      end
      endpoint_dmaLogic_enumDef_VALIDATION : begin
      end
      endpoint_dmaLogic_enumDef_CALC_CMD : begin
      end
      endpoint_dmaLogic_enumDef_READ_CMD : begin
      end
      endpoint_dmaLogic_enumDef_WRITE_CMD : begin
        ioDma_cmd_payload_fragment_data = endpoint_dmaLogic_storage_readRsp_payload;
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    ioDma_cmd_payload_fragment_mask = 4'b0000;
    case(sof_stateReg)
      sof_enumDef_FRAME_TX : begin
      end
      sof_enumDef_FRAME_NUMBER_CMD : begin
        if(when_UsbOhci_l207) begin
          ioDma_cmd_payload_fragment_mask[3 : 0] = 4'b1111;
        end
        if(sof_doInterruptDelay) begin
          if(when_UsbOhci_l207_1) begin
            ioDma_cmd_payload_fragment_mask[3 : 0] = 4'b1111;
          end
        end
      end
      sof_enumDef_FRAME_NUMBER_RSP : begin
      end
      default : begin
      end
    endcase
    case(endpoint_stateReg)
      endpoint_enumDef_ED_READ_CMD : begin
      end
      endpoint_enumDef_ED_READ_RSP : begin
      end
      endpoint_enumDef_ED_ANALYSE : begin
      end
      endpoint_enumDef_TD_READ_CMD : begin
      end
      endpoint_enumDef_TD_READ_RSP : begin
      end
      endpoint_enumDef_TD_READ_DELAY : begin
      end
      endpoint_enumDef_TD_ANALYSE : begin
      end
      endpoint_enumDef_TD_CHECK_TIME : begin
      end
      endpoint_enumDef_BUFFER_READ : begin
      end
      endpoint_enumDef_TOKEN : begin
      end
      endpoint_enumDef_DATA_TX : begin
      end
      endpoint_enumDef_DATA_RX : begin
      end
      endpoint_enumDef_DATA_RX_VALIDATE : begin
      end
      endpoint_enumDef_ACK_RX : begin
      end
      endpoint_enumDef_ACK_TX_0 : begin
      end
      endpoint_enumDef_ACK_TX_1 : begin
      end
      endpoint_enumDef_ACK_TX_EOP : begin
      end
      endpoint_enumDef_DATA_RX_WAIT_DMA : begin
      end
      endpoint_enumDef_UPDATE_TD_PROCESS : begin
      end
      endpoint_enumDef_UPDATE_TD_CMD : begin
        if(endpoint_ED_F) begin
          if(endpoint_TD_isoOverrunReg) begin
            if(when_UsbOhci_l207_2) begin
              ioDma_cmd_payload_fragment_mask[3 : 3] = 1'b1;
            end
          end else begin
            if(endpoint_TD_isoLastReg) begin
              if(when_UsbOhci_l207_3) begin
                ioDma_cmd_payload_fragment_mask[3 : 3] = 1'b1;
              end
            end
            if(when_UsbOhci_l1433) begin
              if(when_UsbOhci_l207_4) begin
                ioDma_cmd_payload_fragment_mask[1 : 0] = 2'b11;
              end
            end
            if(when_UsbOhci_l1433_1) begin
              if(when_UsbOhci_l207_5) begin
                ioDma_cmd_payload_fragment_mask[3 : 2] = 2'b11;
              end
            end
            if(when_UsbOhci_l1433_2) begin
              if(when_UsbOhci_l207_6) begin
                ioDma_cmd_payload_fragment_mask[1 : 0] = 2'b11;
              end
            end
            if(when_UsbOhci_l1433_3) begin
              if(when_UsbOhci_l207_7) begin
                ioDma_cmd_payload_fragment_mask[3 : 2] = 2'b11;
              end
            end
            if(when_UsbOhci_l1433_4) begin
              if(when_UsbOhci_l207_8) begin
                ioDma_cmd_payload_fragment_mask[1 : 0] = 2'b11;
              end
            end
            if(when_UsbOhci_l1433_5) begin
              if(when_UsbOhci_l207_9) begin
                ioDma_cmd_payload_fragment_mask[3 : 2] = 2'b11;
              end
            end
            if(when_UsbOhci_l1433_6) begin
              if(when_UsbOhci_l207_10) begin
                ioDma_cmd_payload_fragment_mask[1 : 0] = 2'b11;
              end
            end
            if(when_UsbOhci_l1433_7) begin
              if(when_UsbOhci_l207_11) begin
                ioDma_cmd_payload_fragment_mask[3 : 2] = 2'b11;
              end
            end
          end
        end else begin
          if(when_UsbOhci_l207_12) begin
            ioDma_cmd_payload_fragment_mask[3 : 3] = 1'b1;
          end
          if(endpoint_TD_upateCBP) begin
            if(when_UsbOhci_l207_13) begin
              ioDma_cmd_payload_fragment_mask[3 : 0] = 4'b1111;
            end
          end
        end
        if(endpoint_TD_retire) begin
          if(when_UsbOhci_l207_14) begin
            ioDma_cmd_payload_fragment_mask[3 : 0] = 4'b1111;
          end
        end
      end
      endpoint_enumDef_UPDATE_ED_CMD : begin
        if(endpoint_TD_retire) begin
          if(when_UsbOhci_l207_15) begin
            ioDma_cmd_payload_fragment_mask[3 : 0] = 4'b1111;
          end
        end
      end
      endpoint_enumDef_UPDATE_SYNC : begin
      end
      endpoint_enumDef_ABORD : begin
      end
      default : begin
      end
    endcase
    case(endpoint_dmaLogic_stateReg)
      endpoint_dmaLogic_enumDef_INIT : begin
      end
      endpoint_dmaLogic_enumDef_TO_USB : begin
      end
      endpoint_dmaLogic_enumDef_FROM_USB : begin
      end
      endpoint_dmaLogic_enumDef_VALIDATION : begin
      end
      endpoint_dmaLogic_enumDef_CALC_CMD : begin
      end
      endpoint_dmaLogic_enumDef_READ_CMD : begin
      end
      endpoint_dmaLogic_enumDef_WRITE_CMD : begin
        ioDma_cmd_payload_fragment_mask = ((((! endpoint_dmaLogic_headHit) ? 4'b1111 : endpoint_dmaLogic_headMask) & ((! endpoint_dmaLogic_lastHit) ? 4'b1111 : endpoint_dmaLogic_lastMask)) & ((endpoint_dmaLogic_headHit || endpoint_dmaLogic_inBurst) ? 4'b1111 : 4'b0000));
      end
      default : begin
      end
    endcase
  end

  assign ioDma_rsp_ready = 1'b1;
  assign dmaRspMux_vec_0 = ioDma_rsp_payload_fragment_data[31 : 0];
  assign dmaRspMux_data = dmaRspMux_vec_0;
  always @(*) begin
    io_phy_tx_valid = 1'b0;
    case(token_stateReg)
      token_enumDef_INIT : begin
      end
      token_enumDef_PID : begin
        io_phy_tx_valid = 1'b1;
      end
      token_enumDef_B1 : begin
        io_phy_tx_valid = 1'b1;
      end
      token_enumDef_B2 : begin
        io_phy_tx_valid = 1'b1;
      end
      token_enumDef_EOP : begin
      end
      default : begin
      end
    endcase
    case(dataTx_stateReg)
      dataTx_enumDef_PID : begin
        io_phy_tx_valid = 1'b1;
      end
      dataTx_enumDef_DATA : begin
        io_phy_tx_valid = 1'b1;
      end
      dataTx_enumDef_CRC_0 : begin
        io_phy_tx_valid = 1'b1;
      end
      dataTx_enumDef_CRC_1 : begin
        io_phy_tx_valid = 1'b1;
      end
      dataTx_enumDef_EOP : begin
      end
      default : begin
      end
    endcase
    case(endpoint_stateReg)
      endpoint_enumDef_ED_READ_CMD : begin
      end
      endpoint_enumDef_ED_READ_RSP : begin
      end
      endpoint_enumDef_ED_ANALYSE : begin
      end
      endpoint_enumDef_TD_READ_CMD : begin
      end
      endpoint_enumDef_TD_READ_RSP : begin
      end
      endpoint_enumDef_TD_READ_DELAY : begin
      end
      endpoint_enumDef_TD_ANALYSE : begin
      end
      endpoint_enumDef_TD_CHECK_TIME : begin
      end
      endpoint_enumDef_BUFFER_READ : begin
      end
      endpoint_enumDef_TOKEN : begin
      end
      endpoint_enumDef_DATA_TX : begin
      end
      endpoint_enumDef_DATA_RX : begin
      end
      endpoint_enumDef_DATA_RX_VALIDATE : begin
      end
      endpoint_enumDef_ACK_RX : begin
      end
      endpoint_enumDef_ACK_TX_0 : begin
      end
      endpoint_enumDef_ACK_TX_1 : begin
        io_phy_tx_valid = 1'b1;
      end
      endpoint_enumDef_ACK_TX_EOP : begin
      end
      endpoint_enumDef_DATA_RX_WAIT_DMA : begin
      end
      endpoint_enumDef_UPDATE_TD_PROCESS : begin
      end
      endpoint_enumDef_UPDATE_TD_CMD : begin
      end
      endpoint_enumDef_UPDATE_ED_CMD : begin
      end
      endpoint_enumDef_UPDATE_SYNC : begin
      end
      endpoint_enumDef_ABORD : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    io_phy_tx_payload_fragment = 8'bxxxxxxxx;
    case(token_stateReg)
      token_enumDef_INIT : begin
      end
      token_enumDef_PID : begin
        io_phy_tx_payload_fragment = {(~ token_pid),token_pid};
      end
      token_enumDef_B1 : begin
        io_phy_tx_payload_fragment = token_data[7 : 0];
      end
      token_enumDef_B2 : begin
        io_phy_tx_payload_fragment = {token_crc5_io_result,token_data[10 : 8]};
      end
      token_enumDef_EOP : begin
      end
      default : begin
      end
    endcase
    case(dataTx_stateReg)
      dataTx_enumDef_PID : begin
        io_phy_tx_payload_fragment = {(~ dataTx_pid),dataTx_pid};
      end
      dataTx_enumDef_DATA : begin
        io_phy_tx_payload_fragment = dataTx_data_payload_fragment;
      end
      dataTx_enumDef_CRC_0 : begin
        io_phy_tx_payload_fragment = dataTx_crc16_io_result[7 : 0];
      end
      dataTx_enumDef_CRC_1 : begin
        io_phy_tx_payload_fragment = dataTx_crc16_io_result[15 : 8];
      end
      dataTx_enumDef_EOP : begin
      end
      default : begin
      end
    endcase
    case(endpoint_stateReg)
      endpoint_enumDef_ED_READ_CMD : begin
      end
      endpoint_enumDef_ED_READ_RSP : begin
      end
      endpoint_enumDef_ED_ANALYSE : begin
      end
      endpoint_enumDef_TD_READ_CMD : begin
      end
      endpoint_enumDef_TD_READ_RSP : begin
      end
      endpoint_enumDef_TD_READ_DELAY : begin
      end
      endpoint_enumDef_TD_ANALYSE : begin
      end
      endpoint_enumDef_TD_CHECK_TIME : begin
      end
      endpoint_enumDef_BUFFER_READ : begin
      end
      endpoint_enumDef_TOKEN : begin
      end
      endpoint_enumDef_DATA_TX : begin
      end
      endpoint_enumDef_DATA_RX : begin
      end
      endpoint_enumDef_DATA_RX_VALIDATE : begin
      end
      endpoint_enumDef_ACK_RX : begin
      end
      endpoint_enumDef_ACK_TX_0 : begin
      end
      endpoint_enumDef_ACK_TX_1 : begin
        io_phy_tx_payload_fragment = 8'hd2;
      end
      endpoint_enumDef_ACK_TX_EOP : begin
      end
      endpoint_enumDef_DATA_RX_WAIT_DMA : begin
      end
      endpoint_enumDef_UPDATE_TD_PROCESS : begin
      end
      endpoint_enumDef_UPDATE_TD_CMD : begin
      end
      endpoint_enumDef_UPDATE_ED_CMD : begin
      end
      endpoint_enumDef_UPDATE_SYNC : begin
      end
      endpoint_enumDef_ABORD : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    io_phy_tx_payload_last = 1'bx;
    case(token_stateReg)
      token_enumDef_INIT : begin
      end
      token_enumDef_PID : begin
        io_phy_tx_payload_last = 1'b0;
      end
      token_enumDef_B1 : begin
        io_phy_tx_payload_last = 1'b0;
      end
      token_enumDef_B2 : begin
        io_phy_tx_payload_last = 1'b1;
      end
      token_enumDef_EOP : begin
      end
      default : begin
      end
    endcase
    case(dataTx_stateReg)
      dataTx_enumDef_PID : begin
        io_phy_tx_payload_last = 1'b0;
      end
      dataTx_enumDef_DATA : begin
        io_phy_tx_payload_last = 1'b0;
      end
      dataTx_enumDef_CRC_0 : begin
        io_phy_tx_payload_last = 1'b0;
      end
      dataTx_enumDef_CRC_1 : begin
        io_phy_tx_payload_last = 1'b1;
      end
      dataTx_enumDef_EOP : begin
      end
      default : begin
      end
    endcase
    case(endpoint_stateReg)
      endpoint_enumDef_ED_READ_CMD : begin
      end
      endpoint_enumDef_ED_READ_RSP : begin
      end
      endpoint_enumDef_ED_ANALYSE : begin
      end
      endpoint_enumDef_TD_READ_CMD : begin
      end
      endpoint_enumDef_TD_READ_RSP : begin
      end
      endpoint_enumDef_TD_READ_DELAY : begin
      end
      endpoint_enumDef_TD_ANALYSE : begin
      end
      endpoint_enumDef_TD_CHECK_TIME : begin
      end
      endpoint_enumDef_BUFFER_READ : begin
      end
      endpoint_enumDef_TOKEN : begin
      end
      endpoint_enumDef_DATA_TX : begin
      end
      endpoint_enumDef_DATA_RX : begin
      end
      endpoint_enumDef_DATA_RX_VALIDATE : begin
      end
      endpoint_enumDef_ACK_RX : begin
      end
      endpoint_enumDef_ACK_TX_0 : begin
      end
      endpoint_enumDef_ACK_TX_1 : begin
        io_phy_tx_payload_last = 1'b1;
      end
      endpoint_enumDef_ACK_TX_EOP : begin
      end
      endpoint_enumDef_DATA_RX_WAIT_DMA : begin
      end
      endpoint_enumDef_UPDATE_TD_PROCESS : begin
      end
      endpoint_enumDef_UPDATE_TD_CMD : begin
      end
      endpoint_enumDef_UPDATE_ED_CMD : begin
      end
      endpoint_enumDef_UPDATE_SYNC : begin
      end
      endpoint_enumDef_ABORD : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    ctrlHalt = 1'b0;
    case(hc_stateReg)
      hc_enumDef_RESET : begin
      end
      hc_enumDef_RESUME : begin
      end
      hc_enumDef_OPERATIONAL : begin
      end
      hc_enumDef_SUSPEND : begin
      end
      hc_enumDef_ANY_TO_RESET : begin
        ctrlHalt = 1'b1;
      end
      hc_enumDef_ANY_TO_SUSPEND : begin
        ctrlHalt = 1'b1;
      end
      default : begin
      end
    endcase
  end

  assign ctrl_readErrorFlag = 1'b0;
  assign ctrl_writeErrorFlag = 1'b0;
  assign ctrl_readHaltTrigger = 1'b0;
  always @(*) begin
    ctrl_writeHaltTrigger = 1'b0;
    if(ctrlHalt) begin
      ctrl_writeHaltTrigger = 1'b1;
    end
  end

  assign _zz_ctrl_rsp_ready = (! (ctrl_readHaltTrigger || ctrl_writeHaltTrigger));
  assign ctrl_rsp_ready = (_zz_ctrl_rsp_ready_1 && _zz_ctrl_rsp_ready);
  always @(*) begin
    _zz_ctrl_rsp_ready_1 = io_ctrl_rsp_ready;
    if(when_Stream_l393) begin
      _zz_ctrl_rsp_ready_1 = 1'b1;
    end
  end

  assign when_Stream_l393 = (! _zz_io_ctrl_rsp_valid);
  assign _zz_io_ctrl_rsp_valid = _zz_io_ctrl_rsp_valid_1;
  assign io_ctrl_rsp_valid = _zz_io_ctrl_rsp_valid;
  assign io_ctrl_rsp_payload_last = _zz_io_ctrl_rsp_payload_last;
  assign io_ctrl_rsp_payload_fragment_opcode = _zz_io_ctrl_rsp_payload_fragment_opcode;
  assign io_ctrl_rsp_payload_fragment_data = _zz_io_ctrl_rsp_payload_fragment_data;
  assign ctrl_askWrite = (io_ctrl_cmd_valid && (io_ctrl_cmd_payload_fragment_opcode == 1'b1));
  assign ctrl_askRead = (io_ctrl_cmd_valid && (io_ctrl_cmd_payload_fragment_opcode == 1'b0));
  assign io_ctrl_cmd_fire = (io_ctrl_cmd_valid && io_ctrl_cmd_ready);
  assign ctrl_doWrite = (io_ctrl_cmd_fire && (io_ctrl_cmd_payload_fragment_opcode == 1'b1));
  assign ctrl_doRead = (io_ctrl_cmd_fire && (io_ctrl_cmd_payload_fragment_opcode == 1'b0));
  assign ctrl_rsp_valid = io_ctrl_cmd_valid;
  assign io_ctrl_cmd_ready = ctrl_rsp_ready;
  assign ctrl_rsp_payload_last = 1'b1;
  assign when_BmbSlaveFactory_l33 = (ctrl_doWrite && ctrl_writeErrorFlag);
  always @(*) begin
    if(when_BmbSlaveFactory_l33) begin
      ctrl_rsp_payload_fragment_opcode = 1'b1;
    end else begin
      if(when_BmbSlaveFactory_l35) begin
        ctrl_rsp_payload_fragment_opcode = 1'b1;
      end else begin
        ctrl_rsp_payload_fragment_opcode = 1'b0;
      end
    end
  end

  assign when_BmbSlaveFactory_l35 = (ctrl_doRead && ctrl_readErrorFlag);
  always @(*) begin
    ctrl_rsp_payload_fragment_data = 32'h0;
    case(io_ctrl_cmd_payload_fragment_address)
      12'h0 : begin
        ctrl_rsp_payload_fragment_data[4 : 0] = reg_hcRevision_REV;
      end
      12'h004 : begin
        ctrl_rsp_payload_fragment_data[1 : 0] = reg_hcControl_CBSR;
        ctrl_rsp_payload_fragment_data[2 : 2] = reg_hcControl_PLE;
        ctrl_rsp_payload_fragment_data[3 : 3] = reg_hcControl_IE;
        ctrl_rsp_payload_fragment_data[4 : 4] = reg_hcControl_CLE;
        ctrl_rsp_payload_fragment_data[5 : 5] = reg_hcControl_BLE;
        ctrl_rsp_payload_fragment_data[7 : 6] = reg_hcControl_HCFS;
        ctrl_rsp_payload_fragment_data[8 : 8] = reg_hcControl_IR;
        ctrl_rsp_payload_fragment_data[9 : 9] = reg_hcControl_RWC;
        ctrl_rsp_payload_fragment_data[10 : 10] = reg_hcControl_RWE;
      end
      12'h008 : begin
        ctrl_rsp_payload_fragment_data[0 : 0] = doSoftReset;
        ctrl_rsp_payload_fragment_data[1 : 1] = reg_hcCommandStatus_CLF;
        ctrl_rsp_payload_fragment_data[2 : 2] = reg_hcCommandStatus_BLF;
        ctrl_rsp_payload_fragment_data[3 : 3] = reg_hcCommandStatus_OCR;
        ctrl_rsp_payload_fragment_data[17 : 16] = reg_hcCommandStatus_SOC;
      end
      12'h010 : begin
        ctrl_rsp_payload_fragment_data[31 : 31] = reg_hcInterrupt_MIE;
        ctrl_rsp_payload_fragment_data[0 : 0] = reg_hcInterrupt_SO_enable;
        ctrl_rsp_payload_fragment_data[1 : 1] = reg_hcInterrupt_WDH_enable;
        ctrl_rsp_payload_fragment_data[2 : 2] = reg_hcInterrupt_SF_enable;
        ctrl_rsp_payload_fragment_data[3 : 3] = reg_hcInterrupt_RD_enable;
        ctrl_rsp_payload_fragment_data[4 : 4] = reg_hcInterrupt_UE_enable;
        ctrl_rsp_payload_fragment_data[5 : 5] = reg_hcInterrupt_FNO_enable;
        ctrl_rsp_payload_fragment_data[6 : 6] = reg_hcInterrupt_RHSC_enable;
        ctrl_rsp_payload_fragment_data[30 : 30] = reg_hcInterrupt_OC_enable;
      end
      12'h014 : begin
        ctrl_rsp_payload_fragment_data[31 : 31] = reg_hcInterrupt_MIE;
        ctrl_rsp_payload_fragment_data[0 : 0] = reg_hcInterrupt_SO_enable;
        ctrl_rsp_payload_fragment_data[1 : 1] = reg_hcInterrupt_WDH_enable;
        ctrl_rsp_payload_fragment_data[2 : 2] = reg_hcInterrupt_SF_enable;
        ctrl_rsp_payload_fragment_data[3 : 3] = reg_hcInterrupt_RD_enable;
        ctrl_rsp_payload_fragment_data[4 : 4] = reg_hcInterrupt_UE_enable;
        ctrl_rsp_payload_fragment_data[5 : 5] = reg_hcInterrupt_FNO_enable;
        ctrl_rsp_payload_fragment_data[6 : 6] = reg_hcInterrupt_RHSC_enable;
        ctrl_rsp_payload_fragment_data[30 : 30] = reg_hcInterrupt_OC_enable;
      end
      12'h00c : begin
        ctrl_rsp_payload_fragment_data[0 : 0] = reg_hcInterrupt_SO_status;
        ctrl_rsp_payload_fragment_data[1 : 1] = reg_hcInterrupt_WDH_status;
        ctrl_rsp_payload_fragment_data[2 : 2] = reg_hcInterrupt_SF_status;
        ctrl_rsp_payload_fragment_data[3 : 3] = reg_hcInterrupt_RD_status;
        ctrl_rsp_payload_fragment_data[4 : 4] = reg_hcInterrupt_UE_status;
        ctrl_rsp_payload_fragment_data[5 : 5] = reg_hcInterrupt_FNO_status;
        ctrl_rsp_payload_fragment_data[6 : 6] = reg_hcInterrupt_RHSC_status;
        ctrl_rsp_payload_fragment_data[30 : 30] = reg_hcInterrupt_OC_status;
      end
      12'h018 : begin
        ctrl_rsp_payload_fragment_data[31 : 8] = reg_hcHCCA_HCCA_reg;
      end
      12'h01c : begin
        ctrl_rsp_payload_fragment_data[31 : 4] = reg_hcPeriodCurrentED_PCED_reg;
      end
      12'h020 : begin
        ctrl_rsp_payload_fragment_data[31 : 4] = reg_hcControlHeadED_CHED_reg;
      end
      12'h024 : begin
        ctrl_rsp_payload_fragment_data[31 : 4] = reg_hcControlCurrentED_CCED_reg;
      end
      12'h028 : begin
        ctrl_rsp_payload_fragment_data[31 : 4] = reg_hcBulkHeadED_BHED_reg;
      end
      12'h02c : begin
        ctrl_rsp_payload_fragment_data[31 : 4] = reg_hcBulkCurrentED_BCED_reg;
      end
      12'h030 : begin
        ctrl_rsp_payload_fragment_data[31 : 4] = reg_hcDoneHead_DH_reg;
      end
      12'h034 : begin
        ctrl_rsp_payload_fragment_data[13 : 0] = reg_hcFmInterval_FI;
        ctrl_rsp_payload_fragment_data[30 : 16] = reg_hcFmInterval_FSMPS;
        ctrl_rsp_payload_fragment_data[31 : 31] = reg_hcFmInterval_FIT;
      end
      12'h038 : begin
        ctrl_rsp_payload_fragment_data[13 : 0] = reg_hcFmRemaining_FR;
        ctrl_rsp_payload_fragment_data[31 : 31] = reg_hcFmRemaining_FRT;
      end
      12'h03c : begin
        ctrl_rsp_payload_fragment_data[15 : 0] = reg_hcFmNumber_FN;
      end
      12'h040 : begin
        ctrl_rsp_payload_fragment_data[13 : 0] = reg_hcPeriodicStart_PS;
      end
      12'h044 : begin
        ctrl_rsp_payload_fragment_data[11 : 0] = reg_hcLSThreshold_LST;
      end
      12'h048 : begin
        ctrl_rsp_payload_fragment_data[7 : 0] = reg_hcRhDescriptorA_NDP;
        ctrl_rsp_payload_fragment_data[8 : 8] = reg_hcRhDescriptorA_PSM;
        ctrl_rsp_payload_fragment_data[9 : 9] = reg_hcRhDescriptorA_NPS;
        ctrl_rsp_payload_fragment_data[11 : 11] = reg_hcRhDescriptorA_OCPM;
        ctrl_rsp_payload_fragment_data[12 : 12] = reg_hcRhDescriptorA_NOCP;
        ctrl_rsp_payload_fragment_data[31 : 24] = reg_hcRhDescriptorA_POTPGT;
      end
      12'h04c : begin
        ctrl_rsp_payload_fragment_data[2 : 1] = reg_hcRhDescriptorB_DR;
        ctrl_rsp_payload_fragment_data[18 : 17] = reg_hcRhDescriptorB_PPCM;
      end
      12'h050 : begin
        ctrl_rsp_payload_fragment_data[1 : 1] = io_phy_overcurrent;
        ctrl_rsp_payload_fragment_data[15 : 15] = reg_hcRhStatus_DRWE;
        ctrl_rsp_payload_fragment_data[17 : 17] = reg_hcRhStatus_CCIC;
      end
      12'h054 : begin
        ctrl_rsp_payload_fragment_data[2 : 2] = reg_hcRhPortStatus_0_PSS;
        ctrl_rsp_payload_fragment_data[8 : 8] = reg_hcRhPortStatus_0_PPS;
        ctrl_rsp_payload_fragment_data[0 : 0] = reg_hcRhPortStatus_0_CCS;
        ctrl_rsp_payload_fragment_data[1 : 1] = reg_hcRhPortStatus_0_PES;
        ctrl_rsp_payload_fragment_data[3 : 3] = io_phy_ports_0_overcurrent;
        ctrl_rsp_payload_fragment_data[4 : 4] = reg_hcRhPortStatus_0_reset;
        ctrl_rsp_payload_fragment_data[9 : 9] = io_phy_ports_0_lowSpeed;
        ctrl_rsp_payload_fragment_data[16 : 16] = reg_hcRhPortStatus_0_CSC_reg;
        ctrl_rsp_payload_fragment_data[17 : 17] = reg_hcRhPortStatus_0_PESC_reg;
        ctrl_rsp_payload_fragment_data[18 : 18] = reg_hcRhPortStatus_0_PSSC_reg;
        ctrl_rsp_payload_fragment_data[19 : 19] = reg_hcRhPortStatus_0_OCIC_reg;
        ctrl_rsp_payload_fragment_data[20 : 20] = reg_hcRhPortStatus_0_PRSC_reg;
      end
      12'h058 : begin
        ctrl_rsp_payload_fragment_data[2 : 2] = reg_hcRhPortStatus_1_PSS;
        ctrl_rsp_payload_fragment_data[8 : 8] = reg_hcRhPortStatus_1_PPS;
        ctrl_rsp_payload_fragment_data[0 : 0] = reg_hcRhPortStatus_1_CCS;
        ctrl_rsp_payload_fragment_data[1 : 1] = reg_hcRhPortStatus_1_PES;
        ctrl_rsp_payload_fragment_data[3 : 3] = io_phy_ports_1_overcurrent;
        ctrl_rsp_payload_fragment_data[4 : 4] = reg_hcRhPortStatus_1_reset;
        ctrl_rsp_payload_fragment_data[9 : 9] = io_phy_ports_1_lowSpeed;
        ctrl_rsp_payload_fragment_data[16 : 16] = reg_hcRhPortStatus_1_CSC_reg;
        ctrl_rsp_payload_fragment_data[17 : 17] = reg_hcRhPortStatus_1_PESC_reg;
        ctrl_rsp_payload_fragment_data[18 : 18] = reg_hcRhPortStatus_1_PSSC_reg;
        ctrl_rsp_payload_fragment_data[19 : 19] = reg_hcRhPortStatus_1_OCIC_reg;
        ctrl_rsp_payload_fragment_data[20 : 20] = reg_hcRhPortStatus_1_PRSC_reg;
      end
      default : begin
      end
    endcase
  end

  assign when_UsbOhci_l224 = (! doUnschedule);
  assign reg_hcRevision_REV = 5'h10;
  always @(*) begin
    reg_hcControl_HCFSWrite_valid = 1'b0;
    case(io_ctrl_cmd_payload_fragment_address)
      12'h004 : begin
        if(ctrl_doWrite) begin
          reg_hcControl_HCFSWrite_valid = 1'b1;
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    reg_hcCommandStatus_startSoftReset = 1'b0;
    if(when_BusSlaveFactory_l377) begin
      if(when_BusSlaveFactory_l379) begin
        reg_hcCommandStatus_startSoftReset = _zz_reg_hcCommandStatus_startSoftReset[0];
      end
    end
  end

  always @(*) begin
    when_BusSlaveFactory_l377 = 1'b0;
    case(io_ctrl_cmd_payload_fragment_address)
      12'h008 : begin
        if(ctrl_doWrite) begin
          when_BusSlaveFactory_l377 = 1'b1;
        end
      end
      default : begin
      end
    endcase
  end

  assign when_BusSlaveFactory_l379 = io_ctrl_cmd_payload_fragment_data[0];
  always @(*) begin
    when_BusSlaveFactory_l377_1 = 1'b0;
    case(io_ctrl_cmd_payload_fragment_address)
      12'h008 : begin
        if(ctrl_doWrite) begin
          when_BusSlaveFactory_l377_1 = 1'b1;
        end
      end
      default : begin
      end
    endcase
  end

  assign when_BusSlaveFactory_l379_1 = io_ctrl_cmd_payload_fragment_data[1];
  always @(*) begin
    when_BusSlaveFactory_l377_2 = 1'b0;
    case(io_ctrl_cmd_payload_fragment_address)
      12'h008 : begin
        if(ctrl_doWrite) begin
          when_BusSlaveFactory_l377_2 = 1'b1;
        end
      end
      default : begin
      end
    endcase
  end

  assign when_BusSlaveFactory_l379_2 = io_ctrl_cmd_payload_fragment_data[2];
  always @(*) begin
    when_BusSlaveFactory_l377_3 = 1'b0;
    case(io_ctrl_cmd_payload_fragment_address)
      12'h008 : begin
        if(ctrl_doWrite) begin
          when_BusSlaveFactory_l377_3 = 1'b1;
        end
      end
      default : begin
      end
    endcase
  end

  assign when_BusSlaveFactory_l379_3 = io_ctrl_cmd_payload_fragment_data[3];
  always @(*) begin
    reg_hcInterrupt_unmaskedPending = 1'b0;
    if(when_UsbOhci_l290) begin
      reg_hcInterrupt_unmaskedPending = 1'b1;
    end
    if(when_UsbOhci_l290_1) begin
      reg_hcInterrupt_unmaskedPending = 1'b1;
    end
    if(when_UsbOhci_l290_2) begin
      reg_hcInterrupt_unmaskedPending = 1'b1;
    end
    if(when_UsbOhci_l290_3) begin
      reg_hcInterrupt_unmaskedPending = 1'b1;
    end
    if(when_UsbOhci_l290_4) begin
      reg_hcInterrupt_unmaskedPending = 1'b1;
    end
    if(when_UsbOhci_l290_5) begin
      reg_hcInterrupt_unmaskedPending = 1'b1;
    end
    if(when_UsbOhci_l290_6) begin
      reg_hcInterrupt_unmaskedPending = 1'b1;
    end
  end

  always @(*) begin
    when_BusSlaveFactory_l377_4 = 1'b0;
    case(io_ctrl_cmd_payload_fragment_address)
      12'h010 : begin
        if(ctrl_doWrite) begin
          when_BusSlaveFactory_l377_4 = 1'b1;
        end
      end
      default : begin
      end
    endcase
  end

  assign when_BusSlaveFactory_l379_4 = io_ctrl_cmd_payload_fragment_data[31];
  always @(*) begin
    when_BusSlaveFactory_l341 = 1'b0;
    case(io_ctrl_cmd_payload_fragment_address)
      12'h014 : begin
        if(ctrl_doWrite) begin
          when_BusSlaveFactory_l341 = 1'b1;
        end
      end
      default : begin
      end
    endcase
  end

  assign when_BusSlaveFactory_l347 = io_ctrl_cmd_payload_fragment_data[31];
  always @(*) begin
    when_BusSlaveFactory_l341_1 = 1'b0;
    case(io_ctrl_cmd_payload_fragment_address)
      12'h00c : begin
        if(ctrl_doWrite) begin
          when_BusSlaveFactory_l341_1 = 1'b1;
        end
      end
      default : begin
      end
    endcase
  end

  assign when_BusSlaveFactory_l347_1 = io_ctrl_cmd_payload_fragment_data[0];
  always @(*) begin
    when_BusSlaveFactory_l377_5 = 1'b0;
    case(io_ctrl_cmd_payload_fragment_address)
      12'h010 : begin
        if(ctrl_doWrite) begin
          when_BusSlaveFactory_l377_5 = 1'b1;
        end
      end
      default : begin
      end
    endcase
  end

  assign when_BusSlaveFactory_l379_5 = io_ctrl_cmd_payload_fragment_data[0];
  always @(*) begin
    when_BusSlaveFactory_l341_2 = 1'b0;
    case(io_ctrl_cmd_payload_fragment_address)
      12'h014 : begin
        if(ctrl_doWrite) begin
          when_BusSlaveFactory_l341_2 = 1'b1;
        end
      end
      default : begin
      end
    endcase
  end

  assign when_BusSlaveFactory_l347_2 = io_ctrl_cmd_payload_fragment_data[0];
  assign when_UsbOhci_l290 = (reg_hcInterrupt_SO_status && reg_hcInterrupt_SO_enable);
  always @(*) begin
    when_BusSlaveFactory_l341_3 = 1'b0;
    case(io_ctrl_cmd_payload_fragment_address)
      12'h00c : begin
        if(ctrl_doWrite) begin
          when_BusSlaveFactory_l341_3 = 1'b1;
        end
      end
      default : begin
      end
    endcase
  end

  assign when_BusSlaveFactory_l347_3 = io_ctrl_cmd_payload_fragment_data[1];
  always @(*) begin
    when_BusSlaveFactory_l377_6 = 1'b0;
    case(io_ctrl_cmd_payload_fragment_address)
      12'h010 : begin
        if(ctrl_doWrite) begin
          when_BusSlaveFactory_l377_6 = 1'b1;
        end
      end
      default : begin
      end
    endcase
  end

  assign when_BusSlaveFactory_l379_6 = io_ctrl_cmd_payload_fragment_data[1];
  always @(*) begin
    when_BusSlaveFactory_l341_4 = 1'b0;
    case(io_ctrl_cmd_payload_fragment_address)
      12'h014 : begin
        if(ctrl_doWrite) begin
          when_BusSlaveFactory_l341_4 = 1'b1;
        end
      end
      default : begin
      end
    endcase
  end

  assign when_BusSlaveFactory_l347_4 = io_ctrl_cmd_payload_fragment_data[1];
  assign when_UsbOhci_l290_1 = (reg_hcInterrupt_WDH_status && reg_hcInterrupt_WDH_enable);
  always @(*) begin
    when_BusSlaveFactory_l341_5 = 1'b0;
    case(io_ctrl_cmd_payload_fragment_address)
      12'h00c : begin
        if(ctrl_doWrite) begin
          when_BusSlaveFactory_l341_5 = 1'b1;
        end
      end
      default : begin
      end
    endcase
  end

  assign when_BusSlaveFactory_l347_5 = io_ctrl_cmd_payload_fragment_data[2];
  always @(*) begin
    when_BusSlaveFactory_l377_7 = 1'b0;
    case(io_ctrl_cmd_payload_fragment_address)
      12'h010 : begin
        if(ctrl_doWrite) begin
          when_BusSlaveFactory_l377_7 = 1'b1;
        end
      end
      default : begin
      end
    endcase
  end

  assign when_BusSlaveFactory_l379_7 = io_ctrl_cmd_payload_fragment_data[2];
  always @(*) begin
    when_BusSlaveFactory_l341_6 = 1'b0;
    case(io_ctrl_cmd_payload_fragment_address)
      12'h014 : begin
        if(ctrl_doWrite) begin
          when_BusSlaveFactory_l341_6 = 1'b1;
        end
      end
      default : begin
      end
    endcase
  end

  assign when_BusSlaveFactory_l347_6 = io_ctrl_cmd_payload_fragment_data[2];
  assign when_UsbOhci_l290_2 = (reg_hcInterrupt_SF_status && reg_hcInterrupt_SF_enable);
  always @(*) begin
    when_BusSlaveFactory_l341_7 = 1'b0;
    case(io_ctrl_cmd_payload_fragment_address)
      12'h00c : begin
        if(ctrl_doWrite) begin
          when_BusSlaveFactory_l341_7 = 1'b1;
        end
      end
      default : begin
      end
    endcase
  end

  assign when_BusSlaveFactory_l347_7 = io_ctrl_cmd_payload_fragment_data[3];
  always @(*) begin
    when_BusSlaveFactory_l377_8 = 1'b0;
    case(io_ctrl_cmd_payload_fragment_address)
      12'h010 : begin
        if(ctrl_doWrite) begin
          when_BusSlaveFactory_l377_8 = 1'b1;
        end
      end
      default : begin
      end
    endcase
  end

  assign when_BusSlaveFactory_l379_8 = io_ctrl_cmd_payload_fragment_data[3];
  always @(*) begin
    when_BusSlaveFactory_l341_8 = 1'b0;
    case(io_ctrl_cmd_payload_fragment_address)
      12'h014 : begin
        if(ctrl_doWrite) begin
          when_BusSlaveFactory_l341_8 = 1'b1;
        end
      end
      default : begin
      end
    endcase
  end

  assign when_BusSlaveFactory_l347_8 = io_ctrl_cmd_payload_fragment_data[3];
  assign when_UsbOhci_l290_3 = (reg_hcInterrupt_RD_status && reg_hcInterrupt_RD_enable);
  always @(*) begin
    when_BusSlaveFactory_l341_9 = 1'b0;
    case(io_ctrl_cmd_payload_fragment_address)
      12'h00c : begin
        if(ctrl_doWrite) begin
          when_BusSlaveFactory_l341_9 = 1'b1;
        end
      end
      default : begin
      end
    endcase
  end

  assign when_BusSlaveFactory_l347_9 = io_ctrl_cmd_payload_fragment_data[4];
  always @(*) begin
    when_BusSlaveFactory_l377_9 = 1'b0;
    case(io_ctrl_cmd_payload_fragment_address)
      12'h010 : begin
        if(ctrl_doWrite) begin
          when_BusSlaveFactory_l377_9 = 1'b1;
        end
      end
      default : begin
      end
    endcase
  end

  assign when_BusSlaveFactory_l379_9 = io_ctrl_cmd_payload_fragment_data[4];
  always @(*) begin
    when_BusSlaveFactory_l341_10 = 1'b0;
    case(io_ctrl_cmd_payload_fragment_address)
      12'h014 : begin
        if(ctrl_doWrite) begin
          when_BusSlaveFactory_l341_10 = 1'b1;
        end
      end
      default : begin
      end
    endcase
  end

  assign when_BusSlaveFactory_l347_10 = io_ctrl_cmd_payload_fragment_data[4];
  assign when_UsbOhci_l290_4 = (reg_hcInterrupt_UE_status && reg_hcInterrupt_UE_enable);
  always @(*) begin
    when_BusSlaveFactory_l341_11 = 1'b0;
    case(io_ctrl_cmd_payload_fragment_address)
      12'h00c : begin
        if(ctrl_doWrite) begin
          when_BusSlaveFactory_l341_11 = 1'b1;
        end
      end
      default : begin
      end
    endcase
  end

  assign when_BusSlaveFactory_l347_11 = io_ctrl_cmd_payload_fragment_data[5];
  always @(*) begin
    when_BusSlaveFactory_l377_10 = 1'b0;
    case(io_ctrl_cmd_payload_fragment_address)
      12'h010 : begin
        if(ctrl_doWrite) begin
          when_BusSlaveFactory_l377_10 = 1'b1;
        end
      end
      default : begin
      end
    endcase
  end

  assign when_BusSlaveFactory_l379_10 = io_ctrl_cmd_payload_fragment_data[5];
  always @(*) begin
    when_BusSlaveFactory_l341_12 = 1'b0;
    case(io_ctrl_cmd_payload_fragment_address)
      12'h014 : begin
        if(ctrl_doWrite) begin
          when_BusSlaveFactory_l341_12 = 1'b1;
        end
      end
      default : begin
      end
    endcase
  end

  assign when_BusSlaveFactory_l347_12 = io_ctrl_cmd_payload_fragment_data[5];
  assign when_UsbOhci_l290_5 = (reg_hcInterrupt_FNO_status && reg_hcInterrupt_FNO_enable);
  always @(*) begin
    when_BusSlaveFactory_l341_13 = 1'b0;
    case(io_ctrl_cmd_payload_fragment_address)
      12'h00c : begin
        if(ctrl_doWrite) begin
          when_BusSlaveFactory_l341_13 = 1'b1;
        end
      end
      default : begin
      end
    endcase
  end

  assign when_BusSlaveFactory_l347_13 = io_ctrl_cmd_payload_fragment_data[6];
  always @(*) begin
    when_BusSlaveFactory_l377_11 = 1'b0;
    case(io_ctrl_cmd_payload_fragment_address)
      12'h010 : begin
        if(ctrl_doWrite) begin
          when_BusSlaveFactory_l377_11 = 1'b1;
        end
      end
      default : begin
      end
    endcase
  end

  assign when_BusSlaveFactory_l379_11 = io_ctrl_cmd_payload_fragment_data[6];
  always @(*) begin
    when_BusSlaveFactory_l341_14 = 1'b0;
    case(io_ctrl_cmd_payload_fragment_address)
      12'h014 : begin
        if(ctrl_doWrite) begin
          when_BusSlaveFactory_l341_14 = 1'b1;
        end
      end
      default : begin
      end
    endcase
  end

  assign when_BusSlaveFactory_l347_14 = io_ctrl_cmd_payload_fragment_data[6];
  assign when_UsbOhci_l290_6 = (reg_hcInterrupt_RHSC_status && reg_hcInterrupt_RHSC_enable);
  always @(*) begin
    when_BusSlaveFactory_l341_15 = 1'b0;
    case(io_ctrl_cmd_payload_fragment_address)
      12'h00c : begin
        if(ctrl_doWrite) begin
          when_BusSlaveFactory_l341_15 = 1'b1;
        end
      end
      default : begin
      end
    endcase
  end

  assign when_BusSlaveFactory_l347_15 = io_ctrl_cmd_payload_fragment_data[30];
  always @(*) begin
    when_BusSlaveFactory_l377_12 = 1'b0;
    case(io_ctrl_cmd_payload_fragment_address)
      12'h010 : begin
        if(ctrl_doWrite) begin
          when_BusSlaveFactory_l377_12 = 1'b1;
        end
      end
      default : begin
      end
    endcase
  end

  assign when_BusSlaveFactory_l379_12 = io_ctrl_cmd_payload_fragment_data[30];
  always @(*) begin
    when_BusSlaveFactory_l341_16 = 1'b0;
    case(io_ctrl_cmd_payload_fragment_address)
      12'h014 : begin
        if(ctrl_doWrite) begin
          when_BusSlaveFactory_l341_16 = 1'b1;
        end
      end
      default : begin
      end
    endcase
  end

  assign when_BusSlaveFactory_l347_16 = io_ctrl_cmd_payload_fragment_data[30];
  assign reg_hcInterrupt_doIrq = (reg_hcInterrupt_unmaskedPending && reg_hcInterrupt_MIE);
  assign io_interrupt = (reg_hcInterrupt_doIrq && (! reg_hcControl_IR));
  assign io_interruptBios = ((reg_hcInterrupt_doIrq && reg_hcControl_IR) || (reg_hcInterrupt_OC_status && reg_hcInterrupt_OC_enable));
  assign reg_hcHCCA_HCCA_address = {reg_hcHCCA_HCCA_reg,8'h0};
  assign reg_hcPeriodCurrentED_PCED_address = {reg_hcPeriodCurrentED_PCED_reg,4'b0000};
  assign reg_hcPeriodCurrentED_isZero = (reg_hcPeriodCurrentED_PCED_reg == 28'h0);
  assign reg_hcControlHeadED_CHED_address = {reg_hcControlHeadED_CHED_reg,4'b0000};
  assign reg_hcControlCurrentED_CCED_address = {reg_hcControlCurrentED_CCED_reg,4'b0000};
  assign reg_hcControlCurrentED_isZero = (reg_hcControlCurrentED_CCED_reg == 28'h0);
  assign reg_hcBulkHeadED_BHED_address = {reg_hcBulkHeadED_BHED_reg,4'b0000};
  assign reg_hcBulkCurrentED_BCED_address = {reg_hcBulkCurrentED_BCED_reg,4'b0000};
  assign reg_hcBulkCurrentED_isZero = (reg_hcBulkCurrentED_BCED_reg == 28'h0);
  assign reg_hcDoneHead_DH_address = {reg_hcDoneHead_DH_reg,4'b0000};
  assign reg_hcFmNumber_FNp1 = (reg_hcFmNumber_FN + 16'h0001);
  assign reg_hcLSThreshold_hit = (reg_hcFmRemaining_FR < _zz_reg_hcLSThreshold_hit);
  assign reg_hcRhDescriptorA_NDP = 8'h02;
  always @(*) begin
    when_BusSlaveFactory_l341_17 = 1'b0;
    case(io_ctrl_cmd_payload_fragment_address)
      12'h050 : begin
        if(ctrl_doWrite) begin
          when_BusSlaveFactory_l341_17 = 1'b1;
        end
      end
      default : begin
      end
    endcase
  end

  assign when_BusSlaveFactory_l347_17 = io_ctrl_cmd_payload_fragment_data[17];
  assign when_UsbOhci_l397 = (io_phy_overcurrent ^ io_phy_overcurrent_regNext);
  always @(*) begin
    reg_hcRhStatus_clearGlobalPower = 1'b0;
    if(when_BusSlaveFactory_l377_13) begin
      if(when_BusSlaveFactory_l379_13) begin
        reg_hcRhStatus_clearGlobalPower = _zz_reg_hcRhStatus_clearGlobalPower[0];
      end
    end
  end

  always @(*) begin
    when_BusSlaveFactory_l377_13 = 1'b0;
    case(io_ctrl_cmd_payload_fragment_address)
      12'h050 : begin
        if(ctrl_doWrite) begin
          when_BusSlaveFactory_l377_13 = 1'b1;
        end
      end
      default : begin
      end
    endcase
  end

  assign when_BusSlaveFactory_l379_13 = io_ctrl_cmd_payload_fragment_data[0];
  always @(*) begin
    reg_hcRhStatus_setRemoteWakeupEnable = 1'b0;
    if(when_BusSlaveFactory_l377_14) begin
      if(when_BusSlaveFactory_l379_14) begin
        reg_hcRhStatus_setRemoteWakeupEnable = _zz_reg_hcRhStatus_setRemoteWakeupEnable[0];
      end
    end
  end

  always @(*) begin
    when_BusSlaveFactory_l377_14 = 1'b0;
    case(io_ctrl_cmd_payload_fragment_address)
      12'h050 : begin
        if(ctrl_doWrite) begin
          when_BusSlaveFactory_l377_14 = 1'b1;
        end
      end
      default : begin
      end
    endcase
  end

  assign when_BusSlaveFactory_l379_14 = io_ctrl_cmd_payload_fragment_data[15];
  always @(*) begin
    reg_hcRhStatus_setGlobalPower = 1'b0;
    if(when_BusSlaveFactory_l377_15) begin
      if(when_BusSlaveFactory_l379_15) begin
        reg_hcRhStatus_setGlobalPower = _zz_reg_hcRhStatus_setGlobalPower[0];
      end
    end
  end

  always @(*) begin
    when_BusSlaveFactory_l377_15 = 1'b0;
    case(io_ctrl_cmd_payload_fragment_address)
      12'h050 : begin
        if(ctrl_doWrite) begin
          when_BusSlaveFactory_l377_15 = 1'b1;
        end
      end
      default : begin
      end
    endcase
  end

  assign when_BusSlaveFactory_l379_15 = io_ctrl_cmd_payload_fragment_data[16];
  always @(*) begin
    reg_hcRhStatus_clearRemoteWakeupEnable = 1'b0;
    if(when_BusSlaveFactory_l377_16) begin
      if(when_BusSlaveFactory_l379_16) begin
        reg_hcRhStatus_clearRemoteWakeupEnable = _zz_reg_hcRhStatus_clearRemoteWakeupEnable[0];
      end
    end
  end

  always @(*) begin
    when_BusSlaveFactory_l377_16 = 1'b0;
    case(io_ctrl_cmd_payload_fragment_address)
      12'h050 : begin
        if(ctrl_doWrite) begin
          when_BusSlaveFactory_l377_16 = 1'b1;
        end
      end
      default : begin
      end
    endcase
  end

  assign when_BusSlaveFactory_l379_16 = io_ctrl_cmd_payload_fragment_data[31];
  always @(*) begin
    reg_hcRhPortStatus_0_clearPortEnable = 1'b0;
    if(when_BusSlaveFactory_l377_17) begin
      if(when_BusSlaveFactory_l379_17) begin
        reg_hcRhPortStatus_0_clearPortEnable = _zz_reg_hcRhPortStatus_0_clearPortEnable[0];
      end
    end
  end

  always @(*) begin
    when_BusSlaveFactory_l377_17 = 1'b0;
    case(io_ctrl_cmd_payload_fragment_address)
      12'h054 : begin
        if(ctrl_doWrite) begin
          when_BusSlaveFactory_l377_17 = 1'b1;
        end
      end
      default : begin
      end
    endcase
  end

  assign when_BusSlaveFactory_l379_17 = io_ctrl_cmd_payload_fragment_data[0];
  always @(*) begin
    reg_hcRhPortStatus_0_setPortEnable = 1'b0;
    if(when_BusSlaveFactory_l377_18) begin
      if(when_BusSlaveFactory_l379_18) begin
        reg_hcRhPortStatus_0_setPortEnable = _zz_reg_hcRhPortStatus_0_setPortEnable[0];
      end
    end
  end

  always @(*) begin
    when_BusSlaveFactory_l377_18 = 1'b0;
    case(io_ctrl_cmd_payload_fragment_address)
      12'h054 : begin
        if(ctrl_doWrite) begin
          when_BusSlaveFactory_l377_18 = 1'b1;
        end
      end
      default : begin
      end
    endcase
  end

  assign when_BusSlaveFactory_l379_18 = io_ctrl_cmd_payload_fragment_data[1];
  always @(*) begin
    reg_hcRhPortStatus_0_setPortSuspend = 1'b0;
    if(when_BusSlaveFactory_l377_19) begin
      if(when_BusSlaveFactory_l379_19) begin
        reg_hcRhPortStatus_0_setPortSuspend = _zz_reg_hcRhPortStatus_0_setPortSuspend[0];
      end
    end
  end

  always @(*) begin
    when_BusSlaveFactory_l377_19 = 1'b0;
    case(io_ctrl_cmd_payload_fragment_address)
      12'h054 : begin
        if(ctrl_doWrite) begin
          when_BusSlaveFactory_l377_19 = 1'b1;
        end
      end
      default : begin
      end
    endcase
  end

  assign when_BusSlaveFactory_l379_19 = io_ctrl_cmd_payload_fragment_data[2];
  always @(*) begin
    reg_hcRhPortStatus_0_clearSuspendStatus = 1'b0;
    if(when_BusSlaveFactory_l377_20) begin
      if(when_BusSlaveFactory_l379_20) begin
        reg_hcRhPortStatus_0_clearSuspendStatus = _zz_reg_hcRhPortStatus_0_clearSuspendStatus[0];
      end
    end
  end

  always @(*) begin
    when_BusSlaveFactory_l377_20 = 1'b0;
    case(io_ctrl_cmd_payload_fragment_address)
      12'h054 : begin
        if(ctrl_doWrite) begin
          when_BusSlaveFactory_l377_20 = 1'b1;
        end
      end
      default : begin
      end
    endcase
  end

  assign when_BusSlaveFactory_l379_20 = io_ctrl_cmd_payload_fragment_data[3];
  always @(*) begin
    reg_hcRhPortStatus_0_setPortReset = 1'b0;
    if(when_BusSlaveFactory_l377_21) begin
      if(when_BusSlaveFactory_l379_21) begin
        reg_hcRhPortStatus_0_setPortReset = _zz_reg_hcRhPortStatus_0_setPortReset[0];
      end
    end
  end

  always @(*) begin
    when_BusSlaveFactory_l377_21 = 1'b0;
    case(io_ctrl_cmd_payload_fragment_address)
      12'h054 : begin
        if(ctrl_doWrite) begin
          when_BusSlaveFactory_l377_21 = 1'b1;
        end
      end
      default : begin
      end
    endcase
  end

  assign when_BusSlaveFactory_l379_21 = io_ctrl_cmd_payload_fragment_data[4];
  always @(*) begin
    reg_hcRhPortStatus_0_setPortPower = 1'b0;
    if(when_BusSlaveFactory_l377_22) begin
      if(when_BusSlaveFactory_l379_22) begin
        reg_hcRhPortStatus_0_setPortPower = _zz_reg_hcRhPortStatus_0_setPortPower[0];
      end
    end
  end

  always @(*) begin
    when_BusSlaveFactory_l377_22 = 1'b0;
    case(io_ctrl_cmd_payload_fragment_address)
      12'h054 : begin
        if(ctrl_doWrite) begin
          when_BusSlaveFactory_l377_22 = 1'b1;
        end
      end
      default : begin
      end
    endcase
  end

  assign when_BusSlaveFactory_l379_22 = io_ctrl_cmd_payload_fragment_data[8];
  always @(*) begin
    reg_hcRhPortStatus_0_clearPortPower = 1'b0;
    if(when_BusSlaveFactory_l377_23) begin
      if(when_BusSlaveFactory_l379_23) begin
        reg_hcRhPortStatus_0_clearPortPower = _zz_reg_hcRhPortStatus_0_clearPortPower[0];
      end
    end
  end

  always @(*) begin
    when_BusSlaveFactory_l377_23 = 1'b0;
    case(io_ctrl_cmd_payload_fragment_address)
      12'h054 : begin
        if(ctrl_doWrite) begin
          when_BusSlaveFactory_l377_23 = 1'b1;
        end
      end
      default : begin
      end
    endcase
  end

  assign when_BusSlaveFactory_l379_23 = io_ctrl_cmd_payload_fragment_data[9];
  assign reg_hcRhPortStatus_0_CCS = ((reg_hcRhPortStatus_0_connected || reg_hcRhDescriptorB_DR[0]) && reg_hcRhPortStatus_0_PPS);
  always @(*) begin
    reg_hcRhPortStatus_0_CSC_clear = 1'b0;
    if(when_BusSlaveFactory_l377_24) begin
      if(when_BusSlaveFactory_l379_24) begin
        reg_hcRhPortStatus_0_CSC_clear = _zz_reg_hcRhPortStatus_0_CSC_clear[0];
      end
    end
  end

  always @(*) begin
    when_BusSlaveFactory_l377_24 = 1'b0;
    case(io_ctrl_cmd_payload_fragment_address)
      12'h054 : begin
        if(ctrl_doWrite) begin
          when_BusSlaveFactory_l377_24 = 1'b1;
        end
      end
      default : begin
      end
    endcase
  end

  assign when_BusSlaveFactory_l379_24 = io_ctrl_cmd_payload_fragment_data[16];
  always @(*) begin
    reg_hcRhPortStatus_0_PESC_clear = 1'b0;
    if(when_BusSlaveFactory_l377_25) begin
      if(when_BusSlaveFactory_l379_25) begin
        reg_hcRhPortStatus_0_PESC_clear = _zz_reg_hcRhPortStatus_0_PESC_clear[0];
      end
    end
  end

  always @(*) begin
    when_BusSlaveFactory_l377_25 = 1'b0;
    case(io_ctrl_cmd_payload_fragment_address)
      12'h054 : begin
        if(ctrl_doWrite) begin
          when_BusSlaveFactory_l377_25 = 1'b1;
        end
      end
      default : begin
      end
    endcase
  end

  assign when_BusSlaveFactory_l379_25 = io_ctrl_cmd_payload_fragment_data[17];
  always @(*) begin
    reg_hcRhPortStatus_0_PSSC_clear = 1'b0;
    if(when_BusSlaveFactory_l377_26) begin
      if(when_BusSlaveFactory_l379_26) begin
        reg_hcRhPortStatus_0_PSSC_clear = _zz_reg_hcRhPortStatus_0_PSSC_clear[0];
      end
    end
    if(reg_hcRhPortStatus_0_PRSC_set) begin
      reg_hcRhPortStatus_0_PSSC_clear = 1'b1;
    end
  end

  always @(*) begin
    when_BusSlaveFactory_l377_26 = 1'b0;
    case(io_ctrl_cmd_payload_fragment_address)
      12'h054 : begin
        if(ctrl_doWrite) begin
          when_BusSlaveFactory_l377_26 = 1'b1;
        end
      end
      default : begin
      end
    endcase
  end

  assign when_BusSlaveFactory_l379_26 = io_ctrl_cmd_payload_fragment_data[18];
  always @(*) begin
    reg_hcRhPortStatus_0_OCIC_clear = 1'b0;
    if(when_BusSlaveFactory_l377_27) begin
      if(when_BusSlaveFactory_l379_27) begin
        reg_hcRhPortStatus_0_OCIC_clear = _zz_reg_hcRhPortStatus_0_OCIC_clear[0];
      end
    end
  end

  always @(*) begin
    when_BusSlaveFactory_l377_27 = 1'b0;
    case(io_ctrl_cmd_payload_fragment_address)
      12'h054 : begin
        if(ctrl_doWrite) begin
          when_BusSlaveFactory_l377_27 = 1'b1;
        end
      end
      default : begin
      end
    endcase
  end

  assign when_BusSlaveFactory_l379_27 = io_ctrl_cmd_payload_fragment_data[19];
  always @(*) begin
    reg_hcRhPortStatus_0_PRSC_clear = 1'b0;
    if(when_BusSlaveFactory_l377_28) begin
      if(when_BusSlaveFactory_l379_28) begin
        reg_hcRhPortStatus_0_PRSC_clear = _zz_reg_hcRhPortStatus_0_PRSC_clear[0];
      end
    end
  end

  always @(*) begin
    when_BusSlaveFactory_l377_28 = 1'b0;
    case(io_ctrl_cmd_payload_fragment_address)
      12'h054 : begin
        if(ctrl_doWrite) begin
          when_BusSlaveFactory_l377_28 = 1'b1;
        end
      end
      default : begin
      end
    endcase
  end

  assign when_BusSlaveFactory_l379_28 = io_ctrl_cmd_payload_fragment_data[20];
  assign when_UsbOhci_l448 = ((reg_hcRhPortStatus_0_clearPortEnable || reg_hcRhPortStatus_0_PESC_set) || (! reg_hcRhPortStatus_0_PPS));
  assign when_UsbOhci_l448_1 = (reg_hcRhPortStatus_0_PRSC_set || reg_hcRhPortStatus_0_PSSC_set);
  assign when_UsbOhci_l448_2 = (reg_hcRhPortStatus_0_setPortEnable && reg_hcRhPortStatus_0_CCS);
  assign when_UsbOhci_l449 = (((reg_hcRhPortStatus_0_PSSC_set || reg_hcRhPortStatus_0_PRSC_set) || (! reg_hcRhPortStatus_0_PPS)) || (reg_hcControl_HCFS == MainState_RESUME));
  assign when_UsbOhci_l449_1 = (reg_hcRhPortStatus_0_setPortSuspend && reg_hcRhPortStatus_0_CCS);
  assign when_UsbOhci_l450 = (reg_hcRhPortStatus_0_setPortSuspend && reg_hcRhPortStatus_0_CCS);
  assign when_UsbOhci_l451 = (reg_hcRhPortStatus_0_clearSuspendStatus && reg_hcRhPortStatus_0_PSS);
  assign when_UsbOhci_l452 = (reg_hcRhPortStatus_0_setPortReset && reg_hcRhPortStatus_0_CCS);
  assign when_UsbOhci_l458 = reg_hcRhDescriptorB_PPCM[0];
  assign reg_hcRhPortStatus_0_CSC_set = ((((reg_hcRhPortStatus_0_CCS ^ reg_hcRhPortStatus_0_CCS_regNext) || (reg_hcRhPortStatus_0_setPortEnable && (! reg_hcRhPortStatus_0_CCS))) || (reg_hcRhPortStatus_0_setPortSuspend && (! reg_hcRhPortStatus_0_CCS))) || (reg_hcRhPortStatus_0_setPortReset && (! reg_hcRhPortStatus_0_CCS)));
  assign reg_hcRhPortStatus_0_PESC_set = io_phy_ports_0_overcurrent;
  assign io_phy_ports_0_suspend_fire = (io_phy_ports_0_suspend_valid && io_phy_ports_0_suspend_ready);
  assign reg_hcRhPortStatus_0_PSSC_set = (io_phy_ports_0_suspend_fire || io_phy_ports_0_remoteResume);
  assign reg_hcRhPortStatus_0_OCIC_set = io_phy_ports_0_overcurrent;
  assign io_phy_ports_0_reset_fire = (io_phy_ports_0_reset_valid && io_phy_ports_0_reset_ready);
  assign reg_hcRhPortStatus_0_PRSC_set = io_phy_ports_0_reset_fire;
  assign io_phy_ports_0_disable_valid = reg_hcRhPortStatus_0_clearPortEnable;
  assign io_phy_ports_0_removable = reg_hcRhDescriptorB_DR[0];
  assign io_phy_ports_0_power = reg_hcRhPortStatus_0_PPS;
  assign io_phy_ports_0_resume_valid = reg_hcRhPortStatus_0_resume;
  assign io_phy_ports_0_resume_fire = (io_phy_ports_0_resume_valid && io_phy_ports_0_resume_ready);
  assign io_phy_ports_0_reset_valid = reg_hcRhPortStatus_0_reset;
  assign io_phy_ports_0_suspend_valid = reg_hcRhPortStatus_0_suspend;
  always @(*) begin
    reg_hcRhPortStatus_1_clearPortEnable = 1'b0;
    if(when_BusSlaveFactory_l377_29) begin
      if(when_BusSlaveFactory_l379_29) begin
        reg_hcRhPortStatus_1_clearPortEnable = _zz_reg_hcRhPortStatus_1_clearPortEnable[0];
      end
    end
  end

  always @(*) begin
    when_BusSlaveFactory_l377_29 = 1'b0;
    case(io_ctrl_cmd_payload_fragment_address)
      12'h058 : begin
        if(ctrl_doWrite) begin
          when_BusSlaveFactory_l377_29 = 1'b1;
        end
      end
      default : begin
      end
    endcase
  end

  assign when_BusSlaveFactory_l379_29 = io_ctrl_cmd_payload_fragment_data[0];
  always @(*) begin
    reg_hcRhPortStatus_1_setPortEnable = 1'b0;
    if(when_BusSlaveFactory_l377_30) begin
      if(when_BusSlaveFactory_l379_30) begin
        reg_hcRhPortStatus_1_setPortEnable = _zz_reg_hcRhPortStatus_1_setPortEnable[0];
      end
    end
  end

  always @(*) begin
    when_BusSlaveFactory_l377_30 = 1'b0;
    case(io_ctrl_cmd_payload_fragment_address)
      12'h058 : begin
        if(ctrl_doWrite) begin
          when_BusSlaveFactory_l377_30 = 1'b1;
        end
      end
      default : begin
      end
    endcase
  end

  assign when_BusSlaveFactory_l379_30 = io_ctrl_cmd_payload_fragment_data[1];
  always @(*) begin
    reg_hcRhPortStatus_1_setPortSuspend = 1'b0;
    if(when_BusSlaveFactory_l377_31) begin
      if(when_BusSlaveFactory_l379_31) begin
        reg_hcRhPortStatus_1_setPortSuspend = _zz_reg_hcRhPortStatus_1_setPortSuspend[0];
      end
    end
  end

  always @(*) begin
    when_BusSlaveFactory_l377_31 = 1'b0;
    case(io_ctrl_cmd_payload_fragment_address)
      12'h058 : begin
        if(ctrl_doWrite) begin
          when_BusSlaveFactory_l377_31 = 1'b1;
        end
      end
      default : begin
      end
    endcase
  end

  assign when_BusSlaveFactory_l379_31 = io_ctrl_cmd_payload_fragment_data[2];
  always @(*) begin
    reg_hcRhPortStatus_1_clearSuspendStatus = 1'b0;
    if(when_BusSlaveFactory_l377_32) begin
      if(when_BusSlaveFactory_l379_32) begin
        reg_hcRhPortStatus_1_clearSuspendStatus = _zz_reg_hcRhPortStatus_1_clearSuspendStatus[0];
      end
    end
  end

  always @(*) begin
    when_BusSlaveFactory_l377_32 = 1'b0;
    case(io_ctrl_cmd_payload_fragment_address)
      12'h058 : begin
        if(ctrl_doWrite) begin
          when_BusSlaveFactory_l377_32 = 1'b1;
        end
      end
      default : begin
      end
    endcase
  end

  assign when_BusSlaveFactory_l379_32 = io_ctrl_cmd_payload_fragment_data[3];
  always @(*) begin
    reg_hcRhPortStatus_1_setPortReset = 1'b0;
    if(when_BusSlaveFactory_l377_33) begin
      if(when_BusSlaveFactory_l379_33) begin
        reg_hcRhPortStatus_1_setPortReset = _zz_reg_hcRhPortStatus_1_setPortReset[0];
      end
    end
  end

  always @(*) begin
    when_BusSlaveFactory_l377_33 = 1'b0;
    case(io_ctrl_cmd_payload_fragment_address)
      12'h058 : begin
        if(ctrl_doWrite) begin
          when_BusSlaveFactory_l377_33 = 1'b1;
        end
      end
      default : begin
      end
    endcase
  end

  assign when_BusSlaveFactory_l379_33 = io_ctrl_cmd_payload_fragment_data[4];
  always @(*) begin
    reg_hcRhPortStatus_1_setPortPower = 1'b0;
    if(when_BusSlaveFactory_l377_34) begin
      if(when_BusSlaveFactory_l379_34) begin
        reg_hcRhPortStatus_1_setPortPower = _zz_reg_hcRhPortStatus_1_setPortPower[0];
      end
    end
  end

  always @(*) begin
    when_BusSlaveFactory_l377_34 = 1'b0;
    case(io_ctrl_cmd_payload_fragment_address)
      12'h058 : begin
        if(ctrl_doWrite) begin
          when_BusSlaveFactory_l377_34 = 1'b1;
        end
      end
      default : begin
      end
    endcase
  end

  assign when_BusSlaveFactory_l379_34 = io_ctrl_cmd_payload_fragment_data[8];
  always @(*) begin
    reg_hcRhPortStatus_1_clearPortPower = 1'b0;
    if(when_BusSlaveFactory_l377_35) begin
      if(when_BusSlaveFactory_l379_35) begin
        reg_hcRhPortStatus_1_clearPortPower = _zz_reg_hcRhPortStatus_1_clearPortPower[0];
      end
    end
  end

  always @(*) begin
    when_BusSlaveFactory_l377_35 = 1'b0;
    case(io_ctrl_cmd_payload_fragment_address)
      12'h058 : begin
        if(ctrl_doWrite) begin
          when_BusSlaveFactory_l377_35 = 1'b1;
        end
      end
      default : begin
      end
    endcase
  end

  assign when_BusSlaveFactory_l379_35 = io_ctrl_cmd_payload_fragment_data[9];
  assign reg_hcRhPortStatus_1_CCS = ((reg_hcRhPortStatus_1_connected || reg_hcRhDescriptorB_DR[1]) && reg_hcRhPortStatus_1_PPS);
  always @(*) begin
    reg_hcRhPortStatus_1_CSC_clear = 1'b0;
    if(when_BusSlaveFactory_l377_36) begin
      if(when_BusSlaveFactory_l379_36) begin
        reg_hcRhPortStatus_1_CSC_clear = _zz_reg_hcRhPortStatus_1_CSC_clear[0];
      end
    end
  end

  always @(*) begin
    when_BusSlaveFactory_l377_36 = 1'b0;
    case(io_ctrl_cmd_payload_fragment_address)
      12'h058 : begin
        if(ctrl_doWrite) begin
          when_BusSlaveFactory_l377_36 = 1'b1;
        end
      end
      default : begin
      end
    endcase
  end

  assign when_BusSlaveFactory_l379_36 = io_ctrl_cmd_payload_fragment_data[16];
  always @(*) begin
    reg_hcRhPortStatus_1_PESC_clear = 1'b0;
    if(when_BusSlaveFactory_l377_37) begin
      if(when_BusSlaveFactory_l379_37) begin
        reg_hcRhPortStatus_1_PESC_clear = _zz_reg_hcRhPortStatus_1_PESC_clear[0];
      end
    end
  end

  always @(*) begin
    when_BusSlaveFactory_l377_37 = 1'b0;
    case(io_ctrl_cmd_payload_fragment_address)
      12'h058 : begin
        if(ctrl_doWrite) begin
          when_BusSlaveFactory_l377_37 = 1'b1;
        end
      end
      default : begin
      end
    endcase
  end

  assign when_BusSlaveFactory_l379_37 = io_ctrl_cmd_payload_fragment_data[17];
  always @(*) begin
    reg_hcRhPortStatus_1_PSSC_clear = 1'b0;
    if(when_BusSlaveFactory_l377_38) begin
      if(when_BusSlaveFactory_l379_38) begin
        reg_hcRhPortStatus_1_PSSC_clear = _zz_reg_hcRhPortStatus_1_PSSC_clear[0];
      end
    end
    if(reg_hcRhPortStatus_1_PRSC_set) begin
      reg_hcRhPortStatus_1_PSSC_clear = 1'b1;
    end
  end

  always @(*) begin
    when_BusSlaveFactory_l377_38 = 1'b0;
    case(io_ctrl_cmd_payload_fragment_address)
      12'h058 : begin
        if(ctrl_doWrite) begin
          when_BusSlaveFactory_l377_38 = 1'b1;
        end
      end
      default : begin
      end
    endcase
  end

  assign when_BusSlaveFactory_l379_38 = io_ctrl_cmd_payload_fragment_data[18];
  always @(*) begin
    reg_hcRhPortStatus_1_OCIC_clear = 1'b0;
    if(when_BusSlaveFactory_l377_39) begin
      if(when_BusSlaveFactory_l379_39) begin
        reg_hcRhPortStatus_1_OCIC_clear = _zz_reg_hcRhPortStatus_1_OCIC_clear[0];
      end
    end
  end

  always @(*) begin
    when_BusSlaveFactory_l377_39 = 1'b0;
    case(io_ctrl_cmd_payload_fragment_address)
      12'h058 : begin
        if(ctrl_doWrite) begin
          when_BusSlaveFactory_l377_39 = 1'b1;
        end
      end
      default : begin
      end
    endcase
  end

  assign when_BusSlaveFactory_l379_39 = io_ctrl_cmd_payload_fragment_data[19];
  always @(*) begin
    reg_hcRhPortStatus_1_PRSC_clear = 1'b0;
    if(when_BusSlaveFactory_l377_40) begin
      if(when_BusSlaveFactory_l379_40) begin
        reg_hcRhPortStatus_1_PRSC_clear = _zz_reg_hcRhPortStatus_1_PRSC_clear[0];
      end
    end
  end

  always @(*) begin
    when_BusSlaveFactory_l377_40 = 1'b0;
    case(io_ctrl_cmd_payload_fragment_address)
      12'h058 : begin
        if(ctrl_doWrite) begin
          when_BusSlaveFactory_l377_40 = 1'b1;
        end
      end
      default : begin
      end
    endcase
  end

  assign when_BusSlaveFactory_l379_40 = io_ctrl_cmd_payload_fragment_data[20];
  assign when_UsbOhci_l448_3 = ((reg_hcRhPortStatus_1_clearPortEnable || reg_hcRhPortStatus_1_PESC_set) || (! reg_hcRhPortStatus_1_PPS));
  assign when_UsbOhci_l448_4 = (reg_hcRhPortStatus_1_PRSC_set || reg_hcRhPortStatus_1_PSSC_set);
  assign when_UsbOhci_l448_5 = (reg_hcRhPortStatus_1_setPortEnable && reg_hcRhPortStatus_1_CCS);
  assign when_UsbOhci_l449_2 = (((reg_hcRhPortStatus_1_PSSC_set || reg_hcRhPortStatus_1_PRSC_set) || (! reg_hcRhPortStatus_1_PPS)) || (reg_hcControl_HCFS == MainState_RESUME));
  assign when_UsbOhci_l449_3 = (reg_hcRhPortStatus_1_setPortSuspend && reg_hcRhPortStatus_1_CCS);
  assign when_UsbOhci_l450_1 = (reg_hcRhPortStatus_1_setPortSuspend && reg_hcRhPortStatus_1_CCS);
  assign when_UsbOhci_l451_1 = (reg_hcRhPortStatus_1_clearSuspendStatus && reg_hcRhPortStatus_1_PSS);
  assign when_UsbOhci_l452_1 = (reg_hcRhPortStatus_1_setPortReset && reg_hcRhPortStatus_1_CCS);
  assign when_UsbOhci_l458_1 = reg_hcRhDescriptorB_PPCM[1];
  assign reg_hcRhPortStatus_1_CSC_set = ((((reg_hcRhPortStatus_1_CCS ^ reg_hcRhPortStatus_1_CCS_regNext) || (reg_hcRhPortStatus_1_setPortEnable && (! reg_hcRhPortStatus_1_CCS))) || (reg_hcRhPortStatus_1_setPortSuspend && (! reg_hcRhPortStatus_1_CCS))) || (reg_hcRhPortStatus_1_setPortReset && (! reg_hcRhPortStatus_1_CCS)));
  assign reg_hcRhPortStatus_1_PESC_set = io_phy_ports_1_overcurrent;
  assign io_phy_ports_1_suspend_fire = (io_phy_ports_1_suspend_valid && io_phy_ports_1_suspend_ready);
  assign reg_hcRhPortStatus_1_PSSC_set = (io_phy_ports_1_suspend_fire || io_phy_ports_1_remoteResume);
  assign reg_hcRhPortStatus_1_OCIC_set = io_phy_ports_1_overcurrent;
  assign io_phy_ports_1_reset_fire = (io_phy_ports_1_reset_valid && io_phy_ports_1_reset_ready);
  assign reg_hcRhPortStatus_1_PRSC_set = io_phy_ports_1_reset_fire;
  assign io_phy_ports_1_disable_valid = reg_hcRhPortStatus_1_clearPortEnable;
  assign io_phy_ports_1_removable = reg_hcRhDescriptorB_DR[1];
  assign io_phy_ports_1_power = reg_hcRhPortStatus_1_PPS;
  assign io_phy_ports_1_resume_valid = reg_hcRhPortStatus_1_resume;
  assign io_phy_ports_1_resume_fire = (io_phy_ports_1_resume_valid && io_phy_ports_1_resume_ready);
  assign io_phy_ports_1_reset_valid = reg_hcRhPortStatus_1_reset;
  assign io_phy_ports_1_suspend_valid = reg_hcRhPortStatus_1_suspend;
  always @(*) begin
    frame_run = 1'b0;
    case(hc_stateReg)
      hc_enumDef_RESET : begin
      end
      hc_enumDef_RESUME : begin
      end
      hc_enumDef_OPERATIONAL : begin
        frame_run = 1'b1;
      end
      hc_enumDef_SUSPEND : begin
      end
      hc_enumDef_ANY_TO_RESET : begin
      end
      hc_enumDef_ANY_TO_SUSPEND : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    frame_reload = 1'b0;
    if(when_UsbOhci_l514) begin
      if(frame_overflow) begin
        frame_reload = 1'b1;
      end
    end
    if(when_StateMachine_l253_7) begin
      frame_reload = 1'b1;
    end
  end

  assign frame_overflow = (reg_hcFmRemaining_FR == 14'h0);
  always @(*) begin
    frame_tick = 1'b0;
    if(when_UsbOhci_l514) begin
      if(frame_overflow) begin
        frame_tick = 1'b1;
      end
    end
  end

  assign frame_section1 = (reg_hcPeriodicStart_PS < reg_hcFmRemaining_FR);
  assign frame_limitHit = (frame_limitCounter == 15'h0);
  assign frame_decrementTimerOverflow = (frame_decrementTimer == 3'b110);
  assign when_UsbOhci_l514 = (frame_run && io_phy_tick);
  assign when_UsbOhci_l516 = ((! frame_limitHit) && (! frame_decrementTimerOverflow));
  assign when_UsbOhci_l528 = (reg_hcFmNumber_FNp1[15] ^ reg_hcFmNumber_FN[15]);
  always @(*) begin
    token_wantExit = 1'b0;
    case(token_stateReg)
      token_enumDef_INIT : begin
      end
      token_enumDef_PID : begin
      end
      token_enumDef_B1 : begin
      end
      token_enumDef_B2 : begin
      end
      token_enumDef_EOP : begin
        if(io_phy_txEop) begin
          token_wantExit = 1'b1;
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    token_wantStart = 1'b0;
    if(when_StateMachine_l237_1) begin
      token_wantStart = 1'b1;
    end
    if(when_StateMachine_l253_1) begin
      token_wantStart = 1'b1;
    end
  end

  always @(*) begin
    token_wantKill = 1'b0;
    if(unscheduleAll_fire) begin
      token_wantKill = 1'b1;
    end
  end

  always @(*) begin
    token_pid = 4'bxxxx;
    case(sof_stateReg)
      sof_enumDef_FRAME_TX : begin
        token_pid = 4'b0101;
      end
      sof_enumDef_FRAME_NUMBER_CMD : begin
      end
      sof_enumDef_FRAME_NUMBER_RSP : begin
      end
      default : begin
      end
    endcase
    case(endpoint_stateReg)
      endpoint_enumDef_ED_READ_CMD : begin
      end
      endpoint_enumDef_ED_READ_RSP : begin
      end
      endpoint_enumDef_ED_ANALYSE : begin
      end
      endpoint_enumDef_TD_READ_CMD : begin
      end
      endpoint_enumDef_TD_READ_RSP : begin
      end
      endpoint_enumDef_TD_READ_DELAY : begin
      end
      endpoint_enumDef_TD_ANALYSE : begin
      end
      endpoint_enumDef_TD_CHECK_TIME : begin
      end
      endpoint_enumDef_BUFFER_READ : begin
      end
      endpoint_enumDef_TOKEN : begin
        case(endpoint_tockenType)
          2'b00 : begin
            token_pid = 4'b1101;
          end
          2'b01 : begin
            token_pid = 4'b0001;
          end
          2'b10 : begin
            token_pid = 4'b1001;
          end
          default : begin
          end
        endcase
      end
      endpoint_enumDef_DATA_TX : begin
      end
      endpoint_enumDef_DATA_RX : begin
      end
      endpoint_enumDef_DATA_RX_VALIDATE : begin
      end
      endpoint_enumDef_ACK_RX : begin
      end
      endpoint_enumDef_ACK_TX_0 : begin
      end
      endpoint_enumDef_ACK_TX_1 : begin
      end
      endpoint_enumDef_ACK_TX_EOP : begin
      end
      endpoint_enumDef_DATA_RX_WAIT_DMA : begin
      end
      endpoint_enumDef_UPDATE_TD_PROCESS : begin
      end
      endpoint_enumDef_UPDATE_TD_CMD : begin
      end
      endpoint_enumDef_UPDATE_ED_CMD : begin
      end
      endpoint_enumDef_UPDATE_SYNC : begin
      end
      endpoint_enumDef_ABORD : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    token_data = 11'bxxxxxxxxxxx;
    case(sof_stateReg)
      sof_enumDef_FRAME_TX : begin
        token_data = _zz_token_data[10:0];
      end
      sof_enumDef_FRAME_NUMBER_CMD : begin
      end
      sof_enumDef_FRAME_NUMBER_RSP : begin
      end
      default : begin
      end
    endcase
    case(endpoint_stateReg)
      endpoint_enumDef_ED_READ_CMD : begin
      end
      endpoint_enumDef_ED_READ_RSP : begin
      end
      endpoint_enumDef_ED_ANALYSE : begin
      end
      endpoint_enumDef_TD_READ_CMD : begin
      end
      endpoint_enumDef_TD_READ_RSP : begin
      end
      endpoint_enumDef_TD_READ_DELAY : begin
      end
      endpoint_enumDef_TD_ANALYSE : begin
      end
      endpoint_enumDef_TD_CHECK_TIME : begin
      end
      endpoint_enumDef_BUFFER_READ : begin
      end
      endpoint_enumDef_TOKEN : begin
        token_data = {endpoint_ED_EN,endpoint_ED_FA};
      end
      endpoint_enumDef_DATA_TX : begin
      end
      endpoint_enumDef_DATA_RX : begin
      end
      endpoint_enumDef_DATA_RX_VALIDATE : begin
      end
      endpoint_enumDef_ACK_RX : begin
      end
      endpoint_enumDef_ACK_TX_0 : begin
      end
      endpoint_enumDef_ACK_TX_1 : begin
      end
      endpoint_enumDef_ACK_TX_EOP : begin
      end
      endpoint_enumDef_DATA_RX_WAIT_DMA : begin
      end
      endpoint_enumDef_UPDATE_TD_PROCESS : begin
      end
      endpoint_enumDef_UPDATE_TD_CMD : begin
      end
      endpoint_enumDef_UPDATE_ED_CMD : begin
      end
      endpoint_enumDef_UPDATE_SYNC : begin
      end
      endpoint_enumDef_ABORD : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    token_crc5_io_flush = 1'b0;
    if(when_StateMachine_l237) begin
      token_crc5_io_flush = 1'b1;
    end
  end

  always @(*) begin
    token_crc5_io_input_valid = 1'b0;
    case(token_stateReg)
      token_enumDef_INIT : begin
        token_crc5_io_input_valid = 1'b1;
      end
      token_enumDef_PID : begin
      end
      token_enumDef_B1 : begin
      end
      token_enumDef_B2 : begin
      end
      token_enumDef_EOP : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    dataTx_wantExit = 1'b0;
    case(dataTx_stateReg)
      dataTx_enumDef_PID : begin
      end
      dataTx_enumDef_DATA : begin
      end
      dataTx_enumDef_CRC_0 : begin
      end
      dataTx_enumDef_CRC_1 : begin
      end
      dataTx_enumDef_EOP : begin
        if(io_phy_txEop) begin
          dataTx_wantExit = 1'b1;
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    dataTx_wantStart = 1'b0;
    if(when_StateMachine_l253_2) begin
      dataTx_wantStart = 1'b1;
    end
  end

  always @(*) begin
    dataTx_wantKill = 1'b0;
    if(unscheduleAll_fire) begin
      dataTx_wantKill = 1'b1;
    end
  end

  always @(*) begin
    dataTx_pid = 4'bxxxx;
    case(endpoint_stateReg)
      endpoint_enumDef_ED_READ_CMD : begin
      end
      endpoint_enumDef_ED_READ_RSP : begin
      end
      endpoint_enumDef_ED_ANALYSE : begin
      end
      endpoint_enumDef_TD_READ_CMD : begin
      end
      endpoint_enumDef_TD_READ_RSP : begin
      end
      endpoint_enumDef_TD_READ_DELAY : begin
      end
      endpoint_enumDef_TD_ANALYSE : begin
      end
      endpoint_enumDef_TD_CHECK_TIME : begin
      end
      endpoint_enumDef_BUFFER_READ : begin
      end
      endpoint_enumDef_TOKEN : begin
      end
      endpoint_enumDef_DATA_TX : begin
        dataTx_pid = {endpoint_dataPhase,3'b011};
      end
      endpoint_enumDef_DATA_RX : begin
      end
      endpoint_enumDef_DATA_RX_VALIDATE : begin
      end
      endpoint_enumDef_ACK_RX : begin
      end
      endpoint_enumDef_ACK_TX_0 : begin
      end
      endpoint_enumDef_ACK_TX_1 : begin
      end
      endpoint_enumDef_ACK_TX_EOP : begin
      end
      endpoint_enumDef_DATA_RX_WAIT_DMA : begin
      end
      endpoint_enumDef_UPDATE_TD_PROCESS : begin
      end
      endpoint_enumDef_UPDATE_TD_CMD : begin
      end
      endpoint_enumDef_UPDATE_ED_CMD : begin
      end
      endpoint_enumDef_UPDATE_SYNC : begin
      end
      endpoint_enumDef_ABORD : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    dataTx_data_valid = 1'b0;
    if(endpoint_dmaLogic_toUsb_run) begin
      if(endpoint_dmaLogic_storage_readRsp_valid) begin
        dataTx_data_valid = 1'b1;
      end
    end
  end

  always @(*) begin
    dataTx_data_payload_last = 1'bx;
    if(endpoint_dmaLogic_toUsb_run) begin
      dataTx_data_payload_last = endpoint_dmaLogic_byteCtx_last;
    end
  end

  always @(*) begin
    dataTx_data_payload_fragment = 8'bxxxxxxxx;
    if(endpoint_dmaLogic_toUsb_run) begin
      dataTx_data_payload_fragment = _zz_dataTx_data_payload_fragment;
    end
  end

  always @(*) begin
    dataTx_data_ready = 1'b0;
    case(dataTx_stateReg)
      dataTx_enumDef_PID : begin
      end
      dataTx_enumDef_DATA : begin
        if(io_phy_tx_ready) begin
          dataTx_data_ready = 1'b1;
        end
      end
      dataTx_enumDef_CRC_0 : begin
      end
      dataTx_enumDef_CRC_1 : begin
      end
      dataTx_enumDef_EOP : begin
      end
      default : begin
      end
    endcase
  end

  assign dataTx_data_fire = (dataTx_data_valid && dataTx_data_ready);
  always @(*) begin
    dataTx_crc16_io_flush = 1'b0;
    case(dataTx_stateReg)
      dataTx_enumDef_PID : begin
        dataTx_crc16_io_flush = 1'b1;
      end
      dataTx_enumDef_DATA : begin
      end
      dataTx_enumDef_CRC_0 : begin
      end
      dataTx_enumDef_CRC_1 : begin
      end
      dataTx_enumDef_EOP : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    rxTimer_clear = 1'b0;
    if(io_phy_rx_active) begin
      rxTimer_clear = 1'b1;
    end
    if(when_StateMachine_l253) begin
      rxTimer_clear = 1'b1;
    end
    if(when_StateMachine_l253_4) begin
      rxTimer_clear = 1'b1;
    end
  end

  assign rxTimer_rxTimeout = (rxTimer_counter == (rxTimer_lowSpeed ? 8'hbf : 8'h17));
  assign rxTimer_ackTx = (rxTimer_counter == _zz_rxTimer_ackTx);
  assign rxPidOk = (io_phy_rx_flow_payload_data[3 : 0] == (~ io_phy_rx_flow_payload_data[7 : 4]));
  assign _zz_2 = io_phy_rx_flow_valid;
  assign _zz_dataRx_pid = io_phy_rx_flow_payload_data;
  assign when_Misc_l87 = (io_phy_rx_flow_valid && io_phy_rx_flow_payload_stuffingError);
  always @(*) begin
    dataRx_wantExit = 1'b0;
    case(dataRx_stateReg)
      dataRx_enumDef_IDLE : begin
        if(!io_phy_rx_active) begin
          if(rxTimer_rxTimeout) begin
            dataRx_wantExit = 1'b1;
          end
        end
      end
      dataRx_enumDef_PID : begin
        if(!_zz_2) begin
          if(when_Misc_l64) begin
            dataRx_wantExit = 1'b1;
          end
        end
      end
      dataRx_enumDef_DATA : begin
        if(when_Misc_l70) begin
          dataRx_wantExit = 1'b1;
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    dataRx_wantStart = 1'b0;
    if(when_StateMachine_l253_3) begin
      dataRx_wantStart = 1'b1;
    end
  end

  always @(*) begin
    dataRx_wantKill = 1'b0;
    if(unscheduleAll_fire) begin
      dataRx_wantKill = 1'b1;
    end
  end

  assign dataRx_history_0 = _zz_dataRx_history_0;
  assign dataRx_history_1 = _zz_dataRx_history_1;
  assign dataRx_hasError = (|{dataRx_crcError,{dataRx_pidError,{dataRx_stuffingError,dataRx_notResponding}}});
  always @(*) begin
    dataRx_data_valid = 1'b0;
    case(dataRx_stateReg)
      dataRx_enumDef_IDLE : begin
      end
      dataRx_enumDef_PID : begin
      end
      dataRx_enumDef_DATA : begin
        if(!when_Misc_l70) begin
          if(_zz_2) begin
            if(when_Misc_l78) begin
              dataRx_data_valid = 1'b1;
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  assign dataRx_data_payload = dataRx_history_1;
  always @(*) begin
    dataRx_crc16_io_input_valid = 1'b0;
    case(dataRx_stateReg)
      dataRx_enumDef_IDLE : begin
      end
      dataRx_enumDef_PID : begin
      end
      dataRx_enumDef_DATA : begin
        if(!when_Misc_l70) begin
          if(_zz_2) begin
            dataRx_crc16_io_input_valid = 1'b1;
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    dataRx_crc16_io_flush = 1'b0;
    case(dataRx_stateReg)
      dataRx_enumDef_IDLE : begin
      end
      dataRx_enumDef_PID : begin
        dataRx_crc16_io_flush = 1'b1;
      end
      dataRx_enumDef_DATA : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    sof_wantExit = 1'b0;
    case(sof_stateReg)
      sof_enumDef_FRAME_TX : begin
      end
      sof_enumDef_FRAME_NUMBER_CMD : begin
      end
      sof_enumDef_FRAME_NUMBER_RSP : begin
        if(ioDma_rsp_valid) begin
          sof_wantExit = 1'b1;
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    sof_wantStart = 1'b0;
    if(when_StateMachine_l253_6) begin
      sof_wantStart = 1'b1;
    end
  end

  always @(*) begin
    sof_wantKill = 1'b0;
    if(unscheduleAll_fire) begin
      sof_wantKill = 1'b1;
    end
  end

  always @(*) begin
    priority_tick = 1'b0;
    case(endpoint_stateReg)
      endpoint_enumDef_ED_READ_CMD : begin
      end
      endpoint_enumDef_ED_READ_RSP : begin
      end
      endpoint_enumDef_ED_ANALYSE : begin
      end
      endpoint_enumDef_TD_READ_CMD : begin
      end
      endpoint_enumDef_TD_READ_RSP : begin
      end
      endpoint_enumDef_TD_READ_DELAY : begin
      end
      endpoint_enumDef_TD_ANALYSE : begin
      end
      endpoint_enumDef_TD_CHECK_TIME : begin
      end
      endpoint_enumDef_BUFFER_READ : begin
      end
      endpoint_enumDef_TOKEN : begin
      end
      endpoint_enumDef_DATA_TX : begin
      end
      endpoint_enumDef_DATA_RX : begin
      end
      endpoint_enumDef_DATA_RX_VALIDATE : begin
      end
      endpoint_enumDef_ACK_RX : begin
      end
      endpoint_enumDef_ACK_TX_0 : begin
      end
      endpoint_enumDef_ACK_TX_1 : begin
      end
      endpoint_enumDef_ACK_TX_EOP : begin
      end
      endpoint_enumDef_DATA_RX_WAIT_DMA : begin
      end
      endpoint_enumDef_UPDATE_TD_PROCESS : begin
      end
      endpoint_enumDef_UPDATE_TD_CMD : begin
      end
      endpoint_enumDef_UPDATE_ED_CMD : begin
      end
      endpoint_enumDef_UPDATE_SYNC : begin
        if(dmaCtx_pendingEmpty) begin
          if(when_UsbOhci_l1473) begin
            priority_tick = 1'b1;
          end
        end
      end
      endpoint_enumDef_ABORD : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    priority_skip = 1'b0;
    if(priority_tick) begin
      if(when_UsbOhci_l651) begin
        priority_skip = 1'b1;
      end
    end
    case(operational_stateReg)
      operational_enumDef_SOF : begin
      end
      operational_enumDef_ARBITER : begin
        if(!operational_askExit) begin
          if(!frame_limitHit) begin
            if(!when_UsbOhci_l1542) begin
              priority_skip = 1'b1;
              if(priority_bulk) begin
                if(operational_allowBulk) begin
                  if(reg_hcBulkCurrentED_isZero) begin
                    if(reg_hcCommandStatus_BLF) begin
                      priority_skip = 1'b0;
                    end
                  end else begin
                    priority_skip = 1'b0;
                  end
                end
              end else begin
                if(operational_allowControl) begin
                  if(reg_hcControlCurrentED_isZero) begin
                    if(reg_hcCommandStatus_CLF) begin
                      priority_skip = 1'b0;
                    end
                  end else begin
                    priority_skip = 1'b0;
                  end
                end
              end
            end
          end
        end
      end
      operational_enumDef_END_POINT : begin
      end
      operational_enumDef_PERIODIC_HEAD_CMD : begin
      end
      operational_enumDef_PERIODIC_HEAD_RSP : begin
      end
      operational_enumDef_WAIT_SOF : begin
      end
      default : begin
      end
    endcase
  end

  assign when_UsbOhci_l651 = (priority_bulk || (priority_counter == reg_hcControl_CBSR));
  always @(*) begin
    interruptDelay_tick = 1'b0;
    case(sof_stateReg)
      sof_enumDef_FRAME_TX : begin
      end
      sof_enumDef_FRAME_NUMBER_CMD : begin
      end
      sof_enumDef_FRAME_NUMBER_RSP : begin
        if(ioDma_rsp_valid) begin
          interruptDelay_tick = 1'b1;
        end
      end
      default : begin
      end
    endcase
  end

  assign interruptDelay_done = (interruptDelay_counter == 3'b000);
  assign interruptDelay_disabled = (interruptDelay_counter == 3'b111);
  always @(*) begin
    interruptDelay_disable = 1'b0;
    case(sof_stateReg)
      sof_enumDef_FRAME_TX : begin
      end
      sof_enumDef_FRAME_NUMBER_CMD : begin
      end
      sof_enumDef_FRAME_NUMBER_RSP : begin
        if(ioDma_rsp_valid) begin
          if(sof_doInterruptDelay) begin
            interruptDelay_disable = 1'b1;
          end
        end
      end
      default : begin
      end
    endcase
    if(when_StateMachine_l237_3) begin
      interruptDelay_disable = 1'b1;
    end
  end

  always @(*) begin
    interruptDelay_load_valid = 1'b0;
    case(endpoint_stateReg)
      endpoint_enumDef_ED_READ_CMD : begin
      end
      endpoint_enumDef_ED_READ_RSP : begin
      end
      endpoint_enumDef_ED_ANALYSE : begin
      end
      endpoint_enumDef_TD_READ_CMD : begin
      end
      endpoint_enumDef_TD_READ_RSP : begin
      end
      endpoint_enumDef_TD_READ_DELAY : begin
      end
      endpoint_enumDef_TD_ANALYSE : begin
      end
      endpoint_enumDef_TD_CHECK_TIME : begin
      end
      endpoint_enumDef_BUFFER_READ : begin
      end
      endpoint_enumDef_TOKEN : begin
      end
      endpoint_enumDef_DATA_TX : begin
      end
      endpoint_enumDef_DATA_RX : begin
      end
      endpoint_enumDef_DATA_RX_VALIDATE : begin
      end
      endpoint_enumDef_ACK_RX : begin
      end
      endpoint_enumDef_ACK_TX_0 : begin
      end
      endpoint_enumDef_ACK_TX_1 : begin
      end
      endpoint_enumDef_ACK_TX_EOP : begin
      end
      endpoint_enumDef_DATA_RX_WAIT_DMA : begin
      end
      endpoint_enumDef_UPDATE_TD_PROCESS : begin
      end
      endpoint_enumDef_UPDATE_TD_CMD : begin
      end
      endpoint_enumDef_UPDATE_ED_CMD : begin
      end
      endpoint_enumDef_UPDATE_SYNC : begin
        if(dmaCtx_pendingEmpty) begin
          if(endpoint_TD_retire) begin
            interruptDelay_load_valid = 1'b1;
          end
        end
      end
      endpoint_enumDef_ABORD : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    interruptDelay_load_payload = 3'bxxx;
    case(endpoint_stateReg)
      endpoint_enumDef_ED_READ_CMD : begin
      end
      endpoint_enumDef_ED_READ_RSP : begin
      end
      endpoint_enumDef_ED_ANALYSE : begin
      end
      endpoint_enumDef_TD_READ_CMD : begin
      end
      endpoint_enumDef_TD_READ_RSP : begin
      end
      endpoint_enumDef_TD_READ_DELAY : begin
      end
      endpoint_enumDef_TD_ANALYSE : begin
      end
      endpoint_enumDef_TD_CHECK_TIME : begin
      end
      endpoint_enumDef_BUFFER_READ : begin
      end
      endpoint_enumDef_TOKEN : begin
      end
      endpoint_enumDef_DATA_TX : begin
      end
      endpoint_enumDef_DATA_RX : begin
      end
      endpoint_enumDef_DATA_RX_VALIDATE : begin
      end
      endpoint_enumDef_ACK_RX : begin
      end
      endpoint_enumDef_ACK_TX_0 : begin
      end
      endpoint_enumDef_ACK_TX_1 : begin
      end
      endpoint_enumDef_ACK_TX_EOP : begin
      end
      endpoint_enumDef_DATA_RX_WAIT_DMA : begin
      end
      endpoint_enumDef_UPDATE_TD_PROCESS : begin
      end
      endpoint_enumDef_UPDATE_TD_CMD : begin
      end
      endpoint_enumDef_UPDATE_ED_CMD : begin
      end
      endpoint_enumDef_UPDATE_SYNC : begin
        if(dmaCtx_pendingEmpty) begin
          if(endpoint_TD_retire) begin
            interruptDelay_load_payload = endpoint_TD_DI;
          end
        end
      end
      endpoint_enumDef_ABORD : begin
      end
      default : begin
      end
    endcase
  end

  assign when_UsbOhci_l673 = ((interruptDelay_tick && (! interruptDelay_done)) && (! interruptDelay_disabled));
  assign when_UsbOhci_l677 = (interruptDelay_load_valid && (interruptDelay_load_payload < interruptDelay_counter));
  always @(*) begin
    endpoint_wantExit = 1'b0;
    case(endpoint_stateReg)
      endpoint_enumDef_ED_READ_CMD : begin
      end
      endpoint_enumDef_ED_READ_RSP : begin
      end
      endpoint_enumDef_ED_ANALYSE : begin
        if(when_UsbOhci_l849) begin
          endpoint_wantExit = 1'b1;
        end
      end
      endpoint_enumDef_TD_READ_CMD : begin
      end
      endpoint_enumDef_TD_READ_RSP : begin
      end
      endpoint_enumDef_TD_READ_DELAY : begin
      end
      endpoint_enumDef_TD_ANALYSE : begin
      end
      endpoint_enumDef_TD_CHECK_TIME : begin
      end
      endpoint_enumDef_BUFFER_READ : begin
      end
      endpoint_enumDef_TOKEN : begin
      end
      endpoint_enumDef_DATA_TX : begin
      end
      endpoint_enumDef_DATA_RX : begin
      end
      endpoint_enumDef_DATA_RX_VALIDATE : begin
      end
      endpoint_enumDef_ACK_RX : begin
      end
      endpoint_enumDef_ACK_TX_0 : begin
      end
      endpoint_enumDef_ACK_TX_1 : begin
      end
      endpoint_enumDef_ACK_TX_EOP : begin
      end
      endpoint_enumDef_DATA_RX_WAIT_DMA : begin
      end
      endpoint_enumDef_UPDATE_TD_PROCESS : begin
      end
      endpoint_enumDef_UPDATE_TD_CMD : begin
      end
      endpoint_enumDef_UPDATE_ED_CMD : begin
      end
      endpoint_enumDef_UPDATE_SYNC : begin
        if(dmaCtx_pendingEmpty) begin
          endpoint_wantExit = 1'b1;
        end
      end
      endpoint_enumDef_ABORD : begin
        endpoint_wantExit = 1'b1;
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    endpoint_wantStart = 1'b0;
    case(operational_stateReg)
      operational_enumDef_SOF : begin
      end
      operational_enumDef_ARBITER : begin
        if(!operational_askExit) begin
          if(!frame_limitHit) begin
            if(when_UsbOhci_l1542) begin
              if(!when_UsbOhci_l1543) begin
                if(!reg_hcPeriodCurrentED_isZero) begin
                  endpoint_wantStart = 1'b1;
                end
              end
            end else begin
              if(priority_bulk) begin
                if(operational_allowBulk) begin
                  if(!reg_hcBulkCurrentED_isZero) begin
                    endpoint_wantStart = 1'b1;
                  end
                end
              end else begin
                if(operational_allowControl) begin
                  if(!reg_hcControlCurrentED_isZero) begin
                    endpoint_wantStart = 1'b1;
                  end
                end
              end
            end
          end
        end
      end
      operational_enumDef_END_POINT : begin
      end
      operational_enumDef_PERIODIC_HEAD_CMD : begin
      end
      operational_enumDef_PERIODIC_HEAD_RSP : begin
      end
      operational_enumDef_WAIT_SOF : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    endpoint_wantKill = 1'b0;
    if(unscheduleAll_fire) begin
      endpoint_wantKill = 1'b1;
    end
  end

  assign endpoint_ED_FA = endpoint_ED_words_0[6 : 0];
  assign endpoint_ED_EN = endpoint_ED_words_0[10 : 7];
  assign endpoint_ED_D = endpoint_ED_words_0[12 : 11];
  assign endpoint_ED_S = endpoint_ED_words_0[13];
  assign endpoint_ED_K = endpoint_ED_words_0[14];
  assign endpoint_ED_F = endpoint_ED_words_0[15];
  assign endpoint_ED_MPS = endpoint_ED_words_0[26 : 16];
  assign endpoint_ED_tailP = endpoint_ED_words_1[31 : 4];
  assign endpoint_ED_H = endpoint_ED_words_2[0];
  assign endpoint_ED_C = endpoint_ED_words_2[1];
  assign endpoint_ED_headP = endpoint_ED_words_2[31 : 4];
  assign endpoint_ED_nextED = endpoint_ED_words_3[31 : 4];
  assign endpoint_ED_tdEmpty = (endpoint_ED_tailP == endpoint_ED_headP);
  assign endpoint_ED_isFs = (! endpoint_ED_S);
  assign endpoint_ED_isoOut = endpoint_ED_D[0];
  assign when_UsbOhci_l738 = (! (endpoint_stateReg == endpoint_enumDef_BOOT));
  assign rxTimer_lowSpeed = endpoint_ED_S;
  assign endpoint_TD_address = ({4'd0,endpoint_ED_headP} <<< 3'd4);
  assign endpoint_TD_CC = endpoint_TD_words_0[31 : 28];
  assign endpoint_TD_EC = endpoint_TD_words_0[27 : 26];
  assign endpoint_TD_T = endpoint_TD_words_0[25 : 24];
  assign endpoint_TD_DI = endpoint_TD_words_0[23 : 21];
  assign endpoint_TD_DP = endpoint_TD_words_0[20 : 19];
  assign endpoint_TD_R = endpoint_TD_words_0[18];
  assign endpoint_TD_CBP = endpoint_TD_words_1[31 : 0];
  assign endpoint_TD_nextTD = endpoint_TD_words_2[31 : 4];
  assign endpoint_TD_BE = endpoint_TD_words_3[31 : 0];
  assign endpoint_TD_FC = endpoint_TD_words_0[26 : 24];
  assign endpoint_TD_SF = endpoint_TD_words_0[15 : 0];
  assign endpoint_TD_isoRelativeFrameNumber = (reg_hcFmNumber_FN - endpoint_TD_SF);
  assign endpoint_TD_tooEarly = endpoint_TD_isoRelativeFrameNumber[15];
  assign endpoint_TD_isoFrameNumber = endpoint_TD_isoRelativeFrameNumber[2 : 0];
  assign endpoint_TD_isoOverrun = ((! endpoint_TD_tooEarly) && (_zz_endpoint_TD_isoOverrun < endpoint_TD_isoRelativeFrameNumber));
  assign endpoint_TD_isoLast = (((! endpoint_TD_isoOverrun) && (! endpoint_TD_tooEarly)) && (endpoint_TD_isoFrameNumber == endpoint_TD_FC));
  assign endpoint_TD_isSinglePage = (endpoint_TD_CBP[31 : 12] == endpoint_TD_BE[31 : 12]);
  assign endpoint_TD_firstOffset = (endpoint_ED_F ? endpoint_TD_isoBase : _zz_endpoint_TD_firstOffset);
  assign endpoint_TD_allowRounding = ((! endpoint_ED_F) && endpoint_TD_R);
  assign endpoint_TD_TNext = (endpoint_TD_dataPhaseUpdate ? {1'b1,(! endpoint_dataPhase)} : endpoint_TD_T);
  assign endpoint_TD_dataPhaseNext = (endpoint_dataPhase ^ endpoint_TD_dataPhaseUpdate);
  assign endpoint_TD_dataPid = (endpoint_dataPhase ? 4'b1011 : 4'b0011);
  assign endpoint_TD_dataPidWrong = (endpoint_dataPhase ? 4'b0011 : 4'b1011);
  always @(*) begin
    endpoint_TD_clear = 1'b0;
    case(endpoint_stateReg)
      endpoint_enumDef_ED_READ_CMD : begin
      end
      endpoint_enumDef_ED_READ_RSP : begin
      end
      endpoint_enumDef_ED_ANALYSE : begin
      end
      endpoint_enumDef_TD_READ_CMD : begin
        endpoint_TD_clear = 1'b1;
      end
      endpoint_enumDef_TD_READ_RSP : begin
      end
      endpoint_enumDef_TD_READ_DELAY : begin
      end
      endpoint_enumDef_TD_ANALYSE : begin
      end
      endpoint_enumDef_TD_CHECK_TIME : begin
      end
      endpoint_enumDef_BUFFER_READ : begin
      end
      endpoint_enumDef_TOKEN : begin
      end
      endpoint_enumDef_DATA_TX : begin
      end
      endpoint_enumDef_DATA_RX : begin
      end
      endpoint_enumDef_DATA_RX_VALIDATE : begin
      end
      endpoint_enumDef_ACK_RX : begin
      end
      endpoint_enumDef_ACK_TX_0 : begin
      end
      endpoint_enumDef_ACK_TX_1 : begin
      end
      endpoint_enumDef_ACK_TX_EOP : begin
      end
      endpoint_enumDef_DATA_RX_WAIT_DMA : begin
      end
      endpoint_enumDef_UPDATE_TD_PROCESS : begin
      end
      endpoint_enumDef_UPDATE_TD_CMD : begin
      end
      endpoint_enumDef_UPDATE_ED_CMD : begin
      end
      endpoint_enumDef_UPDATE_SYNC : begin
      end
      endpoint_enumDef_ABORD : begin
      end
      default : begin
      end
    endcase
  end

  assign endpoint_tockenType = ((endpoint_ED_D[0] != endpoint_ED_D[1]) ? endpoint_ED_D : endpoint_TD_DP);
  assign endpoint_isIn = (endpoint_tockenType == 2'b10);
  always @(*) begin
    endpoint_applyNextED = 1'b0;
    case(endpoint_stateReg)
      endpoint_enumDef_ED_READ_CMD : begin
      end
      endpoint_enumDef_ED_READ_RSP : begin
      end
      endpoint_enumDef_ED_ANALYSE : begin
        if(when_UsbOhci_l849) begin
          endpoint_applyNextED = 1'b1;
        end
      end
      endpoint_enumDef_TD_READ_CMD : begin
      end
      endpoint_enumDef_TD_READ_RSP : begin
      end
      endpoint_enumDef_TD_READ_DELAY : begin
      end
      endpoint_enumDef_TD_ANALYSE : begin
      end
      endpoint_enumDef_TD_CHECK_TIME : begin
      end
      endpoint_enumDef_BUFFER_READ : begin
      end
      endpoint_enumDef_TOKEN : begin
      end
      endpoint_enumDef_DATA_TX : begin
      end
      endpoint_enumDef_DATA_RX : begin
      end
      endpoint_enumDef_DATA_RX_VALIDATE : begin
      end
      endpoint_enumDef_ACK_RX : begin
      end
      endpoint_enumDef_ACK_TX_0 : begin
      end
      endpoint_enumDef_ACK_TX_1 : begin
      end
      endpoint_enumDef_ACK_TX_EOP : begin
      end
      endpoint_enumDef_DATA_RX_WAIT_DMA : begin
      end
      endpoint_enumDef_UPDATE_TD_PROCESS : begin
      end
      endpoint_enumDef_UPDATE_TD_CMD : begin
      end
      endpoint_enumDef_UPDATE_ED_CMD : begin
      end
      endpoint_enumDef_UPDATE_SYNC : begin
        if(dmaCtx_pendingEmpty) begin
          if(when_UsbOhci_l1470) begin
            endpoint_applyNextED = 1'b1;
          end
        end
      end
      endpoint_enumDef_ABORD : begin
      end
      default : begin
      end
    endcase
  end

  assign endpoint_currentAddressFull = {(endpoint_currentAddress[12] ? endpoint_TD_BE[31 : 12] : endpoint_TD_CBP[31 : 12]),endpoint_currentAddress[11 : 0]};
  assign endpoint_currentAddressBmb = ({6'd0,_zz_endpoint_currentAddressBmb} <<< 3'd6);
  assign endpoint_transactionSizeMinusOne = (_zz_endpoint_transactionSizeMinusOne - endpoint_currentAddress);
  assign endpoint_transactionSize = (endpoint_transactionSizeMinusOne + 14'h0001);
  assign endpoint_dataDone = (endpoint_zeroLength || (_zz_endpoint_dataDone < endpoint_currentAddress));
  always @(*) begin
    endpoint_dmaLogic_wantExit = 1'b0;
    case(endpoint_dmaLogic_stateReg)
      endpoint_dmaLogic_enumDef_INIT : begin
      end
      endpoint_dmaLogic_enumDef_TO_USB : begin
      end
      endpoint_dmaLogic_enumDef_FROM_USB : begin
      end
      endpoint_dmaLogic_enumDef_VALIDATION : begin
      end
      endpoint_dmaLogic_enumDef_CALC_CMD : begin
        if(endpoint_isIn) begin
          if(when_UsbOhci_l1047) begin
            endpoint_dmaLogic_wantExit = 1'b1;
          end
        end
      end
      endpoint_dmaLogic_enumDef_READ_CMD : begin
      end
      endpoint_dmaLogic_enumDef_WRITE_CMD : begin
      end
      default : begin
      end
    endcase
    if(endpoint_dmaLogic_toUsb_run) begin
      if(endpoint_dmaLogic_storage_readRsp_valid) begin
        if(dataTx_data_ready) begin
          if(endpoint_dmaLogic_byteCtx_last) begin
            endpoint_dmaLogic_wantExit = 1'b1;
          end
        end
      end
    end
  end

  always @(*) begin
    endpoint_dmaLogic_wantStart = 1'b0;
    case(endpoint_stateReg)
      endpoint_enumDef_ED_READ_CMD : begin
      end
      endpoint_enumDef_ED_READ_RSP : begin
      end
      endpoint_enumDef_ED_ANALYSE : begin
      end
      endpoint_enumDef_TD_READ_CMD : begin
      end
      endpoint_enumDef_TD_READ_RSP : begin
      end
      endpoint_enumDef_TD_READ_DELAY : begin
      end
      endpoint_enumDef_TD_ANALYSE : begin
      end
      endpoint_enumDef_TD_CHECK_TIME : begin
        if(!endpoint_timeCheck) begin
          if(!when_UsbOhci_l1173) begin
            endpoint_dmaLogic_wantStart = 1'b1;
          end
        end
      end
      endpoint_enumDef_BUFFER_READ : begin
      end
      endpoint_enumDef_TOKEN : begin
      end
      endpoint_enumDef_DATA_TX : begin
      end
      endpoint_enumDef_DATA_RX : begin
      end
      endpoint_enumDef_DATA_RX_VALIDATE : begin
      end
      endpoint_enumDef_ACK_RX : begin
      end
      endpoint_enumDef_ACK_TX_0 : begin
      end
      endpoint_enumDef_ACK_TX_1 : begin
      end
      endpoint_enumDef_ACK_TX_EOP : begin
      end
      endpoint_enumDef_DATA_RX_WAIT_DMA : begin
      end
      endpoint_enumDef_UPDATE_TD_PROCESS : begin
      end
      endpoint_enumDef_UPDATE_TD_CMD : begin
      end
      endpoint_enumDef_UPDATE_ED_CMD : begin
      end
      endpoint_enumDef_UPDATE_SYNC : begin
      end
      endpoint_enumDef_ABORD : begin
      end
      default : begin
      end
    endcase
    if(when_StateMachine_l253_3) begin
      endpoint_dmaLogic_wantStart = 1'b1;
    end
  end

  always @(*) begin
    endpoint_dmaLogic_wantKill = 1'b0;
    case(endpoint_stateReg)
      endpoint_enumDef_ED_READ_CMD : begin
      end
      endpoint_enumDef_ED_READ_RSP : begin
      end
      endpoint_enumDef_ED_ANALYSE : begin
      end
      endpoint_enumDef_TD_READ_CMD : begin
      end
      endpoint_enumDef_TD_READ_RSP : begin
      end
      endpoint_enumDef_TD_READ_DELAY : begin
      end
      endpoint_enumDef_TD_ANALYSE : begin
      end
      endpoint_enumDef_TD_CHECK_TIME : begin
      end
      endpoint_enumDef_BUFFER_READ : begin
        if(endpoint_dmaLogic_toUsb_run) begin
          if(endpoint_timeCheck) begin
            endpoint_dmaLogic_wantKill = 1'b1;
          end
        end
      end
      endpoint_enumDef_TOKEN : begin
      end
      endpoint_enumDef_DATA_TX : begin
      end
      endpoint_enumDef_DATA_RX : begin
      end
      endpoint_enumDef_DATA_RX_VALIDATE : begin
      end
      endpoint_enumDef_ACK_RX : begin
      end
      endpoint_enumDef_ACK_TX_0 : begin
      end
      endpoint_enumDef_ACK_TX_1 : begin
      end
      endpoint_enumDef_ACK_TX_EOP : begin
      end
      endpoint_enumDef_DATA_RX_WAIT_DMA : begin
      end
      endpoint_enumDef_UPDATE_TD_PROCESS : begin
      end
      endpoint_enumDef_UPDATE_TD_CMD : begin
      end
      endpoint_enumDef_UPDATE_ED_CMD : begin
      end
      endpoint_enumDef_UPDATE_SYNC : begin
      end
      endpoint_enumDef_ABORD : begin
      end
      default : begin
      end
    endcase
    if(unscheduleAll_fire) begin
      endpoint_dmaLogic_wantKill = 1'b1;
    end
  end

  always @(*) begin
    endpoint_dmaLogic_storage_readCmd_valid = 1'b0;
    case(endpoint_dmaLogic_stateReg)
      endpoint_dmaLogic_enumDef_INIT : begin
      end
      endpoint_dmaLogic_enumDef_TO_USB : begin
      end
      endpoint_dmaLogic_enumDef_FROM_USB : begin
      end
      endpoint_dmaLogic_enumDef_VALIDATION : begin
      end
      endpoint_dmaLogic_enumDef_CALC_CMD : begin
      end
      endpoint_dmaLogic_enumDef_READ_CMD : begin
      end
      endpoint_dmaLogic_enumDef_WRITE_CMD : begin
        if(when_UsbOhci_l1093) begin
          endpoint_dmaLogic_storage_readCmd_valid = 1'b1;
        end
      end
      default : begin
      end
    endcase
    if(endpoint_dmaLogic_toUsb_run) begin
      endpoint_dmaLogic_storage_readCmd_valid = 1'b1;
    end
  end

  always @(*) begin
    endpoint_dmaLogic_storage_readCmd_payload = 6'bxxxxxx;
    case(endpoint_dmaLogic_stateReg)
      endpoint_dmaLogic_enumDef_INIT : begin
      end
      endpoint_dmaLogic_enumDef_TO_USB : begin
      end
      endpoint_dmaLogic_enumDef_FROM_USB : begin
      end
      endpoint_dmaLogic_enumDef_VALIDATION : begin
      end
      endpoint_dmaLogic_enumDef_CALC_CMD : begin
      end
      endpoint_dmaLogic_enumDef_READ_CMD : begin
      end
      endpoint_dmaLogic_enumDef_WRITE_CMD : begin
        if(when_UsbOhci_l1093) begin
          endpoint_dmaLogic_storage_readCmd_payload = endpoint_dmaLogic_storage_readPtr[5:0];
        end
      end
      default : begin
      end
    endcase
    if(endpoint_dmaLogic_toUsb_run) begin
      endpoint_dmaLogic_storage_readCmd_payload = endpoint_dmaLogic_storage_readPtr[5:0];
    end
  end

  assign endpoint_dmaLogic_storage_readCmd_fire = (endpoint_dmaLogic_storage_readCmd_valid && endpoint_dmaLogic_storage_readCmd_ready);
  assign endpoint_dmaLogic_storage_readRsp_isFree = ((! endpoint_dmaLogic_storage_readRsp_valid) || endpoint_dmaLogic_storage_readRsp_ready);
  assign endpoint_dmaLogic_storage_readCmd_ready = endpoint_dmaLogic_storage_readRsp_isFree;
  assign endpoint_dmaLogic_storage_readRsp_valid = _zz_endpoint_dmaLogic_storage_readRsp_valid;
  assign endpoint_dmaLogic_storage_readRsp_payload = endpoint_dmaLogic_storage_ram_spinal_port0;
  always @(*) begin
    endpoint_dmaLogic_storage_readRsp_ready = (endpoint_dmaLogic_stateReg == endpoint_dmaLogic_enumDef_BOOT);
    case(endpoint_dmaLogic_stateReg)
      endpoint_dmaLogic_enumDef_INIT : begin
      end
      endpoint_dmaLogic_enumDef_TO_USB : begin
      end
      endpoint_dmaLogic_enumDef_FROM_USB : begin
      end
      endpoint_dmaLogic_enumDef_VALIDATION : begin
      end
      endpoint_dmaLogic_enumDef_CALC_CMD : begin
      end
      endpoint_dmaLogic_enumDef_READ_CMD : begin
      end
      endpoint_dmaLogic_enumDef_WRITE_CMD : begin
        if(ioDma_cmd_ready) begin
          endpoint_dmaLogic_storage_readRsp_ready = 1'b1;
        end
      end
      default : begin
      end
    endcase
    if(endpoint_dmaLogic_toUsb_run) begin
      if(endpoint_dmaLogic_storage_readRsp_valid) begin
        if(dataTx_data_ready) begin
          if(when_UsbOhci_l973) begin
            endpoint_dmaLogic_storage_readRsp_ready = 1'b1;
          end
        end
      end
    end
  end

  always @(*) begin
    endpoint_dmaLogic_storage_write_valid = 1'b0;
    if(when_UsbOhci_l937) begin
      endpoint_dmaLogic_storage_write_valid = 1'b1;
    end
    if(endpoint_dmaLogic_fromUsb_push) begin
      endpoint_dmaLogic_storage_write_valid = 1'b1;
    end
  end

  always @(*) begin
    endpoint_dmaLogic_storage_write_payload_address = 6'bxxxxxx;
    if(when_UsbOhci_l937) begin
      endpoint_dmaLogic_storage_write_payload_address = endpoint_dmaLogic_storage_writePtr[5:0];
    end
    if(endpoint_dmaLogic_fromUsb_push) begin
      endpoint_dmaLogic_storage_write_payload_address = endpoint_dmaLogic_storage_writePtr[5:0];
    end
  end

  always @(*) begin
    endpoint_dmaLogic_storage_write_payload_data = 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
    if(when_UsbOhci_l937) begin
      endpoint_dmaLogic_storage_write_payload_data = ioDma_rsp_payload_fragment_data;
    end
    if(endpoint_dmaLogic_fromUsb_push) begin
      endpoint_dmaLogic_storage_write_payload_data = endpoint_dmaLogic_fromUsb_buffer;
    end
  end

  assign _zz_endpoint_dmaLogic_storage_full = endpoint_dmaLogic_storage_readPtr[6 : 4];
  assign endpoint_dmaLogic_storage_full = ({(! _zz_endpoint_dmaLogic_storage_full[2]),_zz_endpoint_dmaLogic_storage_full[1 : 0]} == _zz_endpoint_dmaLogic_storage_full_1);
  always @(*) begin
    endpoint_dmaLogic_validated = 1'b0;
    case(endpoint_stateReg)
      endpoint_enumDef_ED_READ_CMD : begin
      end
      endpoint_enumDef_ED_READ_RSP : begin
      end
      endpoint_enumDef_ED_ANALYSE : begin
      end
      endpoint_enumDef_TD_READ_CMD : begin
      end
      endpoint_enumDef_TD_READ_RSP : begin
      end
      endpoint_enumDef_TD_READ_DELAY : begin
      end
      endpoint_enumDef_TD_ANALYSE : begin
      end
      endpoint_enumDef_TD_CHECK_TIME : begin
      end
      endpoint_enumDef_BUFFER_READ : begin
      end
      endpoint_enumDef_TOKEN : begin
      end
      endpoint_enumDef_DATA_TX : begin
      end
      endpoint_enumDef_DATA_RX : begin
      end
      endpoint_enumDef_DATA_RX_VALIDATE : begin
        endpoint_dmaLogic_validated = 1'b1;
      end
      endpoint_enumDef_ACK_RX : begin
      end
      endpoint_enumDef_ACK_TX_0 : begin
      end
      endpoint_enumDef_ACK_TX_1 : begin
      end
      endpoint_enumDef_ACK_TX_EOP : begin
      end
      endpoint_enumDef_DATA_RX_WAIT_DMA : begin
      end
      endpoint_enumDef_UPDATE_TD_PROCESS : begin
      end
      endpoint_enumDef_UPDATE_TD_CMD : begin
      end
      endpoint_enumDef_UPDATE_ED_CMD : begin
      end
      endpoint_enumDef_UPDATE_SYNC : begin
      end
      endpoint_enumDef_ABORD : begin
      end
      default : begin
      end
    endcase
  end

  assign endpoint_dmaLogic_lengthMax = (~ _zz_endpoint_dmaLogic_lengthMax);
  assign endpoint_dmaLogic_lengthCalc = _zz_endpoint_dmaLogic_lengthCalc[5:0];
  assign endpoint_dmaLogic_beatCount = _zz_endpoint_dmaLogic_beatCount[6 : 2];
  assign endpoint_dmaLogic_underflowError = (endpoint_dmaLogic_underflow && (! endpoint_TD_allowRounding));
  assign when_UsbOhci_l937 = (((! (endpoint_dmaLogic_stateReg == endpoint_dmaLogic_enumDef_BOOT)) && (! endpoint_isIn)) && ioDma_rsp_valid);
  assign endpoint_dmaLogic_byteCtx_last = (endpoint_dmaLogic_byteCtx_counter == endpoint_lastAddress);
  assign endpoint_dmaLogic_byteCtx_sel = endpoint_dmaLogic_byteCtx_counter[1:0];
  always @(*) begin
    endpoint_dmaLogic_byteCtx_increment = 1'b0;
    if(endpoint_dmaLogic_fromUsb_run) begin
      if(dataRx_data_valid) begin
        endpoint_dmaLogic_byteCtx_increment = 1'b1;
      end
    end
    if(endpoint_dmaLogic_toUsb_run) begin
      if(endpoint_dmaLogic_storage_readRsp_valid) begin
        if(dataTx_data_ready) begin
          endpoint_dmaLogic_byteCtx_increment = 1'b1;
        end
      end
    end
  end

  always @(*) begin
    endpoint_dmaLogic_toUsb_dmaReady = 1'b0;
    case(endpoint_dmaLogic_stateReg)
      endpoint_dmaLogic_enumDef_INIT : begin
      end
      endpoint_dmaLogic_enumDef_TO_USB : begin
      end
      endpoint_dmaLogic_enumDef_FROM_USB : begin
      end
      endpoint_dmaLogic_enumDef_VALIDATION : begin
      end
      endpoint_dmaLogic_enumDef_CALC_CMD : begin
        if(!endpoint_isIn) begin
          if(endpoint_dataDone) begin
            if(dmaCtx_pendingEmpty) begin
              endpoint_dmaLogic_toUsb_dmaReady = 1'b1;
            end
          end else begin
            if(!when_UsbOhci_l1057) begin
              if(dmaCtx_pendingEmpty) begin
                endpoint_dmaLogic_toUsb_dmaReady = 1'b1;
              end
            end
          end
        end
      end
      endpoint_dmaLogic_enumDef_READ_CMD : begin
      end
      endpoint_dmaLogic_enumDef_WRITE_CMD : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    endpoint_dmaLogic_fromUsb_start = 1'b0;
    case(endpoint_dmaLogic_stateReg)
      endpoint_dmaLogic_enumDef_INIT : begin
        if(endpoint_isIn) begin
          endpoint_dmaLogic_fromUsb_start = 1'b1;
        end
      end
      endpoint_dmaLogic_enumDef_TO_USB : begin
      end
      endpoint_dmaLogic_enumDef_FROM_USB : begin
      end
      endpoint_dmaLogic_enumDef_VALIDATION : begin
      end
      endpoint_dmaLogic_enumDef_CALC_CMD : begin
      end
      endpoint_dmaLogic_enumDef_READ_CMD : begin
      end
      endpoint_dmaLogic_enumDef_WRITE_CMD : begin
      end
      default : begin
      end
    endcase
  end

  assign endpoint_dmaLogic_fromUsb_dmaReady = ((_zz_endpoint_dmaLogic_fromUsb_dmaReady[6 : 4] != 3'b000) || ((! endpoint_dmaLogic_fromUsb_run) && (! endpoint_dmaLogic_fromUsb_push)));
  assign when_UsbOhci_l1011 = (_zz_when_UsbOhci_l1011 < endpoint_dmaLogic_fromUsb_transactionSizeMax);
  assign _zz_5 = ({3'd0,1'b1} <<< endpoint_dmaLogic_byteCtx_sel);
  assign when_UsbOhci_l1020 = (&endpoint_dmaLogic_byteCtx_sel);
  assign endpoint_dmaLogic_headMask = {(endpoint_currentAddress[1 : 0] <= 2'b11),{(endpoint_currentAddress[1 : 0] <= 2'b10),{(endpoint_currentAddress[1 : 0] <= 2'b01),(endpoint_currentAddress[1 : 0] <= 2'b00)}}};
  assign endpoint_dmaLogic_lastMask = {(2'b11 <= _zz_endpoint_dmaLogic_lastMask[1 : 0]),{(2'b10 <= _zz_endpoint_dmaLogic_lastMask_2[1 : 0]),{(2'b01 <= _zz_endpoint_dmaLogic_lastMask_4[1 : 0]),(2'b00 <= _zz_endpoint_dmaLogic_lastMask_6[1 : 0])}}};
  assign endpoint_dmaLogic_fullMask = 4'b1111;
  assign endpoint_dmaLogic_beatLast = (dmaCtx_beatCounter == 4'b1111);
  assign endpoint_dmaLogic_headHit = (_zz_endpoint_dmaLogic_headHit == dmaCtx_beatCounter);
  assign endpoint_dmaLogic_lastHit = (_zz_endpoint_dmaLogic_lastHit == dmaCtx_beatCounter);
  assign endpoint_byteCountCalc = (_zz_endpoint_byteCountCalc + 14'h0001);
  assign endpoint_fsTimeCheck = (endpoint_zeroLength ? (frame_limitCounter == 15'h0) : (_zz_endpoint_fsTimeCheck <= _zz_endpoint_fsTimeCheck_1));
  assign endpoint_timeCheck = ((endpoint_ED_isFs && endpoint_fsTimeCheck) || (endpoint_ED_S && reg_hcLSThreshold_hit));
  assign endpoint_tdUpdateAddress = ((endpoint_TD_retire && (! ((endpoint_isIn && ((endpoint_TD_CC == 4'b0000) || (endpoint_TD_CC == 4'b1001))) && endpoint_dmaLogic_underflow))) ? 32'h0 : endpoint_currentAddressFull);
  always @(*) begin
    operational_wantExit = 1'b0;
    case(operational_stateReg)
      operational_enumDef_SOF : begin
      end
      operational_enumDef_ARBITER : begin
        if(operational_askExit) begin
          operational_wantExit = 1'b1;
        end
      end
      operational_enumDef_END_POINT : begin
      end
      operational_enumDef_PERIODIC_HEAD_CMD : begin
      end
      operational_enumDef_PERIODIC_HEAD_RSP : begin
      end
      operational_enumDef_WAIT_SOF : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    operational_wantStart = 1'b0;
    if(when_StateMachine_l253_7) begin
      operational_wantStart = 1'b1;
    end
  end

  always @(*) begin
    operational_wantKill = 1'b0;
    if(unscheduleAll_fire) begin
      operational_wantKill = 1'b1;
    end
  end

  always @(*) begin
    operational_askExit = 1'b0;
    case(hc_stateReg)
      hc_enumDef_RESET : begin
      end
      hc_enumDef_RESUME : begin
      end
      hc_enumDef_OPERATIONAL : begin
      end
      hc_enumDef_SUSPEND : begin
      end
      hc_enumDef_ANY_TO_RESET : begin
      end
      hc_enumDef_ANY_TO_SUSPEND : begin
        operational_askExit = 1'b1;
      end
      default : begin
      end
    endcase
  end

  assign hc_wantExit = 1'b0;
  always @(*) begin
    hc_wantStart = 1'b0;
    case(hc_stateReg)
      hc_enumDef_RESET : begin
      end
      hc_enumDef_RESUME : begin
      end
      hc_enumDef_OPERATIONAL : begin
      end
      hc_enumDef_SUSPEND : begin
      end
      hc_enumDef_ANY_TO_RESET : begin
      end
      hc_enumDef_ANY_TO_SUSPEND : begin
      end
      default : begin
        hc_wantStart = 1'b1;
      end
    endcase
  end

  assign hc_wantKill = 1'b0;
  always @(*) begin
    reg_hcControl_HCFS = MainState_RESET;
    case(hc_stateReg)
      hc_enumDef_RESET : begin
      end
      hc_enumDef_RESUME : begin
        reg_hcControl_HCFS = MainState_RESUME;
      end
      hc_enumDef_OPERATIONAL : begin
        reg_hcControl_HCFS = MainState_OPERATIONAL;
      end
      hc_enumDef_SUSPEND : begin
        reg_hcControl_HCFS = MainState_SUSPEND;
      end
      hc_enumDef_ANY_TO_RESET : begin
        reg_hcControl_HCFS = MainState_RESET;
      end
      hc_enumDef_ANY_TO_SUSPEND : begin
        reg_hcControl_HCFS = MainState_SUSPEND;
      end
      default : begin
      end
    endcase
  end

  assign io_phy_usbReset = (reg_hcControl_HCFS == MainState_RESET);
  assign io_phy_usbResume = (reg_hcControl_HCFS == MainState_RESUME);
  always @(*) begin
    hc_error = 1'b0;
    case(hc_stateReg)
      hc_enumDef_RESET : begin
        if(reg_hcControl_HCFSWrite_valid) begin
          case(reg_hcControl_HCFSWrite_payload)
            MainState_OPERATIONAL : begin
            end
            default : begin
              hc_error = 1'b1;
            end
          endcase
        end
      end
      hc_enumDef_RESUME : begin
      end
      hc_enumDef_OPERATIONAL : begin
      end
      hc_enumDef_SUSPEND : begin
      end
      hc_enumDef_ANY_TO_RESET : begin
      end
      hc_enumDef_ANY_TO_SUSPEND : begin
      end
      default : begin
      end
    endcase
  end

  assign _zz_reg_hcControl_HCFSWrite_payload = io_ctrl_cmd_payload_fragment_data[7 : 6];
  assign reg_hcControl_HCFSWrite_payload = _zz_reg_hcControl_HCFSWrite_payload;
  assign when_BusSlaveFactory_l1041 = io_ctrl_cmd_payload_fragment_mask[0];
  assign when_BusSlaveFactory_l1041_1 = io_ctrl_cmd_payload_fragment_mask[0];
  assign when_BusSlaveFactory_l1041_2 = io_ctrl_cmd_payload_fragment_mask[0];
  assign when_BusSlaveFactory_l1041_3 = io_ctrl_cmd_payload_fragment_mask[0];
  assign when_BusSlaveFactory_l1041_4 = io_ctrl_cmd_payload_fragment_mask[0];
  assign when_BusSlaveFactory_l1041_5 = io_ctrl_cmd_payload_fragment_mask[1];
  assign when_BusSlaveFactory_l1041_6 = io_ctrl_cmd_payload_fragment_mask[1];
  assign when_BusSlaveFactory_l1041_7 = io_ctrl_cmd_payload_fragment_mask[1];
  assign when_BusSlaveFactory_l1041_8 = io_ctrl_cmd_payload_fragment_mask[1];
  assign when_BusSlaveFactory_l1041_9 = io_ctrl_cmd_payload_fragment_mask[2];
  assign when_BusSlaveFactory_l1041_10 = io_ctrl_cmd_payload_fragment_mask[3];
  assign when_BusSlaveFactory_l1041_11 = io_ctrl_cmd_payload_fragment_mask[0];
  assign when_BusSlaveFactory_l1041_12 = io_ctrl_cmd_payload_fragment_mask[1];
  assign when_BusSlaveFactory_l1041_13 = io_ctrl_cmd_payload_fragment_mask[2];
  assign when_BusSlaveFactory_l1041_14 = io_ctrl_cmd_payload_fragment_mask[3];
  assign when_BusSlaveFactory_l1041_15 = io_ctrl_cmd_payload_fragment_mask[0];
  assign when_BusSlaveFactory_l1041_16 = io_ctrl_cmd_payload_fragment_mask[1];
  assign when_BusSlaveFactory_l1041_17 = io_ctrl_cmd_payload_fragment_mask[2];
  assign when_BusSlaveFactory_l1041_18 = io_ctrl_cmd_payload_fragment_mask[3];
  assign when_BusSlaveFactory_l1041_19 = io_ctrl_cmd_payload_fragment_mask[0];
  assign when_BusSlaveFactory_l1041_20 = io_ctrl_cmd_payload_fragment_mask[1];
  assign when_BusSlaveFactory_l1041_21 = io_ctrl_cmd_payload_fragment_mask[2];
  assign when_BusSlaveFactory_l1041_22 = io_ctrl_cmd_payload_fragment_mask[3];
  assign when_BusSlaveFactory_l1041_23 = io_ctrl_cmd_payload_fragment_mask[0];
  assign when_BusSlaveFactory_l1041_24 = io_ctrl_cmd_payload_fragment_mask[1];
  assign when_BusSlaveFactory_l1041_25 = io_ctrl_cmd_payload_fragment_mask[2];
  assign when_BusSlaveFactory_l1041_26 = io_ctrl_cmd_payload_fragment_mask[3];
  assign when_BusSlaveFactory_l1041_27 = io_ctrl_cmd_payload_fragment_mask[0];
  assign when_BusSlaveFactory_l1041_28 = io_ctrl_cmd_payload_fragment_mask[1];
  assign when_BusSlaveFactory_l1041_29 = io_ctrl_cmd_payload_fragment_mask[2];
  assign when_BusSlaveFactory_l1041_30 = io_ctrl_cmd_payload_fragment_mask[3];
  assign when_BusSlaveFactory_l1041_31 = io_ctrl_cmd_payload_fragment_mask[0];
  assign when_BusSlaveFactory_l1041_32 = io_ctrl_cmd_payload_fragment_mask[1];
  assign when_BusSlaveFactory_l1041_33 = io_ctrl_cmd_payload_fragment_mask[2];
  assign when_BusSlaveFactory_l1041_34 = io_ctrl_cmd_payload_fragment_mask[3];
  assign when_BusSlaveFactory_l1041_35 = io_ctrl_cmd_payload_fragment_mask[3];
  assign when_BusSlaveFactory_l1041_36 = io_ctrl_cmd_payload_fragment_mask[0];
  assign when_BusSlaveFactory_l1041_37 = io_ctrl_cmd_payload_fragment_mask[1];
  assign when_BusSlaveFactory_l1041_38 = io_ctrl_cmd_payload_fragment_mask[0];
  assign when_BusSlaveFactory_l1041_39 = io_ctrl_cmd_payload_fragment_mask[1];
  assign when_BusSlaveFactory_l1041_40 = io_ctrl_cmd_payload_fragment_mask[1];
  assign when_BusSlaveFactory_l1041_41 = io_ctrl_cmd_payload_fragment_mask[1];
  assign when_BusSlaveFactory_l1041_42 = io_ctrl_cmd_payload_fragment_mask[1];
  assign when_BusSlaveFactory_l1041_43 = io_ctrl_cmd_payload_fragment_mask[1];
  assign when_BusSlaveFactory_l1041_44 = io_ctrl_cmd_payload_fragment_mask[3];
  assign when_BusSlaveFactory_l1041_45 = io_ctrl_cmd_payload_fragment_mask[0];
  assign when_BusSlaveFactory_l1041_46 = io_ctrl_cmd_payload_fragment_mask[2];
  assign when_UsbOhci_l241 = (doSoftReset || _zz_when_UsbOhci_l241);
  always @(*) begin
    token_stateNext = token_stateReg;
    case(token_stateReg)
      token_enumDef_INIT : begin
        token_stateNext = token_enumDef_PID;
      end
      token_enumDef_PID : begin
        if(io_phy_tx_ready) begin
          token_stateNext = token_enumDef_B1;
        end
      end
      token_enumDef_B1 : begin
        if(io_phy_tx_ready) begin
          token_stateNext = token_enumDef_B2;
        end
      end
      token_enumDef_B2 : begin
        if(io_phy_tx_ready) begin
          token_stateNext = token_enumDef_EOP;
        end
      end
      token_enumDef_EOP : begin
        if(io_phy_txEop) begin
          token_stateNext = token_enumDef_BOOT;
        end
      end
      default : begin
      end
    endcase
    if(token_wantStart) begin
      token_stateNext = token_enumDef_INIT;
    end
    if(token_wantKill) begin
      token_stateNext = token_enumDef_BOOT;
    end
  end

  assign when_StateMachine_l237 = ((token_stateReg == token_enumDef_BOOT) && (! (token_stateNext == token_enumDef_BOOT)));
  assign unscheduleAll_fire = (unscheduleAll_valid && unscheduleAll_ready);
  always @(*) begin
    dataTx_stateNext = dataTx_stateReg;
    case(dataTx_stateReg)
      dataTx_enumDef_PID : begin
        if(io_phy_tx_ready) begin
          if(dataTx_data_valid) begin
            dataTx_stateNext = dataTx_enumDef_DATA;
          end else begin
            dataTx_stateNext = dataTx_enumDef_CRC_0;
          end
        end
      end
      dataTx_enumDef_DATA : begin
        if(io_phy_tx_ready) begin
          if(dataTx_data_payload_last) begin
            dataTx_stateNext = dataTx_enumDef_CRC_0;
          end
        end
      end
      dataTx_enumDef_CRC_0 : begin
        if(io_phy_tx_ready) begin
          dataTx_stateNext = dataTx_enumDef_CRC_1;
        end
      end
      dataTx_enumDef_CRC_1 : begin
        if(io_phy_tx_ready) begin
          dataTx_stateNext = dataTx_enumDef_EOP;
        end
      end
      dataTx_enumDef_EOP : begin
        if(io_phy_txEop) begin
          dataTx_stateNext = dataTx_enumDef_BOOT;
        end
      end
      default : begin
      end
    endcase
    if(dataTx_wantStart) begin
      dataTx_stateNext = dataTx_enumDef_PID;
    end
    if(dataTx_wantKill) begin
      dataTx_stateNext = dataTx_enumDef_BOOT;
    end
  end

  always @(*) begin
    dataRx_stateNext = dataRx_stateReg;
    case(dataRx_stateReg)
      dataRx_enumDef_IDLE : begin
        if(io_phy_rx_active) begin
          dataRx_stateNext = dataRx_enumDef_PID;
        end else begin
          if(rxTimer_rxTimeout) begin
            dataRx_stateNext = dataRx_enumDef_BOOT;
          end
        end
      end
      dataRx_enumDef_PID : begin
        if(_zz_2) begin
          dataRx_stateNext = dataRx_enumDef_DATA;
        end else begin
          if(when_Misc_l64) begin
            dataRx_stateNext = dataRx_enumDef_BOOT;
          end
        end
      end
      dataRx_enumDef_DATA : begin
        if(when_Misc_l70) begin
          dataRx_stateNext = dataRx_enumDef_BOOT;
        end
      end
      default : begin
      end
    endcase
    if(dataRx_wantStart) begin
      dataRx_stateNext = dataRx_enumDef_IDLE;
    end
    if(dataRx_wantKill) begin
      dataRx_stateNext = dataRx_enumDef_BOOT;
    end
  end

  assign when_Misc_l64 = (! io_phy_rx_active);
  assign when_Misc_l70 = (! io_phy_rx_active);
  assign when_Misc_l71 = ((! (&dataRx_valids)) || (dataRx_crc16_io_result != 16'h800d));
  assign when_Misc_l78 = (&dataRx_valids);
  assign when_StateMachine_l253 = ((! (dataRx_stateReg == dataRx_enumDef_IDLE)) && (dataRx_stateNext == dataRx_enumDef_IDLE));
  assign when_Misc_l85 = (! (dataRx_stateReg == dataRx_enumDef_BOOT));
  always @(*) begin
    sof_stateNext = sof_stateReg;
    case(sof_stateReg)
      sof_enumDef_FRAME_TX : begin
        if(token_wantExit) begin
          sof_stateNext = sof_enumDef_FRAME_NUMBER_CMD;
        end
      end
      sof_enumDef_FRAME_NUMBER_CMD : begin
        if(when_UsbOhci_l614) begin
          sof_stateNext = sof_enumDef_FRAME_NUMBER_RSP;
        end
      end
      sof_enumDef_FRAME_NUMBER_RSP : begin
        if(ioDma_rsp_valid) begin
          sof_stateNext = sof_enumDef_BOOT;
        end
      end
      default : begin
      end
    endcase
    if(sof_wantStart) begin
      sof_stateNext = sof_enumDef_FRAME_TX;
    end
    if(sof_wantKill) begin
      sof_stateNext = sof_enumDef_BOOT;
    end
  end

  assign when_UsbOhci_l207 = (dmaWriteCtx_counter == 4'b0000);
  assign when_UsbOhci_l207_1 = (dmaWriteCtx_counter == 4'b0001);
  assign when_UsbOhci_l614 = (ioDma_cmd_ready && ioDma_cmd_payload_last);
  assign when_StateMachine_l237_1 = ((sof_stateReg == sof_enumDef_BOOT) && (! (sof_stateNext == sof_enumDef_BOOT)));
  always @(*) begin
    endpoint_stateNext = endpoint_stateReg;
    case(endpoint_stateReg)
      endpoint_enumDef_ED_READ_CMD : begin
        if(ioDma_cmd_ready) begin
          endpoint_stateNext = endpoint_enumDef_ED_READ_RSP;
        end
      end
      endpoint_enumDef_ED_READ_RSP : begin
        if(when_UsbOhci_l843) begin
          endpoint_stateNext = endpoint_enumDef_ED_ANALYSE;
        end
      end
      endpoint_enumDef_ED_ANALYSE : begin
        if(when_UsbOhci_l849) begin
          endpoint_stateNext = endpoint_enumDef_BOOT;
        end else begin
          endpoint_stateNext = endpoint_enumDef_TD_READ_CMD;
        end
      end
      endpoint_enumDef_TD_READ_CMD : begin
        if(ioDma_cmd_ready) begin
          endpoint_stateNext = endpoint_enumDef_TD_READ_RSP;
        end
      end
      endpoint_enumDef_TD_READ_RSP : begin
        if(when_UsbOhci_l886) begin
          endpoint_stateNext = endpoint_enumDef_TD_READ_DELAY;
        end
      end
      endpoint_enumDef_TD_READ_DELAY : begin
        endpoint_stateNext = endpoint_enumDef_TD_ANALYSE;
      end
      endpoint_enumDef_TD_ANALYSE : begin
        endpoint_stateNext = endpoint_enumDef_TD_CHECK_TIME;
        if(endpoint_ED_F) begin
          if(endpoint_TD_tooEarlyReg) begin
            endpoint_stateNext = endpoint_enumDef_UPDATE_SYNC;
          end
          if(endpoint_TD_isoOverrunReg) begin
            endpoint_stateNext = endpoint_enumDef_UPDATE_TD_CMD;
          end
        end
      end
      endpoint_enumDef_TD_CHECK_TIME : begin
        if(endpoint_timeCheck) begin
          endpoint_stateNext = endpoint_enumDef_ABORD;
        end else begin
          if(when_UsbOhci_l1173) begin
            endpoint_stateNext = endpoint_enumDef_TOKEN;
          end else begin
            endpoint_stateNext = endpoint_enumDef_BUFFER_READ;
          end
        end
      end
      endpoint_enumDef_BUFFER_READ : begin
        if(endpoint_dmaLogic_toUsb_run) begin
          endpoint_stateNext = endpoint_enumDef_TOKEN;
          if(endpoint_timeCheck) begin
            endpoint_stateNext = endpoint_enumDef_ABORD;
          end
        end
      end
      endpoint_enumDef_TOKEN : begin
        if(token_wantExit) begin
          if(endpoint_isIn) begin
            endpoint_stateNext = endpoint_enumDef_DATA_RX;
          end else begin
            endpoint_stateNext = endpoint_enumDef_DATA_TX;
          end
        end
      end
      endpoint_enumDef_DATA_TX : begin
        if(dataTx_wantExit) begin
          if(endpoint_ED_F) begin
            endpoint_stateNext = endpoint_enumDef_UPDATE_TD_PROCESS;
          end else begin
            endpoint_stateNext = endpoint_enumDef_ACK_RX;
          end
        end
      end
      endpoint_enumDef_DATA_RX : begin
        if(dataRx_wantExit) begin
          endpoint_stateNext = endpoint_enumDef_DATA_RX_VALIDATE;
        end
      end
      endpoint_enumDef_DATA_RX_VALIDATE : begin
        endpoint_stateNext = endpoint_enumDef_DATA_RX_WAIT_DMA;
        if(!dataRx_notResponding) begin
          if(!dataRx_stuffingError) begin
            if(!dataRx_pidError) begin
              if(!endpoint_ED_F) begin
                case(dataRx_pid)
                  4'b1010 : begin
                  end
                  4'b1110 : begin
                  end
                  4'b0011, 4'b1011 : begin
                    if(when_UsbOhci_l1318) begin
                      endpoint_stateNext = endpoint_enumDef_ACK_TX_0;
                    end
                  end
                  default : begin
                  end
                endcase
              end
              if(when_UsbOhci_l1329) begin
                if(!dataRx_crcError) begin
                  if(when_UsbOhci_l1338) begin
                    endpoint_stateNext = endpoint_enumDef_ACK_TX_0;
                  end
                end
              end
            end
          end
        end
      end
      endpoint_enumDef_ACK_RX : begin
        if(when_UsbOhci_l1260) begin
          endpoint_stateNext = endpoint_enumDef_UPDATE_TD_PROCESS;
          if(!when_UsbOhci_l1262) begin
            if(!endpoint_ackRxStuffing) begin
              if(!endpoint_ackRxPidFailure) begin
                case(endpoint_ackRxPid)
                  4'b0010 : begin
                  end
                  4'b1010 : begin
                    endpoint_stateNext = endpoint_enumDef_UPDATE_SYNC;
                  end
                  4'b1110 : begin
                  end
                  default : begin
                  end
                endcase
              end
            end
          end
        end
        if(rxTimer_rxTimeout) begin
          endpoint_stateNext = endpoint_enumDef_UPDATE_TD_PROCESS;
        end
      end
      endpoint_enumDef_ACK_TX_0 : begin
        if(rxTimer_ackTx) begin
          endpoint_stateNext = endpoint_enumDef_ACK_TX_1;
        end
      end
      endpoint_enumDef_ACK_TX_1 : begin
        if(io_phy_tx_ready) begin
          endpoint_stateNext = endpoint_enumDef_ACK_TX_EOP;
        end
      end
      endpoint_enumDef_ACK_TX_EOP : begin
        if(io_phy_txEop) begin
          endpoint_stateNext = endpoint_enumDef_DATA_RX_WAIT_DMA;
        end
      end
      endpoint_enumDef_DATA_RX_WAIT_DMA : begin
        if(when_UsbOhci_l1366) begin
          endpoint_stateNext = endpoint_enumDef_UPDATE_TD_PROCESS;
        end
      end
      endpoint_enumDef_UPDATE_TD_PROCESS : begin
        endpoint_stateNext = endpoint_enumDef_UPDATE_TD_CMD;
        if(!endpoint_ED_F) begin
          if(endpoint_TD_noUpdate) begin
            endpoint_stateNext = endpoint_enumDef_UPDATE_SYNC;
          end
        end
      end
      endpoint_enumDef_UPDATE_TD_CMD : begin
        if(when_UsbOhci_l1448) begin
          endpoint_stateNext = endpoint_enumDef_UPDATE_ED_CMD;
        end
      end
      endpoint_enumDef_UPDATE_ED_CMD : begin
        if(when_UsbOhci_l1463) begin
          endpoint_stateNext = endpoint_enumDef_UPDATE_SYNC;
        end
      end
      endpoint_enumDef_UPDATE_SYNC : begin
        if(dmaCtx_pendingEmpty) begin
          endpoint_stateNext = endpoint_enumDef_BOOT;
        end
      end
      endpoint_enumDef_ABORD : begin
        endpoint_stateNext = endpoint_enumDef_BOOT;
      end
      default : begin
      end
    endcase
    if(endpoint_wantStart) begin
      endpoint_stateNext = endpoint_enumDef_ED_READ_CMD;
    end
    if(endpoint_wantKill) begin
      endpoint_stateNext = endpoint_enumDef_BOOT;
    end
  end

  assign when_UsbOhci_l189 = (ioDma_rsp_valid && (dmaReadCtx_counter == 4'b0000));
  assign when_UsbOhci_l189_1 = (ioDma_rsp_valid && (dmaReadCtx_counter == 4'b0001));
  assign when_UsbOhci_l189_2 = (ioDma_rsp_valid && (dmaReadCtx_counter == 4'b0010));
  assign when_UsbOhci_l189_3 = (ioDma_rsp_valid && (dmaReadCtx_counter == 4'b0011));
  assign when_UsbOhci_l843 = (ioDma_rsp_valid && ioDma_rsp_payload_last);
  assign when_UsbOhci_l849 = ((endpoint_ED_H || endpoint_ED_K) || endpoint_ED_tdEmpty);
  assign when_UsbOhci_l189_4 = (ioDma_rsp_valid && (dmaReadCtx_counter == 4'b0000));
  assign when_UsbOhci_l189_5 = (ioDma_rsp_valid && (dmaReadCtx_counter == 4'b0001));
  assign when_UsbOhci_l189_6 = (ioDma_rsp_valid && (dmaReadCtx_counter == 4'b0010));
  assign when_UsbOhci_l189_7 = (ioDma_rsp_valid && (dmaReadCtx_counter == 4'b0011));
  assign when_UsbOhci_l879 = (endpoint_TD_isoFrameNumber == 3'b000);
  assign when_UsbOhci_l189_8 = (ioDma_rsp_valid && (dmaReadCtx_counter == 4'b0100));
  assign when_UsbOhci_l189_9 = (ioDma_rsp_valid && (dmaReadCtx_counter == 4'b0100));
  assign when_UsbOhci_l879_1 = (endpoint_TD_isoFrameNumber == 3'b001);
  assign when_UsbOhci_l189_10 = (ioDma_rsp_valid && (dmaReadCtx_counter == 4'b0100));
  assign when_UsbOhci_l189_11 = (ioDma_rsp_valid && (dmaReadCtx_counter == 4'b0101));
  assign when_UsbOhci_l879_2 = (endpoint_TD_isoFrameNumber == 3'b010);
  assign when_UsbOhci_l189_12 = (ioDma_rsp_valid && (dmaReadCtx_counter == 4'b0101));
  assign when_UsbOhci_l189_13 = (ioDma_rsp_valid && (dmaReadCtx_counter == 4'b0101));
  assign when_UsbOhci_l879_3 = (endpoint_TD_isoFrameNumber == 3'b011);
  assign when_UsbOhci_l189_14 = (ioDma_rsp_valid && (dmaReadCtx_counter == 4'b0101));
  assign when_UsbOhci_l189_15 = (ioDma_rsp_valid && (dmaReadCtx_counter == 4'b0110));
  assign when_UsbOhci_l879_4 = (endpoint_TD_isoFrameNumber == 3'b100);
  assign when_UsbOhci_l189_16 = (ioDma_rsp_valid && (dmaReadCtx_counter == 4'b0110));
  assign when_UsbOhci_l189_17 = (ioDma_rsp_valid && (dmaReadCtx_counter == 4'b0110));
  assign when_UsbOhci_l879_5 = (endpoint_TD_isoFrameNumber == 3'b101);
  assign when_UsbOhci_l189_18 = (ioDma_rsp_valid && (dmaReadCtx_counter == 4'b0110));
  assign when_UsbOhci_l189_19 = (ioDma_rsp_valid && (dmaReadCtx_counter == 4'b0111));
  assign when_UsbOhci_l879_6 = (endpoint_TD_isoFrameNumber == 3'b110);
  assign when_UsbOhci_l189_20 = (ioDma_rsp_valid && (dmaReadCtx_counter == 4'b0111));
  assign when_UsbOhci_l189_21 = (ioDma_rsp_valid && (dmaReadCtx_counter == 4'b0111));
  assign when_UsbOhci_l879_7 = (endpoint_TD_isoFrameNumber == 3'b111);
  assign when_UsbOhci_l189_22 = (ioDma_rsp_valid && (dmaReadCtx_counter == 4'b0111));
  assign when_UsbOhci_l886 = (ioDma_rsp_fire && ioDma_rsp_payload_last);
  assign _zz_endpoint_lastAddress = (_zz__zz_endpoint_lastAddress - 14'h0001);
  assign when_UsbOhci_l1173 = (endpoint_isIn || endpoint_zeroLength);
  always @(*) begin
    when_UsbOhci_l1329 = 1'b0;
    if(endpoint_ED_F) begin
      case(dataRx_pid)
        4'b1110, 4'b1010 : begin
        end
        4'b0011, 4'b1011 : begin
          when_UsbOhci_l1329 = 1'b1;
        end
        default : begin
        end
      endcase
    end else begin
      case(dataRx_pid)
        4'b1010 : begin
        end
        4'b1110 : begin
        end
        4'b0011, 4'b1011 : begin
          if(!when_UsbOhci_l1318) begin
            when_UsbOhci_l1329 = 1'b1;
          end
        end
        default : begin
        end
      endcase
    end
  end

  assign when_UsbOhci_l1318 = (dataRx_pid == endpoint_TD_dataPidWrong);
  assign when_UsbOhci_l1338 = (! endpoint_ED_F);
  assign when_UsbOhci_l1255 = ((! rxPidOk) || endpoint_ackRxFired);
  assign when_UsbOhci_l1260 = ((! io_phy_rx_active) && endpoint_ackRxActivated);
  assign when_UsbOhci_l1262 = (! endpoint_ackRxFired);
  assign when_UsbOhci_l1386 = ((endpoint_dmaLogic_underflow || (_zz_when_UsbOhci_l1386 < endpoint_currentAddress)) || endpoint_zeroLength);
  assign when_UsbOhci_l1401 = (endpoint_TD_EC != 2'b10);
  assign when_UsbOhci_l207_2 = (dmaWriteCtx_counter == 4'b0000);
  assign when_UsbOhci_l207_3 = (dmaWriteCtx_counter == 4'b0000);
  assign _zz_ioDma_cmd_payload_fragment_data = {endpoint_TD_CC,_zz__zz_ioDma_cmd_payload_fragment_data};
  assign when_UsbOhci_l1433 = (endpoint_TD_isoFrameNumber == 3'b000);
  assign when_UsbOhci_l207_4 = (dmaWriteCtx_counter == 4'b0100);
  assign when_UsbOhci_l1433_1 = (endpoint_TD_isoFrameNumber == 3'b001);
  assign when_UsbOhci_l207_5 = (dmaWriteCtx_counter == 4'b0100);
  assign when_UsbOhci_l1433_2 = (endpoint_TD_isoFrameNumber == 3'b010);
  assign when_UsbOhci_l207_6 = (dmaWriteCtx_counter == 4'b0101);
  assign when_UsbOhci_l1433_3 = (endpoint_TD_isoFrameNumber == 3'b011);
  assign when_UsbOhci_l207_7 = (dmaWriteCtx_counter == 4'b0101);
  assign when_UsbOhci_l1433_4 = (endpoint_TD_isoFrameNumber == 3'b100);
  assign when_UsbOhci_l207_8 = (dmaWriteCtx_counter == 4'b0110);
  assign when_UsbOhci_l1433_5 = (endpoint_TD_isoFrameNumber == 3'b101);
  assign when_UsbOhci_l207_9 = (dmaWriteCtx_counter == 4'b0110);
  assign when_UsbOhci_l1433_6 = (endpoint_TD_isoFrameNumber == 3'b110);
  assign when_UsbOhci_l207_10 = (dmaWriteCtx_counter == 4'b0111);
  assign when_UsbOhci_l1433_7 = (endpoint_TD_isoFrameNumber == 3'b111);
  assign when_UsbOhci_l207_11 = (dmaWriteCtx_counter == 4'b0111);
  assign when_UsbOhci_l207_12 = (dmaWriteCtx_counter == 4'b0000);
  assign when_UsbOhci_l207_13 = (dmaWriteCtx_counter == 4'b0001);
  assign when_UsbOhci_l207_14 = (dmaWriteCtx_counter == 4'b0010);
  assign when_UsbOhci_l1448 = (ioDma_cmd_ready && ioDma_cmd_payload_last);
  assign when_UsbOhci_l207_15 = (dmaWriteCtx_counter == 4'b0010);
  assign when_UsbOhci_l1463 = (ioDma_cmd_ready && ioDma_cmd_payload_last);
  assign when_UsbOhci_l1470 = (! (endpoint_ED_F && endpoint_TD_isoOverrunReg));
  assign when_UsbOhci_l1473 = (endpoint_flowType != FlowType_PERIODIC);
  assign when_StateMachine_l237_2 = ((endpoint_stateReg == endpoint_enumDef_BOOT) && (! (endpoint_stateNext == endpoint_enumDef_BOOT)));
  assign when_StateMachine_l253_1 = ((! (endpoint_stateReg == endpoint_enumDef_TOKEN)) && (endpoint_stateNext == endpoint_enumDef_TOKEN));
  assign when_StateMachine_l253_2 = ((! (endpoint_stateReg == endpoint_enumDef_DATA_TX)) && (endpoint_stateNext == endpoint_enumDef_DATA_TX));
  assign when_StateMachine_l253_3 = ((! (endpoint_stateReg == endpoint_enumDef_DATA_RX)) && (endpoint_stateNext == endpoint_enumDef_DATA_RX));
  assign when_StateMachine_l253_4 = ((! (endpoint_stateReg == endpoint_enumDef_ACK_RX)) && (endpoint_stateNext == endpoint_enumDef_ACK_RX));
  always @(*) begin
    endpoint_dmaLogic_stateNext = endpoint_dmaLogic_stateReg;
    case(endpoint_dmaLogic_stateReg)
      endpoint_dmaLogic_enumDef_INIT : begin
        if(endpoint_isIn) begin
          endpoint_dmaLogic_stateNext = endpoint_dmaLogic_enumDef_CALC_CMD;
        end else begin
          endpoint_dmaLogic_stateNext = endpoint_dmaLogic_enumDef_CALC_CMD;
        end
      end
      endpoint_dmaLogic_enumDef_TO_USB : begin
      end
      endpoint_dmaLogic_enumDef_FROM_USB : begin
      end
      endpoint_dmaLogic_enumDef_VALIDATION : begin
      end
      endpoint_dmaLogic_enumDef_CALC_CMD : begin
        if(endpoint_isIn) begin
          if(when_UsbOhci_l1047) begin
            endpoint_dmaLogic_stateNext = endpoint_dmaLogic_enumDef_BOOT;
          end else begin
            if(endpoint_dmaLogic_fromUsb_dmaReady) begin
              endpoint_dmaLogic_stateNext = endpoint_dmaLogic_enumDef_WRITE_CMD;
            end
          end
        end else begin
          if(!endpoint_dataDone) begin
            if(when_UsbOhci_l1057) begin
              endpoint_dmaLogic_stateNext = endpoint_dmaLogic_enumDef_READ_CMD;
            end
          end
        end
      end
      endpoint_dmaLogic_enumDef_READ_CMD : begin
        if(ioDma_cmd_ready) begin
          endpoint_dmaLogic_stateNext = endpoint_dmaLogic_enumDef_CALC_CMD;
        end
      end
      endpoint_dmaLogic_enumDef_WRITE_CMD : begin
        if(ioDma_cmd_ready) begin
          if(endpoint_dmaLogic_beatLast) begin
            endpoint_dmaLogic_stateNext = endpoint_dmaLogic_enumDef_CALC_CMD;
          end
        end
      end
      default : begin
      end
    endcase
    if(endpoint_dmaLogic_toUsb_run) begin
      if(endpoint_dmaLogic_storage_readRsp_valid) begin
        if(dataTx_data_ready) begin
          if(endpoint_dmaLogic_byteCtx_last) begin
            endpoint_dmaLogic_stateNext = endpoint_dmaLogic_enumDef_BOOT;
          end
        end
      end
    end
    if(endpoint_dmaLogic_wantStart) begin
      endpoint_dmaLogic_stateNext = endpoint_dmaLogic_enumDef_INIT;
    end
    if(endpoint_dmaLogic_wantKill) begin
      endpoint_dmaLogic_stateNext = endpoint_dmaLogic_enumDef_BOOT;
    end
  end

  assign when_UsbOhci_l1047 = ((! endpoint_dmaLogic_fromUsb_run) && (endpoint_dataDone || (endpoint_dmaLogic_fromUsbCounter == 11'h0)));
  assign when_UsbOhci_l1057 = (! endpoint_dmaLogic_storage_full);
  assign when_UsbOhci_l1093 = (! endpoint_dmaLogic_storageReadDone);
  assign when_UsbOhci_l1098 = (&endpoint_dmaLogic_storage_readPtr[3 : 0]);
  assign when_StateMachine_l253_5 = ((! (endpoint_dmaLogic_stateReg == endpoint_dmaLogic_enumDef_WRITE_CMD)) && (endpoint_dmaLogic_stateNext == endpoint_dmaLogic_enumDef_WRITE_CMD));
  assign when_UsbOhci_l973 = (&endpoint_dmaLogic_byteCtx_sel);
  assign when_UsbOhci_l958 = ((endpoint_dmaLogic_stateNext == endpoint_dmaLogic_enumDef_BOOT) && (endpoint_dmaLogic_stateReg != endpoint_dmaLogic_enumDef_BOOT));
  assign when_UsbOhci_l997 = ((endpoint_dmaLogic_stateNext == endpoint_dmaLogic_enumDef_BOOT) && (endpoint_dmaLogic_stateReg != endpoint_dmaLogic_enumDef_BOOT));
  assign endpoint_dmaLogic_fsmStopped = (endpoint_dmaLogic_stateReg == endpoint_dmaLogic_enumDef_BOOT);
  assign when_UsbOhci_l1366 = (endpoint_dmaLogic_stateReg == endpoint_dmaLogic_enumDef_BOOT);
  always @(*) begin
    operational_stateNext = operational_stateReg;
    case(operational_stateReg)
      operational_enumDef_SOF : begin
        if(sof_wantExit) begin
          operational_stateNext = operational_enumDef_ARBITER;
        end
      end
      operational_enumDef_ARBITER : begin
        if(operational_askExit) begin
          operational_stateNext = operational_enumDef_BOOT;
        end else begin
          if(frame_limitHit) begin
            operational_stateNext = operational_enumDef_WAIT_SOF;
          end else begin
            if(when_UsbOhci_l1542) begin
              if(when_UsbOhci_l1543) begin
                operational_stateNext = operational_enumDef_PERIODIC_HEAD_CMD;
              end else begin
                if(!reg_hcPeriodCurrentED_isZero) begin
                  operational_stateNext = operational_enumDef_END_POINT;
                end
              end
            end else begin
              if(priority_bulk) begin
                if(operational_allowBulk) begin
                  if(!reg_hcBulkCurrentED_isZero) begin
                    operational_stateNext = operational_enumDef_END_POINT;
                  end
                end
              end else begin
                if(operational_allowControl) begin
                  if(!reg_hcControlCurrentED_isZero) begin
                    operational_stateNext = operational_enumDef_END_POINT;
                  end
                end
              end
            end
          end
        end
      end
      operational_enumDef_END_POINT : begin
        if(endpoint_wantExit) begin
          case(endpoint_status_1)
            endpoint_Status_OK : begin
              operational_stateNext = operational_enumDef_ARBITER;
            end
            default : begin
              operational_stateNext = operational_enumDef_WAIT_SOF;
            end
          endcase
        end
      end
      operational_enumDef_PERIODIC_HEAD_CMD : begin
        if(ioDma_cmd_ready) begin
          operational_stateNext = operational_enumDef_PERIODIC_HEAD_RSP;
        end
      end
      operational_enumDef_PERIODIC_HEAD_RSP : begin
        if(ioDma_rsp_valid) begin
          operational_stateNext = operational_enumDef_ARBITER;
        end
      end
      operational_enumDef_WAIT_SOF : begin
        if(frame_tick) begin
          operational_stateNext = operational_enumDef_SOF;
        end
      end
      default : begin
      end
    endcase
    if(operational_wantStart) begin
      operational_stateNext = operational_enumDef_WAIT_SOF;
    end
    if(operational_wantKill) begin
      operational_stateNext = operational_enumDef_BOOT;
    end
  end

  assign when_UsbOhci_l1516 = (operational_allowPeriodic && (! operational_periodicDone));
  assign when_UsbOhci_l1543 = (! operational_periodicHeadFetched);
  assign when_UsbOhci_l1542 = ((operational_allowPeriodic && (! operational_periodicDone)) && (! frame_section1));
  assign when_StateMachine_l237_3 = ((operational_stateReg == operational_enumDef_BOOT) && (! (operational_stateNext == operational_enumDef_BOOT)));
  assign when_StateMachine_l253_6 = ((! (operational_stateReg == operational_enumDef_SOF)) && (operational_stateNext == operational_enumDef_SOF));
  assign hc_operationalIsDone = (operational_stateReg == operational_enumDef_BOOT);
  always @(*) begin
    hc_stateNext = hc_stateReg;
    case(hc_stateReg)
      hc_enumDef_RESET : begin
        if(reg_hcControl_HCFSWrite_valid) begin
          case(reg_hcControl_HCFSWrite_payload)
            MainState_OPERATIONAL : begin
              hc_stateNext = hc_enumDef_OPERATIONAL;
            end
            default : begin
            end
          endcase
        end
      end
      hc_enumDef_RESUME : begin
        if(when_UsbOhci_l1671) begin
          hc_stateNext = hc_enumDef_OPERATIONAL;
        end
      end
      hc_enumDef_OPERATIONAL : begin
      end
      hc_enumDef_SUSPEND : begin
        if(when_UsbOhci_l1680) begin
          hc_stateNext = hc_enumDef_RESUME;
        end else begin
          if(when_UsbOhci_l1683) begin
            hc_stateNext = hc_enumDef_OPERATIONAL;
          end
        end
      end
      hc_enumDef_ANY_TO_RESET : begin
        if(when_UsbOhci_l1694) begin
          hc_stateNext = hc_enumDef_RESET;
        end
      end
      hc_enumDef_ANY_TO_SUSPEND : begin
        if(when_UsbOhci_l1707) begin
          hc_stateNext = hc_enumDef_SUSPEND;
        end
      end
      default : begin
      end
    endcase
    if(when_UsbOhci_l1714) begin
      hc_stateNext = hc_enumDef_ANY_TO_RESET;
    end
    if(reg_hcCommandStatus_startSoftReset) begin
      hc_stateNext = hc_enumDef_ANY_TO_SUSPEND;
    end
    if(hc_wantStart) begin
      hc_stateNext = hc_enumDef_RESET;
    end
    if(hc_wantKill) begin
      hc_stateNext = hc_enumDef_BOOT;
    end
  end

  assign when_UsbOhci_l1671 = (reg_hcControl_HCFSWrite_valid && (reg_hcControl_HCFSWrite_payload == MainState_OPERATIONAL));
  assign when_UsbOhci_l1680 = (reg_hcRhStatus_DRWE && (|{reg_hcRhPortStatus_1_CSC_reg,reg_hcRhPortStatus_0_CSC_reg}));
  assign when_UsbOhci_l1683 = (reg_hcControl_HCFSWrite_valid && (reg_hcControl_HCFSWrite_payload == MainState_OPERATIONAL));
  assign when_UsbOhci_l1694 = (! doUnschedule);
  assign when_UsbOhci_l1707 = (((! doUnschedule) && (! doSoftReset)) && hc_operationalIsDone);
  assign when_StateMachine_l253_7 = ((! (hc_stateReg == hc_enumDef_OPERATIONAL)) && (hc_stateNext == hc_enumDef_OPERATIONAL));
  assign when_StateMachine_l253_8 = ((! (hc_stateReg == hc_enumDef_ANY_TO_RESET)) && (hc_stateNext == hc_enumDef_ANY_TO_RESET));
  assign when_StateMachine_l253_9 = ((! (hc_stateReg == hc_enumDef_ANY_TO_SUSPEND)) && (hc_stateNext == hc_enumDef_ANY_TO_SUSPEND));
  assign when_UsbOhci_l1714 = (reg_hcControl_HCFSWrite_valid && (reg_hcControl_HCFSWrite_payload == MainState_RESET));
  always @(posedge clk_peripheral or posedge reset_peripheral) begin
    if(reset_peripheral) begin
      dmaCtx_pendingCounter <= 4'b0000;
      dmaCtx_beatCounter <= 4'b0000;
      io_dma_cmd_payload_first <= 1'b1;
      dmaReadCtx_counter <= 4'b0000;
      dmaWriteCtx_counter <= 4'b0000;
      _zz_io_ctrl_rsp_valid_1 <= 1'b0;
      doUnschedule <= 1'b0;
      doSoftReset <= 1'b0;
      reg_hcControl_IR <= 1'b0;
      reg_hcControl_RWC <= 1'b0;
      reg_hcFmNumber_overflow <= 1'b0;
      reg_hcPeriodicStart_PS <= 14'h0;
      io_phy_overcurrent_regNext <= 1'b0;
      reg_hcRhPortStatus_0_connected <= 1'b0;
      reg_hcRhPortStatus_0_CCS_regNext <= 1'b0;
      reg_hcRhPortStatus_1_connected <= 1'b0;
      reg_hcRhPortStatus_1_CCS_regNext <= 1'b0;
      interruptDelay_counter <= 3'b111;
      _zz_endpoint_dmaLogic_storage_readRsp_valid <= 1'b0;
      endpoint_dmaLogic_toUsb_run <= 1'b0;
      endpoint_dmaLogic_fromUsb_push <= 1'b0;
      endpoint_dmaLogic_fromUsb_run <= 1'b0;
      endpoint_dmaLogic_inBurst <= 1'b0;
      _zz_when_UsbOhci_l241 <= 1'b1;
      token_stateReg <= token_enumDef_BOOT;
      dataTx_stateReg <= dataTx_enumDef_BOOT;
      dataRx_stateReg <= dataRx_enumDef_BOOT;
      sof_stateReg <= sof_enumDef_BOOT;
      endpoint_stateReg <= endpoint_enumDef_BOOT;
      endpoint_dmaLogic_stateReg <= endpoint_dmaLogic_enumDef_BOOT;
      operational_stateReg <= operational_enumDef_BOOT;
      hc_stateReg <= hc_enumDef_BOOT;
    end else begin
      dmaCtx_pendingCounter <= (_zz_dmaCtx_pendingCounter - _zz_dmaCtx_pendingCounter_3);
      if(ioDma_cmd_fire) begin
        dmaCtx_beatCounter <= (dmaCtx_beatCounter + 4'b0001);
        if(io_dma_cmd_payload_last) begin
          dmaCtx_beatCounter <= 4'b0000;
        end
      end
      if(io_dma_cmd_fire) begin
        io_dma_cmd_payload_first <= io_dma_cmd_payload_last;
      end
      if(ioDma_rsp_fire) begin
        dmaReadCtx_counter <= (dmaReadCtx_counter + 4'b0001);
        if(ioDma_rsp_payload_last) begin
          dmaReadCtx_counter <= 4'b0000;
        end
      end
      if(ioDma_cmd_fire) begin
        dmaWriteCtx_counter <= (dmaWriteCtx_counter + 4'b0001);
        if(ioDma_cmd_payload_last) begin
          dmaWriteCtx_counter <= 4'b0000;
        end
      end
      if(_zz_ctrl_rsp_ready_1) begin
        _zz_io_ctrl_rsp_valid_1 <= (ctrl_rsp_valid && _zz_ctrl_rsp_ready);
      end
      if(unscheduleAll_ready) begin
        doUnschedule <= 1'b0;
      end
      if(when_UsbOhci_l224) begin
        doSoftReset <= 1'b0;
      end
      io_phy_overcurrent_regNext <= io_phy_overcurrent;
      if(io_phy_ports_0_connect) begin
        reg_hcRhPortStatus_0_connected <= 1'b1;
      end
      if(io_phy_ports_0_disconnect) begin
        reg_hcRhPortStatus_0_connected <= 1'b0;
      end
      reg_hcRhPortStatus_0_CCS_regNext <= reg_hcRhPortStatus_0_CCS;
      if(io_phy_ports_1_connect) begin
        reg_hcRhPortStatus_1_connected <= 1'b1;
      end
      if(io_phy_ports_1_disconnect) begin
        reg_hcRhPortStatus_1_connected <= 1'b0;
      end
      reg_hcRhPortStatus_1_CCS_regNext <= reg_hcRhPortStatus_1_CCS;
      if(frame_reload) begin
        if(when_UsbOhci_l528) begin
          reg_hcFmNumber_overflow <= 1'b1;
        end
      end
      if(when_UsbOhci_l673) begin
        interruptDelay_counter <= (interruptDelay_counter - 3'b001);
      end
      if(when_UsbOhci_l677) begin
        interruptDelay_counter <= interruptDelay_load_payload;
      end
      if(interruptDelay_disable) begin
        interruptDelay_counter <= 3'b111;
      end
      if(endpoint_dmaLogic_storage_readRsp_ready) begin
        _zz_endpoint_dmaLogic_storage_readRsp_valid <= 1'b0;
      end
      if(endpoint_dmaLogic_storage_readCmd_ready) begin
        _zz_endpoint_dmaLogic_storage_readRsp_valid <= endpoint_dmaLogic_storage_readCmd_valid;
      end
      if(endpoint_dmaLogic_toUsb_dmaReady) begin
        endpoint_dmaLogic_toUsb_run <= 1'b1;
      end
      if(when_UsbOhci_l958) begin
        endpoint_dmaLogic_toUsb_run <= 1'b0;
      end
      endpoint_dmaLogic_fromUsb_push <= 1'b0;
      if(endpoint_dmaLogic_fromUsb_start) begin
        endpoint_dmaLogic_fromUsb_run <= 1'b1;
      end
      if(when_UsbOhci_l997) begin
        endpoint_dmaLogic_fromUsb_run <= 1'b0;
      end
      if(endpoint_dmaLogic_fromUsb_run) begin
        if(dataRx_wantExit) begin
          endpoint_dmaLogic_fromUsb_push <= (|endpoint_dmaLogic_byteCtx_sel);
          endpoint_dmaLogic_fromUsb_run <= 1'b0;
        end
        if(dataRx_data_valid) begin
          if(when_UsbOhci_l1020) begin
            endpoint_dmaLogic_fromUsb_push <= 1'b1;
          end
        end
      end
      case(io_ctrl_cmd_payload_fragment_address)
        12'h004 : begin
          if(ctrl_doWrite) begin
            if(when_BusSlaveFactory_l1041_5) begin
              reg_hcControl_IR <= io_ctrl_cmd_payload_fragment_data[8];
            end
            if(when_BusSlaveFactory_l1041_6) begin
              reg_hcControl_RWC <= io_ctrl_cmd_payload_fragment_data[9];
            end
          end
        end
        12'h040 : begin
          if(ctrl_doWrite) begin
            if(when_BusSlaveFactory_l1041_36) begin
              reg_hcPeriodicStart_PS[7 : 0] <= io_ctrl_cmd_payload_fragment_data[7 : 0];
            end
            if(when_BusSlaveFactory_l1041_37) begin
              reg_hcPeriodicStart_PS[13 : 8] <= io_ctrl_cmd_payload_fragment_data[13 : 8];
            end
          end
        end
        default : begin
        end
      endcase
      _zz_when_UsbOhci_l241 <= 1'b0;
      token_stateReg <= token_stateNext;
      dataTx_stateReg <= dataTx_stateNext;
      dataRx_stateReg <= dataRx_stateNext;
      sof_stateReg <= sof_stateNext;
      case(sof_stateReg)
        sof_enumDef_FRAME_TX : begin
        end
        sof_enumDef_FRAME_NUMBER_CMD : begin
        end
        sof_enumDef_FRAME_NUMBER_RSP : begin
          if(ioDma_rsp_valid) begin
            reg_hcFmNumber_overflow <= 1'b0;
          end
        end
        default : begin
        end
      endcase
      endpoint_stateReg <= endpoint_stateNext;
      endpoint_dmaLogic_stateReg <= endpoint_dmaLogic_stateNext;
      case(endpoint_dmaLogic_stateReg)
        endpoint_dmaLogic_enumDef_INIT : begin
        end
        endpoint_dmaLogic_enumDef_TO_USB : begin
        end
        endpoint_dmaLogic_enumDef_FROM_USB : begin
        end
        endpoint_dmaLogic_enumDef_VALIDATION : begin
        end
        endpoint_dmaLogic_enumDef_CALC_CMD : begin
        end
        endpoint_dmaLogic_enumDef_READ_CMD : begin
        end
        endpoint_dmaLogic_enumDef_WRITE_CMD : begin
          if(ioDma_cmd_ready) begin
            if(endpoint_dmaLogic_headHit) begin
              endpoint_dmaLogic_inBurst <= 1'b1;
            end
            if(endpoint_dmaLogic_lastHit) begin
              endpoint_dmaLogic_inBurst <= 1'b0;
            end
          end
        end
        default : begin
        end
      endcase
      if(when_StateMachine_l253_5) begin
        endpoint_dmaLogic_inBurst <= 1'b0;
      end
      operational_stateReg <= operational_stateNext;
      hc_stateReg <= hc_stateNext;
      if(when_StateMachine_l253_8) begin
        doUnschedule <= 1'b1;
      end
      if(when_StateMachine_l253_9) begin
        doUnschedule <= 1'b1;
      end
      if(reg_hcCommandStatus_startSoftReset) begin
        doSoftReset <= 1'b1;
      end
    end
  end

  always @(posedge clk_peripheral) begin
    if(_zz_ctrl_rsp_ready_1) begin
      _zz_io_ctrl_rsp_payload_last <= ctrl_rsp_payload_last;
      _zz_io_ctrl_rsp_payload_fragment_opcode <= ctrl_rsp_payload_fragment_opcode;
      _zz_io_ctrl_rsp_payload_fragment_data <= ctrl_rsp_payload_fragment_data;
    end
    if(when_BusSlaveFactory_l377_1) begin
      if(when_BusSlaveFactory_l379_1) begin
        reg_hcCommandStatus_CLF <= _zz_reg_hcCommandStatus_CLF[0];
      end
    end
    if(when_BusSlaveFactory_l377_2) begin
      if(when_BusSlaveFactory_l379_2) begin
        reg_hcCommandStatus_BLF <= _zz_reg_hcCommandStatus_BLF[0];
      end
    end
    if(when_BusSlaveFactory_l377_3) begin
      if(when_BusSlaveFactory_l379_3) begin
        reg_hcCommandStatus_OCR <= _zz_reg_hcCommandStatus_OCR[0];
      end
    end
    if(when_BusSlaveFactory_l377_4) begin
      if(when_BusSlaveFactory_l379_4) begin
        reg_hcInterrupt_MIE <= _zz_reg_hcInterrupt_MIE[0];
      end
    end
    if(when_BusSlaveFactory_l341) begin
      if(when_BusSlaveFactory_l347) begin
        reg_hcInterrupt_MIE <= _zz_reg_hcInterrupt_MIE_1[0];
      end
    end
    if(when_BusSlaveFactory_l341_1) begin
      if(when_BusSlaveFactory_l347_1) begin
        reg_hcInterrupt_SO_status <= _zz_reg_hcInterrupt_SO_status[0];
      end
    end
    if(when_BusSlaveFactory_l377_5) begin
      if(when_BusSlaveFactory_l379_5) begin
        reg_hcInterrupt_SO_enable <= _zz_reg_hcInterrupt_SO_enable[0];
      end
    end
    if(when_BusSlaveFactory_l341_2) begin
      if(when_BusSlaveFactory_l347_2) begin
        reg_hcInterrupt_SO_enable <= _zz_reg_hcInterrupt_SO_enable_1[0];
      end
    end
    if(when_BusSlaveFactory_l341_3) begin
      if(when_BusSlaveFactory_l347_3) begin
        reg_hcInterrupt_WDH_status <= _zz_reg_hcInterrupt_WDH_status[0];
      end
    end
    if(when_BusSlaveFactory_l377_6) begin
      if(when_BusSlaveFactory_l379_6) begin
        reg_hcInterrupt_WDH_enable <= _zz_reg_hcInterrupt_WDH_enable[0];
      end
    end
    if(when_BusSlaveFactory_l341_4) begin
      if(when_BusSlaveFactory_l347_4) begin
        reg_hcInterrupt_WDH_enable <= _zz_reg_hcInterrupt_WDH_enable_1[0];
      end
    end
    if(when_BusSlaveFactory_l341_5) begin
      if(when_BusSlaveFactory_l347_5) begin
        reg_hcInterrupt_SF_status <= _zz_reg_hcInterrupt_SF_status[0];
      end
    end
    if(when_BusSlaveFactory_l377_7) begin
      if(when_BusSlaveFactory_l379_7) begin
        reg_hcInterrupt_SF_enable <= _zz_reg_hcInterrupt_SF_enable[0];
      end
    end
    if(when_BusSlaveFactory_l341_6) begin
      if(when_BusSlaveFactory_l347_6) begin
        reg_hcInterrupt_SF_enable <= _zz_reg_hcInterrupt_SF_enable_1[0];
      end
    end
    if(when_BusSlaveFactory_l341_7) begin
      if(when_BusSlaveFactory_l347_7) begin
        reg_hcInterrupt_RD_status <= _zz_reg_hcInterrupt_RD_status[0];
      end
    end
    if(when_BusSlaveFactory_l377_8) begin
      if(when_BusSlaveFactory_l379_8) begin
        reg_hcInterrupt_RD_enable <= _zz_reg_hcInterrupt_RD_enable[0];
      end
    end
    if(when_BusSlaveFactory_l341_8) begin
      if(when_BusSlaveFactory_l347_8) begin
        reg_hcInterrupt_RD_enable <= _zz_reg_hcInterrupt_RD_enable_1[0];
      end
    end
    if(when_BusSlaveFactory_l341_9) begin
      if(when_BusSlaveFactory_l347_9) begin
        reg_hcInterrupt_UE_status <= _zz_reg_hcInterrupt_UE_status[0];
      end
    end
    if(when_BusSlaveFactory_l377_9) begin
      if(when_BusSlaveFactory_l379_9) begin
        reg_hcInterrupt_UE_enable <= _zz_reg_hcInterrupt_UE_enable[0];
      end
    end
    if(when_BusSlaveFactory_l341_10) begin
      if(when_BusSlaveFactory_l347_10) begin
        reg_hcInterrupt_UE_enable <= _zz_reg_hcInterrupt_UE_enable_1[0];
      end
    end
    if(when_BusSlaveFactory_l341_11) begin
      if(when_BusSlaveFactory_l347_11) begin
        reg_hcInterrupt_FNO_status <= _zz_reg_hcInterrupt_FNO_status[0];
      end
    end
    if(when_BusSlaveFactory_l377_10) begin
      if(when_BusSlaveFactory_l379_10) begin
        reg_hcInterrupt_FNO_enable <= _zz_reg_hcInterrupt_FNO_enable[0];
      end
    end
    if(when_BusSlaveFactory_l341_12) begin
      if(when_BusSlaveFactory_l347_12) begin
        reg_hcInterrupt_FNO_enable <= _zz_reg_hcInterrupt_FNO_enable_1[0];
      end
    end
    if(when_BusSlaveFactory_l341_13) begin
      if(when_BusSlaveFactory_l347_13) begin
        reg_hcInterrupt_RHSC_status <= _zz_reg_hcInterrupt_RHSC_status[0];
      end
    end
    if(when_BusSlaveFactory_l377_11) begin
      if(when_BusSlaveFactory_l379_11) begin
        reg_hcInterrupt_RHSC_enable <= _zz_reg_hcInterrupt_RHSC_enable[0];
      end
    end
    if(when_BusSlaveFactory_l341_14) begin
      if(when_BusSlaveFactory_l347_14) begin
        reg_hcInterrupt_RHSC_enable <= _zz_reg_hcInterrupt_RHSC_enable_1[0];
      end
    end
    if(when_BusSlaveFactory_l341_15) begin
      if(when_BusSlaveFactory_l347_15) begin
        reg_hcInterrupt_OC_status <= _zz_reg_hcInterrupt_OC_status[0];
      end
    end
    if(when_BusSlaveFactory_l377_12) begin
      if(when_BusSlaveFactory_l379_12) begin
        reg_hcInterrupt_OC_enable <= _zz_reg_hcInterrupt_OC_enable[0];
      end
    end
    if(when_BusSlaveFactory_l341_16) begin
      if(when_BusSlaveFactory_l347_16) begin
        reg_hcInterrupt_OC_enable <= _zz_reg_hcInterrupt_OC_enable_1[0];
      end
    end
    if(reg_hcCommandStatus_OCR) begin
      reg_hcInterrupt_OC_status <= 1'b1;
    end
    if(when_BusSlaveFactory_l341_17) begin
      if(when_BusSlaveFactory_l347_17) begin
        reg_hcRhStatus_CCIC <= _zz_reg_hcRhStatus_CCIC[0];
      end
    end
    if(when_UsbOhci_l397) begin
      reg_hcRhStatus_CCIC <= 1'b1;
    end
    if(reg_hcRhStatus_setRemoteWakeupEnable) begin
      reg_hcRhStatus_DRWE <= 1'b1;
    end
    if(reg_hcRhStatus_clearRemoteWakeupEnable) begin
      reg_hcRhStatus_DRWE <= 1'b0;
    end
    if(reg_hcRhPortStatus_0_CSC_clear) begin
      reg_hcRhPortStatus_0_CSC_reg <= 1'b0;
    end
    if(reg_hcRhPortStatus_0_CSC_set) begin
      reg_hcRhPortStatus_0_CSC_reg <= 1'b1;
    end
    if(reg_hcRhPortStatus_0_CSC_set) begin
      reg_hcInterrupt_RHSC_status <= 1'b1;
    end
    if(reg_hcRhPortStatus_0_PESC_clear) begin
      reg_hcRhPortStatus_0_PESC_reg <= 1'b0;
    end
    if(reg_hcRhPortStatus_0_PESC_set) begin
      reg_hcRhPortStatus_0_PESC_reg <= 1'b1;
    end
    if(reg_hcRhPortStatus_0_PESC_set) begin
      reg_hcInterrupt_RHSC_status <= 1'b1;
    end
    if(reg_hcRhPortStatus_0_PSSC_clear) begin
      reg_hcRhPortStatus_0_PSSC_reg <= 1'b0;
    end
    if(reg_hcRhPortStatus_0_PSSC_set) begin
      reg_hcRhPortStatus_0_PSSC_reg <= 1'b1;
    end
    if(reg_hcRhPortStatus_0_PSSC_set) begin
      reg_hcInterrupt_RHSC_status <= 1'b1;
    end
    if(reg_hcRhPortStatus_0_OCIC_clear) begin
      reg_hcRhPortStatus_0_OCIC_reg <= 1'b0;
    end
    if(reg_hcRhPortStatus_0_OCIC_set) begin
      reg_hcRhPortStatus_0_OCIC_reg <= 1'b1;
    end
    if(reg_hcRhPortStatus_0_OCIC_set) begin
      reg_hcInterrupt_RHSC_status <= 1'b1;
    end
    if(reg_hcRhPortStatus_0_PRSC_clear) begin
      reg_hcRhPortStatus_0_PRSC_reg <= 1'b0;
    end
    if(reg_hcRhPortStatus_0_PRSC_set) begin
      reg_hcRhPortStatus_0_PRSC_reg <= 1'b1;
    end
    if(reg_hcRhPortStatus_0_PRSC_set) begin
      reg_hcInterrupt_RHSC_status <= 1'b1;
    end
    if(when_UsbOhci_l448) begin
      reg_hcRhPortStatus_0_PES <= 1'b0;
    end
    if(when_UsbOhci_l448_1) begin
      reg_hcRhPortStatus_0_PES <= 1'b1;
    end
    if(when_UsbOhci_l448_2) begin
      reg_hcRhPortStatus_0_PES <= 1'b1;
    end
    if(when_UsbOhci_l449) begin
      reg_hcRhPortStatus_0_PSS <= 1'b0;
    end
    if(when_UsbOhci_l449_1) begin
      reg_hcRhPortStatus_0_PSS <= 1'b1;
    end
    if(when_UsbOhci_l450) begin
      reg_hcRhPortStatus_0_suspend <= 1'b1;
    end
    if(when_UsbOhci_l451) begin
      reg_hcRhPortStatus_0_resume <= 1'b1;
    end
    if(when_UsbOhci_l452) begin
      reg_hcRhPortStatus_0_reset <= 1'b1;
    end
    if(reg_hcRhDescriptorA_NPS) begin
      reg_hcRhPortStatus_0_PPS <= 1'b1;
    end else begin
      if(reg_hcRhDescriptorA_PSM) begin
        if(when_UsbOhci_l458) begin
          if(reg_hcRhPortStatus_0_clearPortPower) begin
            reg_hcRhPortStatus_0_PPS <= 1'b0;
          end
          if(reg_hcRhPortStatus_0_setPortPower) begin
            reg_hcRhPortStatus_0_PPS <= 1'b1;
          end
        end else begin
          if(reg_hcRhStatus_clearGlobalPower) begin
            reg_hcRhPortStatus_0_PPS <= 1'b0;
          end
          if(reg_hcRhStatus_setGlobalPower) begin
            reg_hcRhPortStatus_0_PPS <= 1'b1;
          end
        end
      end else begin
        if(reg_hcRhStatus_clearGlobalPower) begin
          reg_hcRhPortStatus_0_PPS <= 1'b0;
        end
        if(reg_hcRhStatus_setGlobalPower) begin
          reg_hcRhPortStatus_0_PPS <= 1'b1;
        end
      end
    end
    if(io_phy_ports_0_resume_fire) begin
      reg_hcRhPortStatus_0_resume <= 1'b0;
    end
    if(io_phy_ports_0_reset_fire) begin
      reg_hcRhPortStatus_0_reset <= 1'b0;
    end
    if(io_phy_ports_0_suspend_fire) begin
      reg_hcRhPortStatus_0_suspend <= 1'b0;
    end
    if(reg_hcRhPortStatus_1_CSC_clear) begin
      reg_hcRhPortStatus_1_CSC_reg <= 1'b0;
    end
    if(reg_hcRhPortStatus_1_CSC_set) begin
      reg_hcRhPortStatus_1_CSC_reg <= 1'b1;
    end
    if(reg_hcRhPortStatus_1_CSC_set) begin
      reg_hcInterrupt_RHSC_status <= 1'b1;
    end
    if(reg_hcRhPortStatus_1_PESC_clear) begin
      reg_hcRhPortStatus_1_PESC_reg <= 1'b0;
    end
    if(reg_hcRhPortStatus_1_PESC_set) begin
      reg_hcRhPortStatus_1_PESC_reg <= 1'b1;
    end
    if(reg_hcRhPortStatus_1_PESC_set) begin
      reg_hcInterrupt_RHSC_status <= 1'b1;
    end
    if(reg_hcRhPortStatus_1_PSSC_clear) begin
      reg_hcRhPortStatus_1_PSSC_reg <= 1'b0;
    end
    if(reg_hcRhPortStatus_1_PSSC_set) begin
      reg_hcRhPortStatus_1_PSSC_reg <= 1'b1;
    end
    if(reg_hcRhPortStatus_1_PSSC_set) begin
      reg_hcInterrupt_RHSC_status <= 1'b1;
    end
    if(reg_hcRhPortStatus_1_OCIC_clear) begin
      reg_hcRhPortStatus_1_OCIC_reg <= 1'b0;
    end
    if(reg_hcRhPortStatus_1_OCIC_set) begin
      reg_hcRhPortStatus_1_OCIC_reg <= 1'b1;
    end
    if(reg_hcRhPortStatus_1_OCIC_set) begin
      reg_hcInterrupt_RHSC_status <= 1'b1;
    end
    if(reg_hcRhPortStatus_1_PRSC_clear) begin
      reg_hcRhPortStatus_1_PRSC_reg <= 1'b0;
    end
    if(reg_hcRhPortStatus_1_PRSC_set) begin
      reg_hcRhPortStatus_1_PRSC_reg <= 1'b1;
    end
    if(reg_hcRhPortStatus_1_PRSC_set) begin
      reg_hcInterrupt_RHSC_status <= 1'b1;
    end
    if(when_UsbOhci_l448_3) begin
      reg_hcRhPortStatus_1_PES <= 1'b0;
    end
    if(when_UsbOhci_l448_4) begin
      reg_hcRhPortStatus_1_PES <= 1'b1;
    end
    if(when_UsbOhci_l448_5) begin
      reg_hcRhPortStatus_1_PES <= 1'b1;
    end
    if(when_UsbOhci_l449_2) begin
      reg_hcRhPortStatus_1_PSS <= 1'b0;
    end
    if(when_UsbOhci_l449_3) begin
      reg_hcRhPortStatus_1_PSS <= 1'b1;
    end
    if(when_UsbOhci_l450_1) begin
      reg_hcRhPortStatus_1_suspend <= 1'b1;
    end
    if(when_UsbOhci_l451_1) begin
      reg_hcRhPortStatus_1_resume <= 1'b1;
    end
    if(when_UsbOhci_l452_1) begin
      reg_hcRhPortStatus_1_reset <= 1'b1;
    end
    if(reg_hcRhDescriptorA_NPS) begin
      reg_hcRhPortStatus_1_PPS <= 1'b1;
    end else begin
      if(reg_hcRhDescriptorA_PSM) begin
        if(when_UsbOhci_l458_1) begin
          if(reg_hcRhPortStatus_1_clearPortPower) begin
            reg_hcRhPortStatus_1_PPS <= 1'b0;
          end
          if(reg_hcRhPortStatus_1_setPortPower) begin
            reg_hcRhPortStatus_1_PPS <= 1'b1;
          end
        end else begin
          if(reg_hcRhStatus_clearGlobalPower) begin
            reg_hcRhPortStatus_1_PPS <= 1'b0;
          end
          if(reg_hcRhStatus_setGlobalPower) begin
            reg_hcRhPortStatus_1_PPS <= 1'b1;
          end
        end
      end else begin
        if(reg_hcRhStatus_clearGlobalPower) begin
          reg_hcRhPortStatus_1_PPS <= 1'b0;
        end
        if(reg_hcRhStatus_setGlobalPower) begin
          reg_hcRhPortStatus_1_PPS <= 1'b1;
        end
      end
    end
    if(io_phy_ports_1_resume_fire) begin
      reg_hcRhPortStatus_1_resume <= 1'b0;
    end
    if(io_phy_ports_1_reset_fire) begin
      reg_hcRhPortStatus_1_reset <= 1'b0;
    end
    if(io_phy_ports_1_suspend_fire) begin
      reg_hcRhPortStatus_1_suspend <= 1'b0;
    end
    frame_decrementTimer <= (frame_decrementTimer + 3'b001);
    if(frame_decrementTimerOverflow) begin
      frame_decrementTimer <= 3'b000;
    end
    if(when_UsbOhci_l514) begin
      reg_hcFmRemaining_FR <= (reg_hcFmRemaining_FR - 14'h0001);
      if(when_UsbOhci_l516) begin
        frame_limitCounter <= (frame_limitCounter - 15'h0001);
      end
    end
    if(frame_reload) begin
      reg_hcFmRemaining_FR <= reg_hcFmInterval_FI;
      reg_hcFmRemaining_FRT <= reg_hcFmInterval_FIT;
      reg_hcFmNumber_FN <= reg_hcFmNumber_FNp1;
      frame_limitCounter <= reg_hcFmInterval_FSMPS;
      frame_decrementTimer <= 3'b000;
    end
    if(io_phy_tick) begin
      rxTimer_counter <= (rxTimer_counter + 8'h01);
    end
    if(rxTimer_clear) begin
      rxTimer_counter <= 8'h0;
    end
    if(_zz_2) begin
      _zz_dataRx_history_0 <= _zz_dataRx_pid;
    end
    if(_zz_2) begin
      _zz_dataRx_history_1 <= _zz_dataRx_history_0;
    end
    if(priority_tick) begin
      priority_counter <= (priority_counter + 2'b01);
    end
    if(priority_skip) begin
      priority_bulk <= (! priority_bulk);
      priority_counter <= 2'b00;
    end
    endpoint_TD_isoOverrunReg <= endpoint_TD_isoOverrun;
    endpoint_TD_isoZero <= (endpoint_TD_isoLast ? (endpoint_TD_isoBaseNext < endpoint_TD_isoBase) : (endpoint_TD_isoBase == endpoint_TD_isoBaseNext));
    endpoint_TD_isoLastReg <= endpoint_TD_isoLast;
    endpoint_TD_tooEarlyReg <= endpoint_TD_tooEarly;
    endpoint_TD_lastOffset <= (endpoint_ED_F ? _zz_endpoint_TD_lastOffset : {(! endpoint_TD_isSinglePage),endpoint_TD_BE[11 : 0]});
    if(endpoint_TD_clear) begin
      endpoint_TD_retire <= 1'b0;
      endpoint_TD_dataPhaseUpdate <= 1'b0;
      endpoint_TD_upateCBP <= 1'b0;
      endpoint_TD_noUpdate <= 1'b0;
    end
    if(endpoint_applyNextED) begin
      case(endpoint_flowType)
        FlowType_BULK : begin
          reg_hcBulkCurrentED_BCED_reg <= endpoint_ED_nextED;
        end
        FlowType_CONTROL : begin
          reg_hcControlCurrentED_CCED_reg <= endpoint_ED_nextED;
        end
        default : begin
          reg_hcPeriodCurrentED_PCED_reg <= endpoint_ED_nextED;
        end
      endcase
    end
    if(when_UsbOhci_l937) begin
      endpoint_dmaLogic_storage_writePtr <= (endpoint_dmaLogic_storage_writePtr + 7'h01);
    end
    if(endpoint_dmaLogic_byteCtx_increment) begin
      endpoint_dmaLogic_byteCtx_counter <= (endpoint_dmaLogic_byteCtx_counter + 13'h0001);
    end
    if(endpoint_dmaLogic_fromUsb_push) begin
      endpoint_dmaLogic_storage_writePtr <= (endpoint_dmaLogic_storage_writePtr + 7'h01);
    end
    if(endpoint_dmaLogic_fromUsb_run) begin
      if(dataRx_wantExit) begin
        endpoint_dmaLogic_underflow <= when_UsbOhci_l1011;
        endpoint_dmaLogic_overflow <= ((! when_UsbOhci_l1011) && (_zz_endpoint_dmaLogic_overflow != endpoint_dmaLogic_fromUsb_transactionSizeMax));
        if(endpoint_zeroLength) begin
          endpoint_dmaLogic_underflow <= 1'b0;
          endpoint_dmaLogic_overflow <= (endpoint_dmaLogic_fromUsbCounter != 11'h0);
        end
        if(when_UsbOhci_l1011) begin
          endpoint_lastAddress <= (_zz_endpoint_lastAddress_1 - 13'h0001);
        end
      end
      if(dataRx_data_valid) begin
        endpoint_dmaLogic_fromUsbCounter <= (endpoint_dmaLogic_fromUsbCounter + _zz_endpoint_dmaLogic_fromUsbCounter);
        if(_zz_5[0]) begin
          endpoint_dmaLogic_fromUsb_buffer[7 : 0] <= dataRx_data_payload;
        end
        if(_zz_5[1]) begin
          endpoint_dmaLogic_fromUsb_buffer[15 : 8] <= dataRx_data_payload;
        end
        if(_zz_5[2]) begin
          endpoint_dmaLogic_fromUsb_buffer[23 : 16] <= dataRx_data_payload;
        end
        if(_zz_5[3]) begin
          endpoint_dmaLogic_fromUsb_buffer[31 : 24] <= dataRx_data_payload;
        end
      end
    end
    case(io_ctrl_cmd_payload_fragment_address)
      12'h004 : begin
        if(ctrl_doWrite) begin
          if(when_BusSlaveFactory_l1041) begin
            reg_hcControl_CBSR[1 : 0] <= io_ctrl_cmd_payload_fragment_data[1 : 0];
          end
          if(when_BusSlaveFactory_l1041_1) begin
            reg_hcControl_PLE <= io_ctrl_cmd_payload_fragment_data[2];
          end
          if(when_BusSlaveFactory_l1041_2) begin
            reg_hcControl_IE <= io_ctrl_cmd_payload_fragment_data[3];
          end
          if(when_BusSlaveFactory_l1041_3) begin
            reg_hcControl_CLE <= io_ctrl_cmd_payload_fragment_data[4];
          end
          if(when_BusSlaveFactory_l1041_4) begin
            reg_hcControl_BLE <= io_ctrl_cmd_payload_fragment_data[5];
          end
          if(when_BusSlaveFactory_l1041_7) begin
            reg_hcControl_RWE <= io_ctrl_cmd_payload_fragment_data[10];
          end
        end
      end
      12'h018 : begin
        if(ctrl_doWrite) begin
          if(when_BusSlaveFactory_l1041_8) begin
            reg_hcHCCA_HCCA_reg[7 : 0] <= io_ctrl_cmd_payload_fragment_data[15 : 8];
          end
          if(when_BusSlaveFactory_l1041_9) begin
            reg_hcHCCA_HCCA_reg[15 : 8] <= io_ctrl_cmd_payload_fragment_data[23 : 16];
          end
          if(when_BusSlaveFactory_l1041_10) begin
            reg_hcHCCA_HCCA_reg[23 : 16] <= io_ctrl_cmd_payload_fragment_data[31 : 24];
          end
        end
      end
      12'h020 : begin
        if(ctrl_doWrite) begin
          if(when_BusSlaveFactory_l1041_11) begin
            reg_hcControlHeadED_CHED_reg[3 : 0] <= io_ctrl_cmd_payload_fragment_data[7 : 4];
          end
          if(when_BusSlaveFactory_l1041_12) begin
            reg_hcControlHeadED_CHED_reg[11 : 4] <= io_ctrl_cmd_payload_fragment_data[15 : 8];
          end
          if(when_BusSlaveFactory_l1041_13) begin
            reg_hcControlHeadED_CHED_reg[19 : 12] <= io_ctrl_cmd_payload_fragment_data[23 : 16];
          end
          if(when_BusSlaveFactory_l1041_14) begin
            reg_hcControlHeadED_CHED_reg[27 : 20] <= io_ctrl_cmd_payload_fragment_data[31 : 24];
          end
        end
      end
      12'h024 : begin
        if(ctrl_doWrite) begin
          if(when_BusSlaveFactory_l1041_15) begin
            reg_hcControlCurrentED_CCED_reg[3 : 0] <= io_ctrl_cmd_payload_fragment_data[7 : 4];
          end
          if(when_BusSlaveFactory_l1041_16) begin
            reg_hcControlCurrentED_CCED_reg[11 : 4] <= io_ctrl_cmd_payload_fragment_data[15 : 8];
          end
          if(when_BusSlaveFactory_l1041_17) begin
            reg_hcControlCurrentED_CCED_reg[19 : 12] <= io_ctrl_cmd_payload_fragment_data[23 : 16];
          end
          if(when_BusSlaveFactory_l1041_18) begin
            reg_hcControlCurrentED_CCED_reg[27 : 20] <= io_ctrl_cmd_payload_fragment_data[31 : 24];
          end
        end
      end
      12'h028 : begin
        if(ctrl_doWrite) begin
          if(when_BusSlaveFactory_l1041_19) begin
            reg_hcBulkHeadED_BHED_reg[3 : 0] <= io_ctrl_cmd_payload_fragment_data[7 : 4];
          end
          if(when_BusSlaveFactory_l1041_20) begin
            reg_hcBulkHeadED_BHED_reg[11 : 4] <= io_ctrl_cmd_payload_fragment_data[15 : 8];
          end
          if(when_BusSlaveFactory_l1041_21) begin
            reg_hcBulkHeadED_BHED_reg[19 : 12] <= io_ctrl_cmd_payload_fragment_data[23 : 16];
          end
          if(when_BusSlaveFactory_l1041_22) begin
            reg_hcBulkHeadED_BHED_reg[27 : 20] <= io_ctrl_cmd_payload_fragment_data[31 : 24];
          end
        end
      end
      12'h02c : begin
        if(ctrl_doWrite) begin
          if(when_BusSlaveFactory_l1041_23) begin
            reg_hcBulkCurrentED_BCED_reg[3 : 0] <= io_ctrl_cmd_payload_fragment_data[7 : 4];
          end
          if(when_BusSlaveFactory_l1041_24) begin
            reg_hcBulkCurrentED_BCED_reg[11 : 4] <= io_ctrl_cmd_payload_fragment_data[15 : 8];
          end
          if(when_BusSlaveFactory_l1041_25) begin
            reg_hcBulkCurrentED_BCED_reg[19 : 12] <= io_ctrl_cmd_payload_fragment_data[23 : 16];
          end
          if(when_BusSlaveFactory_l1041_26) begin
            reg_hcBulkCurrentED_BCED_reg[27 : 20] <= io_ctrl_cmd_payload_fragment_data[31 : 24];
          end
        end
      end
      12'h030 : begin
        if(ctrl_doWrite) begin
          if(when_BusSlaveFactory_l1041_27) begin
            reg_hcDoneHead_DH_reg[3 : 0] <= io_ctrl_cmd_payload_fragment_data[7 : 4];
          end
          if(when_BusSlaveFactory_l1041_28) begin
            reg_hcDoneHead_DH_reg[11 : 4] <= io_ctrl_cmd_payload_fragment_data[15 : 8];
          end
          if(when_BusSlaveFactory_l1041_29) begin
            reg_hcDoneHead_DH_reg[19 : 12] <= io_ctrl_cmd_payload_fragment_data[23 : 16];
          end
          if(when_BusSlaveFactory_l1041_30) begin
            reg_hcDoneHead_DH_reg[27 : 20] <= io_ctrl_cmd_payload_fragment_data[31 : 24];
          end
        end
      end
      12'h034 : begin
        if(ctrl_doWrite) begin
          if(when_BusSlaveFactory_l1041_31) begin
            reg_hcFmInterval_FI[7 : 0] <= io_ctrl_cmd_payload_fragment_data[7 : 0];
          end
          if(when_BusSlaveFactory_l1041_32) begin
            reg_hcFmInterval_FI[13 : 8] <= io_ctrl_cmd_payload_fragment_data[13 : 8];
          end
          if(when_BusSlaveFactory_l1041_33) begin
            reg_hcFmInterval_FSMPS[7 : 0] <= io_ctrl_cmd_payload_fragment_data[23 : 16];
          end
          if(when_BusSlaveFactory_l1041_34) begin
            reg_hcFmInterval_FSMPS[14 : 8] <= io_ctrl_cmd_payload_fragment_data[30 : 24];
          end
          if(when_BusSlaveFactory_l1041_35) begin
            reg_hcFmInterval_FIT <= io_ctrl_cmd_payload_fragment_data[31];
          end
        end
      end
      12'h044 : begin
        if(ctrl_doWrite) begin
          if(when_BusSlaveFactory_l1041_38) begin
            reg_hcLSThreshold_LST[7 : 0] <= io_ctrl_cmd_payload_fragment_data[7 : 0];
          end
          if(when_BusSlaveFactory_l1041_39) begin
            reg_hcLSThreshold_LST[11 : 8] <= io_ctrl_cmd_payload_fragment_data[11 : 8];
          end
        end
      end
      12'h048 : begin
        if(ctrl_doWrite) begin
          if(when_BusSlaveFactory_l1041_40) begin
            reg_hcRhDescriptorA_PSM <= io_ctrl_cmd_payload_fragment_data[8];
          end
          if(when_BusSlaveFactory_l1041_41) begin
            reg_hcRhDescriptorA_NPS <= io_ctrl_cmd_payload_fragment_data[9];
          end
          if(when_BusSlaveFactory_l1041_42) begin
            reg_hcRhDescriptorA_OCPM <= io_ctrl_cmd_payload_fragment_data[11];
          end
          if(when_BusSlaveFactory_l1041_43) begin
            reg_hcRhDescriptorA_NOCP <= io_ctrl_cmd_payload_fragment_data[12];
          end
          if(when_BusSlaveFactory_l1041_44) begin
            reg_hcRhDescriptorA_POTPGT[7 : 0] <= io_ctrl_cmd_payload_fragment_data[31 : 24];
          end
        end
      end
      12'h04c : begin
        if(ctrl_doWrite) begin
          if(when_BusSlaveFactory_l1041_45) begin
            reg_hcRhDescriptorB_DR[1 : 0] <= io_ctrl_cmd_payload_fragment_data[2 : 1];
          end
          if(when_BusSlaveFactory_l1041_46) begin
            reg_hcRhDescriptorB_PPCM[1 : 0] <= io_ctrl_cmd_payload_fragment_data[18 : 17];
          end
        end
      end
      default : begin
      end
    endcase
    if(when_UsbOhci_l241) begin
      reg_hcControl_CBSR <= 2'b00;
      reg_hcControl_PLE <= 1'b0;
      reg_hcControl_IE <= 1'b0;
      reg_hcControl_CLE <= 1'b0;
      reg_hcControl_BLE <= 1'b0;
      reg_hcControl_RWE <= 1'b0;
      reg_hcCommandStatus_CLF <= 1'b0;
      reg_hcCommandStatus_BLF <= 1'b0;
      reg_hcCommandStatus_OCR <= 1'b0;
      reg_hcCommandStatus_SOC <= 2'b00;
      reg_hcInterrupt_MIE <= 1'b0;
      reg_hcInterrupt_SO_status <= 1'b0;
      reg_hcInterrupt_SO_enable <= 1'b0;
      reg_hcInterrupt_WDH_status <= 1'b0;
      reg_hcInterrupt_WDH_enable <= 1'b0;
      reg_hcInterrupt_SF_status <= 1'b0;
      reg_hcInterrupt_SF_enable <= 1'b0;
      reg_hcInterrupt_RD_status <= 1'b0;
      reg_hcInterrupt_RD_enable <= 1'b0;
      reg_hcInterrupt_UE_status <= 1'b0;
      reg_hcInterrupt_UE_enable <= 1'b0;
      reg_hcInterrupt_FNO_status <= 1'b0;
      reg_hcInterrupt_FNO_enable <= 1'b0;
      reg_hcInterrupt_RHSC_status <= 1'b0;
      reg_hcInterrupt_RHSC_enable <= 1'b0;
      reg_hcInterrupt_OC_status <= 1'b0;
      reg_hcInterrupt_OC_enable <= 1'b0;
      reg_hcHCCA_HCCA_reg <= 24'h0;
      reg_hcPeriodCurrentED_PCED_reg <= 28'h0;
      reg_hcControlHeadED_CHED_reg <= 28'h0;
      reg_hcControlCurrentED_CCED_reg <= 28'h0;
      reg_hcBulkHeadED_BHED_reg <= 28'h0;
      reg_hcBulkCurrentED_BCED_reg <= 28'h0;
      reg_hcDoneHead_DH_reg <= 28'h0;
      reg_hcFmInterval_FI <= 14'h2edf;
      reg_hcFmInterval_FIT <= 1'b0;
      reg_hcFmRemaining_FR <= 14'h0;
      reg_hcFmRemaining_FRT <= 1'b0;
      reg_hcFmNumber_FN <= 16'h0;
      reg_hcLSThreshold_LST <= 12'h628;
      reg_hcRhDescriptorA_PSM <= 1'b1;
      reg_hcRhDescriptorA_NPS <= 1'b1;
      reg_hcRhDescriptorA_OCPM <= 1'b1;
      reg_hcRhDescriptorA_NOCP <= 1'b1;
      reg_hcRhDescriptorA_POTPGT <= 8'h0a;
      reg_hcRhDescriptorB_DR <= {1'b0,1'b0};
      reg_hcRhDescriptorB_PPCM <= {1'b1,1'b1};
      reg_hcRhStatus_DRWE <= 1'b0;
      reg_hcRhStatus_CCIC <= 1'b0;
      reg_hcRhPortStatus_0_resume <= 1'b0;
      reg_hcRhPortStatus_0_reset <= 1'b0;
      reg_hcRhPortStatus_0_suspend <= 1'b0;
      reg_hcRhPortStatus_0_PSS <= 1'b0;
      reg_hcRhPortStatus_0_PPS <= 1'b0;
      reg_hcRhPortStatus_0_PES <= 1'b0;
      reg_hcRhPortStatus_0_CSC_reg <= 1'b0;
      reg_hcRhPortStatus_0_PESC_reg <= 1'b0;
      reg_hcRhPortStatus_0_PSSC_reg <= 1'b0;
      reg_hcRhPortStatus_0_OCIC_reg <= 1'b0;
      reg_hcRhPortStatus_0_PRSC_reg <= 1'b0;
      reg_hcRhPortStatus_1_resume <= 1'b0;
      reg_hcRhPortStatus_1_reset <= 1'b0;
      reg_hcRhPortStatus_1_suspend <= 1'b0;
      reg_hcRhPortStatus_1_PSS <= 1'b0;
      reg_hcRhPortStatus_1_PPS <= 1'b0;
      reg_hcRhPortStatus_1_PES <= 1'b0;
      reg_hcRhPortStatus_1_CSC_reg <= 1'b0;
      reg_hcRhPortStatus_1_PESC_reg <= 1'b0;
      reg_hcRhPortStatus_1_PSSC_reg <= 1'b0;
      reg_hcRhPortStatus_1_OCIC_reg <= 1'b0;
      reg_hcRhPortStatus_1_PRSC_reg <= 1'b0;
    end
    case(dataRx_stateReg)
      dataRx_enumDef_IDLE : begin
        if(!io_phy_rx_active) begin
          if(rxTimer_rxTimeout) begin
            dataRx_notResponding <= 1'b1;
          end
        end
      end
      dataRx_enumDef_PID : begin
        dataRx_valids <= 2'b00;
        dataRx_pidError <= 1'b1;
        if(_zz_2) begin
          dataRx_pid <= _zz_dataRx_pid[3 : 0];
          dataRx_pidError <= (_zz_dataRx_pid[3 : 0] != (~ _zz_dataRx_pid[7 : 4]));
        end
      end
      dataRx_enumDef_DATA : begin
        if(when_Misc_l70) begin
          if(when_Misc_l71) begin
            dataRx_crcError <= 1'b1;
          end
        end else begin
          if(_zz_2) begin
            dataRx_valids <= {dataRx_valids[0],1'b1};
          end
        end
      end
      default : begin
      end
    endcase
    if(when_StateMachine_l253) begin
      dataRx_notResponding <= 1'b0;
      dataRx_stuffingError <= 1'b0;
      dataRx_pidError <= 1'b0;
      dataRx_crcError <= 1'b0;
    end
    if(when_Misc_l85) begin
      if(_zz_2) begin
        if(when_Misc_l87) begin
          dataRx_stuffingError <= 1'b1;
        end
      end
    end
    case(sof_stateReg)
      sof_enumDef_FRAME_TX : begin
        sof_doInterruptDelay <= (interruptDelay_done && (! reg_hcInterrupt_WDH_status));
      end
      sof_enumDef_FRAME_NUMBER_CMD : begin
      end
      sof_enumDef_FRAME_NUMBER_RSP : begin
        if(ioDma_rsp_valid) begin
          reg_hcInterrupt_SF_status <= 1'b1;
          if(reg_hcFmNumber_overflow) begin
            reg_hcInterrupt_FNO_status <= 1'b1;
          end
          if(sof_doInterruptDelay) begin
            reg_hcInterrupt_WDH_status <= 1'b1;
            reg_hcDoneHead_DH_reg <= 28'h0;
          end
        end
      end
      default : begin
      end
    endcase
    case(endpoint_stateReg)
      endpoint_enumDef_ED_READ_CMD : begin
      end
      endpoint_enumDef_ED_READ_RSP : begin
        if(when_UsbOhci_l189) begin
          endpoint_ED_words_0 <= dmaRspMux_vec_0[31 : 0];
        end
        if(when_UsbOhci_l189_1) begin
          endpoint_ED_words_1 <= dmaRspMux_vec_0[31 : 0];
        end
        if(when_UsbOhci_l189_2) begin
          endpoint_ED_words_2 <= dmaRspMux_vec_0[31 : 0];
        end
        if(when_UsbOhci_l189_3) begin
          endpoint_ED_words_3 <= dmaRspMux_vec_0[31 : 0];
        end
      end
      endpoint_enumDef_ED_ANALYSE : begin
      end
      endpoint_enumDef_TD_READ_CMD : begin
      end
      endpoint_enumDef_TD_READ_RSP : begin
        if(when_UsbOhci_l189_4) begin
          endpoint_TD_words_0 <= dmaRspMux_vec_0[31 : 0];
        end
        if(when_UsbOhci_l189_5) begin
          endpoint_TD_words_1 <= dmaRspMux_vec_0[31 : 0];
        end
        if(when_UsbOhci_l189_6) begin
          endpoint_TD_words_2 <= dmaRspMux_vec_0[31 : 0];
        end
        if(when_UsbOhci_l189_7) begin
          endpoint_TD_words_3 <= dmaRspMux_vec_0[31 : 0];
        end
        if(when_UsbOhci_l879) begin
          if(when_UsbOhci_l189_8) begin
            endpoint_TD_isoBase <= dmaRspMux_vec_0[12 : 0];
          end
          if(when_UsbOhci_l189_9) begin
            endpoint_TD_isoBaseNext <= dmaRspMux_vec_0[28 : 16];
          end
        end
        if(when_UsbOhci_l879_1) begin
          if(when_UsbOhci_l189_10) begin
            endpoint_TD_isoBase <= dmaRspMux_vec_0[28 : 16];
          end
          if(when_UsbOhci_l189_11) begin
            endpoint_TD_isoBaseNext <= dmaRspMux_vec_0[12 : 0];
          end
        end
        if(when_UsbOhci_l879_2) begin
          if(when_UsbOhci_l189_12) begin
            endpoint_TD_isoBase <= dmaRspMux_vec_0[12 : 0];
          end
          if(when_UsbOhci_l189_13) begin
            endpoint_TD_isoBaseNext <= dmaRspMux_vec_0[28 : 16];
          end
        end
        if(when_UsbOhci_l879_3) begin
          if(when_UsbOhci_l189_14) begin
            endpoint_TD_isoBase <= dmaRspMux_vec_0[28 : 16];
          end
          if(when_UsbOhci_l189_15) begin
            endpoint_TD_isoBaseNext <= dmaRspMux_vec_0[12 : 0];
          end
        end
        if(when_UsbOhci_l879_4) begin
          if(when_UsbOhci_l189_16) begin
            endpoint_TD_isoBase <= dmaRspMux_vec_0[12 : 0];
          end
          if(when_UsbOhci_l189_17) begin
            endpoint_TD_isoBaseNext <= dmaRspMux_vec_0[28 : 16];
          end
        end
        if(when_UsbOhci_l879_5) begin
          if(when_UsbOhci_l189_18) begin
            endpoint_TD_isoBase <= dmaRspMux_vec_0[28 : 16];
          end
          if(when_UsbOhci_l189_19) begin
            endpoint_TD_isoBaseNext <= dmaRspMux_vec_0[12 : 0];
          end
        end
        if(when_UsbOhci_l879_6) begin
          if(when_UsbOhci_l189_20) begin
            endpoint_TD_isoBase <= dmaRspMux_vec_0[12 : 0];
          end
          if(when_UsbOhci_l189_21) begin
            endpoint_TD_isoBaseNext <= dmaRspMux_vec_0[28 : 16];
          end
        end
        if(when_UsbOhci_l879_7) begin
          if(when_UsbOhci_l189_22) begin
            endpoint_TD_isoBase <= dmaRspMux_vec_0[28 : 16];
          end
        end
        if(endpoint_TD_isoLast) begin
          endpoint_TD_isoBaseNext <= {(! endpoint_TD_isSinglePage),endpoint_TD_BE[11 : 0]};
        end
      end
      endpoint_enumDef_TD_READ_DELAY : begin
      end
      endpoint_enumDef_TD_ANALYSE : begin
        case(endpoint_flowType)
          FlowType_CONTROL : begin
            reg_hcCommandStatus_CLF <= 1'b1;
          end
          FlowType_BULK : begin
            reg_hcCommandStatus_BLF <= 1'b1;
          end
          default : begin
          end
        endcase
        endpoint_dmaLogic_byteCtx_counter <= endpoint_TD_firstOffset;
        endpoint_currentAddress <= {1'd0, endpoint_TD_firstOffset};
        endpoint_lastAddress <= _zz_endpoint_lastAddress_3[12:0];
        endpoint_zeroLength <= (endpoint_ED_F ? endpoint_TD_isoZero : (endpoint_TD_CBP == 32'h0));
        endpoint_dataPhase <= (endpoint_ED_F ? 1'b0 : (endpoint_TD_T[1] ? endpoint_TD_T[0] : endpoint_ED_C));
        if(endpoint_ED_F) begin
          if(endpoint_TD_isoOverrunReg) begin
            endpoint_TD_retire <= 1'b1;
          end
        end
      end
      endpoint_enumDef_TD_CHECK_TIME : begin
        if(endpoint_timeCheck) begin
          endpoint_status_1 <= endpoint_Status_FRAME_TIME;
        end
      end
      endpoint_enumDef_BUFFER_READ : begin
        if(endpoint_dmaLogic_toUsb_run) begin
          if(endpoint_timeCheck) begin
            endpoint_status_1 <= endpoint_Status_FRAME_TIME;
          end
        end
      end
      endpoint_enumDef_TOKEN : begin
      end
      endpoint_enumDef_DATA_TX : begin
        if(dataTx_wantExit) begin
          if(endpoint_ED_F) begin
            endpoint_TD_words_0[31 : 28] <= 4'b0000;
          end
        end
      end
      endpoint_enumDef_DATA_RX : begin
      end
      endpoint_enumDef_DATA_RX_VALIDATE : begin
        endpoint_TD_words_0[31 : 28] <= 4'b0000;
        if(dataRx_notResponding) begin
          endpoint_TD_words_0[31 : 28] <= 4'b0101;
        end else begin
          if(dataRx_stuffingError) begin
            endpoint_TD_words_0[31 : 28] <= 4'b0010;
          end else begin
            if(dataRx_pidError) begin
              endpoint_TD_words_0[31 : 28] <= 4'b0110;
            end else begin
              if(endpoint_ED_F) begin
                case(dataRx_pid)
                  4'b1110, 4'b1010 : begin
                    endpoint_TD_words_0[31 : 28] <= 4'b0100;
                  end
                  4'b0011, 4'b1011 : begin
                  end
                  default : begin
                    endpoint_TD_words_0[31 : 28] <= 4'b0111;
                  end
                endcase
              end else begin
                case(dataRx_pid)
                  4'b1010 : begin
                    endpoint_TD_noUpdate <= 1'b1;
                  end
                  4'b1110 : begin
                    endpoint_TD_words_0[31 : 28] <= 4'b0100;
                  end
                  4'b0011, 4'b1011 : begin
                    if(when_UsbOhci_l1318) begin
                      endpoint_TD_words_0[31 : 28] <= 4'b0011;
                    end
                  end
                  default : begin
                    endpoint_TD_words_0[31 : 28] <= 4'b0111;
                  end
                endcase
              end
              if(when_UsbOhci_l1329) begin
                if(dataRx_crcError) begin
                  endpoint_TD_words_0[31 : 28] <= 4'b0001;
                end else begin
                  if(endpoint_dmaLogic_underflowError) begin
                    endpoint_TD_words_0[31 : 28] <= 4'b1001;
                  end else begin
                    if(endpoint_dmaLogic_overflow) begin
                      endpoint_TD_words_0[31 : 28] <= 4'b1000;
                    end
                  end
                end
              end
            end
          end
        end
      end
      endpoint_enumDef_ACK_RX : begin
        if(io_phy_rx_flow_valid) begin
          endpoint_ackRxFired <= 1'b1;
          endpoint_ackRxPid <= io_phy_rx_flow_payload_data[3 : 0];
          if(io_phy_rx_flow_payload_stuffingError) begin
            endpoint_ackRxStuffing <= 1'b1;
          end
          if(when_UsbOhci_l1255) begin
            endpoint_ackRxPidFailure <= 1'b1;
          end
        end
        if(io_phy_rx_active) begin
          endpoint_ackRxActivated <= 1'b1;
        end
        if(when_UsbOhci_l1260) begin
          if(when_UsbOhci_l1262) begin
            endpoint_TD_words_0[31 : 28] <= 4'b0110;
          end else begin
            if(endpoint_ackRxStuffing) begin
              endpoint_TD_words_0[31 : 28] <= 4'b0010;
            end else begin
              if(endpoint_ackRxPidFailure) begin
                endpoint_TD_words_0[31 : 28] <= 4'b0110;
              end else begin
                case(endpoint_ackRxPid)
                  4'b0010 : begin
                    endpoint_TD_words_0[31 : 28] <= 4'b0000;
                  end
                  4'b1010 : begin
                  end
                  4'b1110 : begin
                    endpoint_TD_words_0[31 : 28] <= 4'b0100;
                  end
                  default : begin
                    endpoint_TD_words_0[31 : 28] <= 4'b0111;
                  end
                endcase
              end
            end
          end
        end
        if(rxTimer_rxTimeout) begin
          endpoint_TD_words_0[31 : 28] <= 4'b0101;
        end
      end
      endpoint_enumDef_ACK_TX_0 : begin
      end
      endpoint_enumDef_ACK_TX_1 : begin
      end
      endpoint_enumDef_ACK_TX_EOP : begin
      end
      endpoint_enumDef_DATA_RX_WAIT_DMA : begin
      end
      endpoint_enumDef_UPDATE_TD_PROCESS : begin
        if(endpoint_ED_F) begin
          if(endpoint_TD_isoLastReg) begin
            endpoint_TD_retire <= 1'b1;
          end
        end else begin
          endpoint_TD_words_0[27 : 26] <= 2'b00;
          case(endpoint_TD_CC)
            4'b0000 : begin
              if(when_UsbOhci_l1386) begin
                endpoint_TD_retire <= 1'b1;
              end
              endpoint_TD_dataPhaseUpdate <= 1'b1;
              endpoint_TD_upateCBP <= 1'b1;
            end
            4'b1001 : begin
              endpoint_TD_retire <= 1'b1;
              endpoint_TD_dataPhaseUpdate <= 1'b1;
              endpoint_TD_upateCBP <= 1'b1;
            end
            4'b1000 : begin
              endpoint_TD_retire <= 1'b1;
              endpoint_TD_dataPhaseUpdate <= 1'b1;
            end
            4'b0010, 4'b0001, 4'b0110, 4'b0101, 4'b0111, 4'b0011 : begin
              endpoint_TD_words_0[27 : 26] <= _zz_endpoint_TD_words_0;
              if(when_UsbOhci_l1401) begin
                endpoint_TD_words_0[31 : 28] <= 4'b0000;
              end else begin
                endpoint_TD_retire <= 1'b1;
              end
            end
            default : begin
              endpoint_TD_retire <= 1'b1;
            end
          endcase
          if(endpoint_TD_noUpdate) begin
            endpoint_TD_retire <= 1'b0;
          end
        end
      end
      endpoint_enumDef_UPDATE_TD_CMD : begin
        endpoint_ED_words_2[0] <= ((! endpoint_ED_F) && (endpoint_TD_CC != 4'b0000));
      end
      endpoint_enumDef_UPDATE_ED_CMD : begin
      end
      endpoint_enumDef_UPDATE_SYNC : begin
        if(dmaCtx_pendingEmpty) begin
          if(endpoint_TD_retire) begin
            reg_hcDoneHead_DH_reg <= endpoint_ED_headP;
          end
        end
      end
      endpoint_enumDef_ABORD : begin
      end
      default : begin
      end
    endcase
    if(when_StateMachine_l237_2) begin
      endpoint_status_1 <= endpoint_Status_OK;
    end
    if(when_StateMachine_l253_4) begin
      endpoint_ackRxFired <= 1'b0;
      endpoint_ackRxActivated <= 1'b0;
      endpoint_ackRxPidFailure <= 1'b0;
      endpoint_ackRxStuffing <= 1'b0;
    end
    case(endpoint_dmaLogic_stateReg)
      endpoint_dmaLogic_enumDef_INIT : begin
        endpoint_dmaLogic_underflow <= 1'b0;
        endpoint_dmaLogic_overflow <= 1'b0;
        if(endpoint_isIn) begin
          endpoint_dmaLogic_fromUsbCounter <= 11'h0;
          endpoint_dmaLogic_storage_writePtr <= _zz_endpoint_dmaLogic_storage_writePtr[6:0];
          endpoint_dmaLogic_storage_readPtr <= _zz_endpoint_dmaLogic_storage_readPtr[6:0];
        end else begin
          endpoint_dmaLogic_storage_writePtr <= _zz_endpoint_dmaLogic_storage_writePtr_1[6:0];
          endpoint_dmaLogic_storage_readPtr <= _zz_endpoint_dmaLogic_storage_readPtr_3[6:0];
        end
        endpoint_dmaLogic_fromUsb_transactionSizeMax <= (_zz_endpoint_dmaLogic_fromUsb_transactionSizeMax + 14'h0001);
      end
      endpoint_dmaLogic_enumDef_TO_USB : begin
      end
      endpoint_dmaLogic_enumDef_FROM_USB : begin
      end
      endpoint_dmaLogic_enumDef_VALIDATION : begin
      end
      endpoint_dmaLogic_enumDef_CALC_CMD : begin
        endpoint_dmaLogic_length <= endpoint_dmaLogic_lengthCalc;
      end
      endpoint_dmaLogic_enumDef_READ_CMD : begin
        if(ioDma_cmd_ready) begin
          endpoint_currentAddress <= (_zz_endpoint_currentAddress + 14'h0001);
        end
      end
      endpoint_dmaLogic_enumDef_WRITE_CMD : begin
        if(when_UsbOhci_l1093) begin
          if(endpoint_dmaLogic_storage_readCmd_ready) begin
            endpoint_dmaLogic_storage_readPtr <= (endpoint_dmaLogic_storage_readPtr + 7'h01);
            if(when_UsbOhci_l1098) begin
              endpoint_dmaLogic_storageReadDone <= 1'b1;
            end
          end
        end
        if(ioDma_cmd_ready) begin
          if(endpoint_dmaLogic_beatLast) begin
            endpoint_currentAddress <= (_zz_endpoint_currentAddress_2 + 14'h0001);
          end
        end
      end
      default : begin
      end
    endcase
    if(when_StateMachine_l253_5) begin
      endpoint_dmaLogic_storageReadDone <= 1'b0;
    end
    if(endpoint_dmaLogic_toUsb_run) begin
      if(endpoint_dmaLogic_storage_readCmd_ready) begin
        endpoint_dmaLogic_storage_readPtr <= (endpoint_dmaLogic_storage_readPtr + 7'h01);
      end
    end
    case(operational_stateReg)
      operational_enumDef_SOF : begin
        if(sof_wantExit) begin
          if(when_UsbOhci_l1516) begin
            reg_hcInterrupt_SO_status <= 1'b1;
            reg_hcCommandStatus_SOC <= (reg_hcCommandStatus_SOC + 2'b01);
          end
          operational_allowBulk <= reg_hcControl_BLE;
          operational_allowControl <= reg_hcControl_CLE;
          operational_allowPeriodic <= reg_hcControl_PLE;
          operational_allowIsochronous <= reg_hcControl_IE;
          operational_periodicDone <= 1'b0;
          operational_periodicHeadFetched <= 1'b0;
          priority_bulk <= 1'b0;
          priority_counter <= 2'b00;
        end
      end
      operational_enumDef_ARBITER : begin
        if(reg_hcControl_BLE) begin
          operational_allowBulk <= 1'b1;
        end
        if(reg_hcControl_CLE) begin
          operational_allowControl <= 1'b1;
        end
        if(!operational_askExit) begin
          if(!frame_limitHit) begin
            if(when_UsbOhci_l1542) begin
              if(!when_UsbOhci_l1543) begin
                if(reg_hcPeriodCurrentED_isZero) begin
                  operational_periodicDone <= 1'b1;
                end else begin
                  endpoint_flowType <= FlowType_PERIODIC;
                  endpoint_ED_address <= reg_hcPeriodCurrentED_PCED_address;
                end
              end
            end else begin
              if(priority_bulk) begin
                if(operational_allowBulk) begin
                  if(reg_hcBulkCurrentED_isZero) begin
                    if(reg_hcCommandStatus_BLF) begin
                      reg_hcBulkCurrentED_BCED_reg <= reg_hcBulkHeadED_BHED_reg;
                      reg_hcCommandStatus_BLF <= 1'b0;
                    end
                  end else begin
                    endpoint_flowType <= FlowType_BULK;
                    endpoint_ED_address <= reg_hcBulkCurrentED_BCED_address;
                  end
                end
              end else begin
                if(operational_allowControl) begin
                  if(reg_hcControlCurrentED_isZero) begin
                    if(reg_hcCommandStatus_CLF) begin
                      reg_hcControlCurrentED_CCED_reg <= reg_hcControlHeadED_CHED_reg;
                      reg_hcCommandStatus_CLF <= 1'b0;
                    end
                  end else begin
                    endpoint_flowType <= FlowType_CONTROL;
                    endpoint_ED_address <= reg_hcControlCurrentED_CCED_address;
                  end
                end
              end
            end
          end
        end
      end
      operational_enumDef_END_POINT : begin
      end
      operational_enumDef_PERIODIC_HEAD_CMD : begin
      end
      operational_enumDef_PERIODIC_HEAD_RSP : begin
        if(ioDma_rsp_valid) begin
          operational_periodicHeadFetched <= 1'b1;
          reg_hcPeriodCurrentED_PCED_reg <= dmaRspMux_data[31 : 4];
        end
      end
      operational_enumDef_WAIT_SOF : begin
      end
      default : begin
      end
    endcase
    if(when_StateMachine_l237_3) begin
      operational_allowPeriodic <= 1'b0;
    end
    case(hc_stateReg)
      hc_enumDef_RESET : begin
      end
      hc_enumDef_RESUME : begin
      end
      hc_enumDef_OPERATIONAL : begin
      end
      hc_enumDef_SUSPEND : begin
        if(when_UsbOhci_l1680) begin
          reg_hcInterrupt_RD_status <= 1'b1;
        end
      end
      hc_enumDef_ANY_TO_RESET : begin
      end
      hc_enumDef_ANY_TO_SUSPEND : begin
      end
      default : begin
      end
    endcase
  end


endmodule

module BufferCC_9 (
  input  wire [1:0]    io_dataIn,
  output wire [1:0]    io_dataOut,
  input  wire          clk_cpu,
  input  wire          ram_axi_cc_toplevel_board_ctrl_reset_ram_synchronized_1
);

  (* async_reg = "true" *) reg        [1:0]    buffers_0;
  (* async_reg = "true" *) reg        [1:0]    buffers_1;

  assign io_dataOut = buffers_1;
  always @(posedge clk_cpu or posedge ram_axi_cc_toplevel_board_ctrl_reset_ram_synchronized_1) begin
    if(ram_axi_cc_toplevel_board_ctrl_reset_ram_synchronized_1) begin
      buffers_0 <= 2'b00;
      buffers_1 <= 2'b00;
    end else begin
      buffers_0 <= io_dataIn;
      buffers_1 <= buffers_0;
    end
  end


endmodule

module BufferCC_8 (
  input  wire [1:0]    io_dataIn,
  output wire [1:0]    io_dataOut,
  input  wire          clk_ram_bus,
  input  wire          reset_ram
);

  (* async_reg = "true" *) reg        [1:0]    buffers_0;
  (* async_reg = "true" *) reg        [1:0]    buffers_1;

  assign io_dataOut = buffers_1;
  always @(posedge clk_ram_bus or posedge reset_ram) begin
    if(reset_ram) begin
      buffers_0 <= 2'b00;
      buffers_1 <= 2'b00;
    end else begin
      buffers_0 <= io_dataIn;
      buffers_1 <= buffers_0;
    end
  end


endmodule

module BufferCC_7 (
  input  wire [4:0]    io_dataIn,
  output wire [4:0]    io_dataOut,
  input  wire          clk_ram_bus,
  input  wire          ram_axi_cc_toplevel_board_ctrl_reset_cpu_synchronized_1
);

  (* async_reg = "true" *) reg        [4:0]    buffers_0;
  (* async_reg = "true" *) reg        [4:0]    buffers_1;

  assign io_dataOut = buffers_1;
  always @(posedge clk_ram_bus or posedge ram_axi_cc_toplevel_board_ctrl_reset_cpu_synchronized_1) begin
    if(ram_axi_cc_toplevel_board_ctrl_reset_cpu_synchronized_1) begin
      buffers_0 <= 5'h0;
      buffers_1 <= 5'h0;
    end else begin
      buffers_0 <= io_dataIn;
      buffers_1 <= buffers_0;
    end
  end


endmodule

module BufferCC_6 (
  input  wire [4:0]    io_dataIn,
  output wire [4:0]    io_dataOut,
  input  wire          clk_cpu,
  input  wire          reset_cpu
);

  (* async_reg = "true" *) reg        [4:0]    buffers_0;
  (* async_reg = "true" *) reg        [4:0]    buffers_1;

  assign io_dataOut = buffers_1;
  always @(posedge clk_cpu or posedge reset_cpu) begin
    if(reset_cpu) begin
      buffers_0 <= 5'h0;
      buffers_1 <= 5'h0;
    end else begin
      buffers_0 <= io_dataIn;
      buffers_1 <= buffers_0;
    end
  end


endmodule

module BufferCC_5 (
  input  wire [7:0]    io_dataIn,
  output wire [7:0]    io_dataOut,
  input  wire          clk_cpu,
  input  wire          ram_axi_cc_toplevel_board_ctrl_reset_ram_synchronized
);

  (* async_reg = "true" *) reg        [7:0]    buffers_0;
  (* async_reg = "true" *) reg        [7:0]    buffers_1;

  assign io_dataOut = buffers_1;
  always @(posedge clk_cpu or posedge ram_axi_cc_toplevel_board_ctrl_reset_ram_synchronized) begin
    if(ram_axi_cc_toplevel_board_ctrl_reset_ram_synchronized) begin
      buffers_0 <= 8'h0;
      buffers_1 <= 8'h0;
    end else begin
      buffers_0 <= io_dataIn;
      buffers_1 <= buffers_0;
    end
  end


endmodule

module BufferCC_4 (
  input  wire          io_dataIn,
  output wire          io_dataOut,
  input  wire          clk_cpu,
  input  wire          reset_ram
);

  (* async_reg = "true" *) reg                 buffers_0;
  (* async_reg = "true" *) reg                 buffers_1;

  assign io_dataOut = buffers_1;
  always @(posedge clk_cpu or posedge reset_ram) begin
    if(reset_ram) begin
      buffers_0 <= 1'b1;
      buffers_1 <= 1'b1;
    end else begin
      buffers_0 <= io_dataIn;
      buffers_1 <= buffers_0;
    end
  end


endmodule

module BufferCC_3 (
  input  wire [7:0]    io_dataIn,
  output wire [7:0]    io_dataOut,
  input  wire          clk_ram_bus,
  input  wire          reset_ram
);

  (* async_reg = "true" *) reg        [7:0]    buffers_0;
  (* async_reg = "true" *) reg        [7:0]    buffers_1;

  assign io_dataOut = buffers_1;
  always @(posedge clk_ram_bus or posedge reset_ram) begin
    if(reset_ram) begin
      buffers_0 <= 8'h0;
      buffers_1 <= 8'h0;
    end else begin
      buffers_0 <= io_dataIn;
      buffers_1 <= buffers_0;
    end
  end


endmodule

module BufferCC_2 (
  input  wire [1:0]    io_dataIn,
  output wire [1:0]    io_dataOut,
  input  wire          clk_ram_bus,
  input  wire          ram_axi_cc_toplevel_board_ctrl_reset_cpu_synchronized
);

  (* async_reg = "true" *) reg        [1:0]    buffers_0;
  (* async_reg = "true" *) reg        [1:0]    buffers_1;

  assign io_dataOut = buffers_1;
  always @(posedge clk_ram_bus or posedge ram_axi_cc_toplevel_board_ctrl_reset_cpu_synchronized) begin
    if(ram_axi_cc_toplevel_board_ctrl_reset_cpu_synchronized) begin
      buffers_0 <= 2'b00;
      buffers_1 <= 2'b00;
    end else begin
      buffers_0 <= io_dataIn;
      buffers_1 <= buffers_0;
    end
  end


endmodule

module BufferCC_1 (
  input  wire          io_dataIn,
  output wire          io_dataOut,
  input  wire          clk_ram_bus,
  input  wire          reset_cpu
);

  (* async_reg = "true" *) reg                 buffers_0;
  (* async_reg = "true" *) reg                 buffers_1;

  assign io_dataOut = buffers_1;
  always @(posedge clk_ram_bus or posedge reset_cpu) begin
    if(reset_cpu) begin
      buffers_0 <= 1'b1;
      buffers_1 <= 1'b1;
    end else begin
      buffers_0 <= io_dataIn;
      buffers_1 <= buffers_0;
    end
  end


endmodule

module BufferCC (
  input  wire [1:0]    io_dataIn,
  output wire [1:0]    io_dataOut,
  input  wire          clk_cpu,
  input  wire          reset_cpu
);

  (* async_reg = "true" *) reg        [1:0]    buffers_0;
  (* async_reg = "true" *) reg        [1:0]    buffers_1;

  assign io_dataOut = buffers_1;
  always @(posedge clk_cpu or posedge reset_cpu) begin
    if(reset_cpu) begin
      buffers_0 <= 2'b00;
      buffers_1 <= 2'b00;
    end else begin
      buffers_0 <= io_dataIn;
      buffers_1 <= buffers_0;
    end
  end


endmodule

module RamSyncMwMux (
  input  wire          io_writes_0_valid,
  input  wire [4:0]    io_writes_0_payload_address,
  input  wire [31:0]   io_writes_0_payload_data,
  input  wire          io_writes_1_valid,
  input  wire [4:0]    io_writes_1_payload_address,
  input  wire [31:0]   io_writes_1_payload_data,
  input  wire          io_read_0_cmd_valid,
  input  wire [4:0]    io_read_0_cmd_payload,
  output wire [31:0]   io_read_0_rsp,
  input  wire          io_read_1_cmd_valid,
  input  wire [4:0]    io_read_1_cmd_payload,
  output wire [31:0]   io_read_1_rsp,
  input  wire          io_read_2_cmd_valid,
  input  wire [4:0]    io_read_2_cmd_payload,
  output wire [31:0]   io_read_2_rsp,
  input  wire          io_read_3_cmd_valid,
  input  wire [4:0]    io_read_3_cmd_payload,
  output wire [31:0]   io_read_3_rsp,
  input  wire          clk_cpu,
  input  wire          reset_cpu
);

  reg        [31:0]   ram_0_spinal_port1;
  reg        [31:0]   ram_0_spinal_port2;
  reg        [31:0]   ram_0_spinal_port3;
  reg        [31:0]   ram_0_spinal_port4;
  reg        [31:0]   ram_1_spinal_port1;
  reg        [31:0]   ram_1_spinal_port2;
  reg        [31:0]   ram_1_spinal_port3;
  reg        [31:0]   ram_1_spinal_port4;
  wire       [0:0]    location_io_read_0_rsp;
  wire       [0:0]    location_io_read_1_rsp;
  wire       [0:0]    location_io_read_2_rsp;
  wire       [0:0]    location_io_read_3_rsp;
  reg        [31:0]   _zz_io_read_0_rsp;
  reg        [31:0]   _zz_io_read_1_rsp;
  reg        [31:0]   _zz_io_read_2_rsp;
  reg        [31:0]   _zz_io_read_3_rsp;
  wire       [31:0]   reads_0_reads_0;
  wire       [31:0]   reads_0_reads_1;
  reg        [4:0]    reads_0_addressReg;
  wire       [31:0]   reads_1_reads_0;
  wire       [31:0]   reads_1_reads_1;
  reg        [4:0]    reads_1_addressReg;
  wire       [31:0]   reads_2_reads_0;
  wire       [31:0]   reads_2_reads_1;
  reg        [4:0]    reads_2_addressReg;
  wire       [31:0]   reads_3_reads_0;
  wire       [31:0]   reads_3_reads_1;
  reg        [4:0]    reads_3_addressReg;
  reg [31:0] ram_0 [0:31];
  reg [31:0] ram_1 [0:31];

  always @(posedge clk_cpu) begin
    if(io_writes_0_valid) begin
      ram_0[io_writes_0_payload_address] <= io_writes_0_payload_data;
    end
  end

  always @(posedge clk_cpu) begin
    if(io_read_0_cmd_valid) begin
      ram_0_spinal_port1 <= ram_0[io_read_0_cmd_payload];
    end
  end

  always @(posedge clk_cpu) begin
    if(io_read_1_cmd_valid) begin
      ram_0_spinal_port2 <= ram_0[io_read_1_cmd_payload];
    end
  end

  always @(posedge clk_cpu) begin
    if(io_read_2_cmd_valid) begin
      ram_0_spinal_port3 <= ram_0[io_read_2_cmd_payload];
    end
  end

  always @(posedge clk_cpu) begin
    if(io_read_3_cmd_valid) begin
      ram_0_spinal_port4 <= ram_0[io_read_3_cmd_payload];
    end
  end

  always @(posedge clk_cpu) begin
    if(io_writes_1_valid) begin
      ram_1[io_writes_1_payload_address] <= io_writes_1_payload_data;
    end
  end

  always @(posedge clk_cpu) begin
    if(io_read_0_cmd_valid) begin
      ram_1_spinal_port1 <= ram_1[io_read_0_cmd_payload];
    end
  end

  always @(posedge clk_cpu) begin
    if(io_read_1_cmd_valid) begin
      ram_1_spinal_port2 <= ram_1[io_read_1_cmd_payload];
    end
  end

  always @(posedge clk_cpu) begin
    if(io_read_2_cmd_valid) begin
      ram_1_spinal_port3 <= ram_1[io_read_2_cmd_payload];
    end
  end

  always @(posedge clk_cpu) begin
    if(io_read_3_cmd_valid) begin
      ram_1_spinal_port4 <= ram_1[io_read_3_cmd_payload];
    end
  end

  RamAsyncMwReg location (
    .io_writes_0_valid           (io_writes_0_valid               ), //i
    .io_writes_0_payload_address (io_writes_0_payload_address[4:0]), //i
    .io_writes_0_payload_data    (1'b0                            ), //i
    .io_writes_1_valid           (io_writes_1_valid               ), //i
    .io_writes_1_payload_address (io_writes_1_payload_address[4:0]), //i
    .io_writes_1_payload_data    (1'b1                            ), //i
    .io_read_0_cmd_valid         (1'b1                            ), //i
    .io_read_0_cmd_payload       (reads_0_addressReg[4:0]         ), //i
    .io_read_0_rsp               (location_io_read_0_rsp          ), //o
    .io_read_1_cmd_valid         (1'b1                            ), //i
    .io_read_1_cmd_payload       (reads_1_addressReg[4:0]         ), //i
    .io_read_1_rsp               (location_io_read_1_rsp          ), //o
    .io_read_2_cmd_valid         (1'b1                            ), //i
    .io_read_2_cmd_payload       (reads_2_addressReg[4:0]         ), //i
    .io_read_2_rsp               (location_io_read_2_rsp          ), //o
    .io_read_3_cmd_valid         (1'b1                            ), //i
    .io_read_3_cmd_payload       (reads_3_addressReg[4:0]         ), //i
    .io_read_3_rsp               (location_io_read_3_rsp          ), //o
    .clk_cpu                     (clk_cpu                         ), //i
    .reset_cpu                   (reset_cpu                       )  //i
  );
  always @(*) begin
    case(location_io_read_0_rsp)
      1'b0 : _zz_io_read_0_rsp = reads_0_reads_0;
      default : _zz_io_read_0_rsp = reads_0_reads_1;
    endcase
  end

  always @(*) begin
    case(location_io_read_1_rsp)
      1'b0 : _zz_io_read_1_rsp = reads_1_reads_0;
      default : _zz_io_read_1_rsp = reads_1_reads_1;
    endcase
  end

  always @(*) begin
    case(location_io_read_2_rsp)
      1'b0 : _zz_io_read_2_rsp = reads_2_reads_0;
      default : _zz_io_read_2_rsp = reads_2_reads_1;
    endcase
  end

  always @(*) begin
    case(location_io_read_3_rsp)
      1'b0 : _zz_io_read_3_rsp = reads_3_reads_0;
      default : _zz_io_read_3_rsp = reads_3_reads_1;
    endcase
  end

  assign reads_0_reads_0 = ram_0_spinal_port1;
  assign reads_0_reads_1 = ram_1_spinal_port1;
  assign io_read_0_rsp = _zz_io_read_0_rsp;
  assign reads_1_reads_0 = ram_0_spinal_port2;
  assign reads_1_reads_1 = ram_1_spinal_port2;
  assign io_read_1_rsp = _zz_io_read_1_rsp;
  assign reads_2_reads_0 = ram_0_spinal_port3;
  assign reads_2_reads_1 = ram_1_spinal_port3;
  assign io_read_2_rsp = _zz_io_read_2_rsp;
  assign reads_3_reads_0 = ram_0_spinal_port4;
  assign reads_3_reads_1 = ram_1_spinal_port4;
  assign io_read_3_rsp = _zz_io_read_3_rsp;
  always @(posedge clk_cpu) begin
    if(io_read_0_cmd_valid) begin
      reads_0_addressReg <= io_read_0_cmd_payload;
    end
    if(io_read_1_cmd_valid) begin
      reads_1_addressReg <= io_read_1_cmd_payload;
    end
    if(io_read_2_cmd_valid) begin
      reads_2_addressReg <= io_read_2_cmd_payload;
    end
    if(io_read_3_cmd_valid) begin
      reads_3_addressReg <= io_read_3_cmd_payload;
    end
  end


endmodule

//UsbLsFsPhyFilter_1 replaced by UsbLsFsPhyFilter

module UsbLsFsPhyFilter (
  input  wire          io_lowSpeed,
  input  wire          io_usb_dp,
  input  wire          io_usb_dm,
  output wire          io_filtred_dp,
  output wire          io_filtred_dm,
  output wire          io_filtred_d,
  output wire          io_filtred_se0,
  output wire          io_filtred_sample,
  input  wire          clk_peripheral,
  input  wire          reset_peripheral
);

  wire       [4:0]    _zz_timer_sampleDo;
  reg                 timer_clear;
  reg        [4:0]    timer_counter;
  wire       [4:0]    timer_counterLimit;
  wire                when_UsbHubPhy_l98;
  wire       [3:0]    timer_sampleAt;
  wire                timer_sampleDo;
  reg                 io_usb_dp_regNext;
  reg                 io_usb_dm_regNext;
  wire                when_UsbHubPhy_l105;

  assign _zz_timer_sampleDo = {1'd0, timer_sampleAt};
  always @(*) begin
    timer_clear = 1'b0;
    if(when_UsbHubPhy_l105) begin
      timer_clear = 1'b1;
    end
  end

  assign timer_counterLimit = (io_lowSpeed ? 5'h1f : 5'h03);
  assign when_UsbHubPhy_l98 = ((timer_counter == timer_counterLimit) || timer_clear);
  assign timer_sampleAt = (io_lowSpeed ? 4'b1110 : 4'b0000);
  assign timer_sampleDo = ((timer_counter == _zz_timer_sampleDo) && (! timer_clear));
  assign when_UsbHubPhy_l105 = ((io_usb_dp ^ io_usb_dp_regNext) || (io_usb_dm ^ io_usb_dm_regNext));
  assign io_filtred_dp = io_usb_dp;
  assign io_filtred_dm = io_usb_dm;
  assign io_filtred_d = io_usb_dp;
  assign io_filtred_sample = timer_sampleDo;
  assign io_filtred_se0 = ((! io_usb_dp) && (! io_usb_dm));
  always @(posedge clk_peripheral) begin
    timer_counter <= (timer_counter + 5'h01);
    if(when_UsbHubPhy_l98) begin
      timer_counter <= 5'h0;
    end
    io_usb_dp_regNext <= io_usb_dp;
    io_usb_dm_regNext <= io_usb_dm;
  end


endmodule

module Crc_2 (
  input  wire          io_flush,
  input  wire          io_input_valid,
  input  wire [7:0]    io_input_payload,
  output wire [15:0]   io_result,
  output wire [15:0]   io_resultNext,
  input  wire          clk_peripheral,
  input  wire          reset_peripheral
);

  wire       [15:0]   _zz_acc_1;
  wire       [15:0]   _zz_acc_2;
  wire       [15:0]   _zz_acc_3;
  wire       [15:0]   _zz_acc_4;
  wire       [15:0]   _zz_acc_5;
  wire       [15:0]   _zz_acc_6;
  wire       [15:0]   _zz_acc_7;
  wire       [15:0]   _zz_acc_8;
  reg        [15:0]   acc_8;
  reg        [15:0]   acc_7;
  reg        [15:0]   acc_6;
  reg        [15:0]   acc_5;
  reg        [15:0]   acc_4;
  reg        [15:0]   acc_3;
  reg        [15:0]   acc_2;
  reg        [15:0]   acc_1;
  reg        [15:0]   state;
  wire       [15:0]   acc;
  wire       [15:0]   stateXor;
  wire       [15:0]   accXor;

  assign _zz_acc_1 = (acc <<< 1);
  assign _zz_acc_2 = (acc_1 <<< 1);
  assign _zz_acc_3 = (acc_2 <<< 1);
  assign _zz_acc_4 = (acc_3 <<< 1);
  assign _zz_acc_5 = (acc_4 <<< 1);
  assign _zz_acc_6 = (acc_5 <<< 1);
  assign _zz_acc_7 = (acc_6 <<< 1);
  assign _zz_acc_8 = (acc_7 <<< 1);
  always @(*) begin
    acc_8 = acc_7;
    acc_8 = (_zz_acc_8 ^ ((io_input_payload[7] ^ acc_7[15]) ? 16'h8005 : 16'h0));
  end

  always @(*) begin
    acc_7 = acc_6;
    acc_7 = (_zz_acc_7 ^ ((io_input_payload[6] ^ acc_6[15]) ? 16'h8005 : 16'h0));
  end

  always @(*) begin
    acc_6 = acc_5;
    acc_6 = (_zz_acc_6 ^ ((io_input_payload[5] ^ acc_5[15]) ? 16'h8005 : 16'h0));
  end

  always @(*) begin
    acc_5 = acc_4;
    acc_5 = (_zz_acc_5 ^ ((io_input_payload[4] ^ acc_4[15]) ? 16'h8005 : 16'h0));
  end

  always @(*) begin
    acc_4 = acc_3;
    acc_4 = (_zz_acc_4 ^ ((io_input_payload[3] ^ acc_3[15]) ? 16'h8005 : 16'h0));
  end

  always @(*) begin
    acc_3 = acc_2;
    acc_3 = (_zz_acc_3 ^ ((io_input_payload[2] ^ acc_2[15]) ? 16'h8005 : 16'h0));
  end

  always @(*) begin
    acc_2 = acc_1;
    acc_2 = (_zz_acc_2 ^ ((io_input_payload[1] ^ acc_1[15]) ? 16'h8005 : 16'h0));
  end

  always @(*) begin
    acc_1 = acc;
    acc_1 = (_zz_acc_1 ^ ((io_input_payload[0] ^ acc[15]) ? 16'h8005 : 16'h0));
  end

  assign acc = state;
  assign stateXor = (state ^ 16'h0);
  assign accXor = (acc_8 ^ 16'h0);
  assign io_result = stateXor;
  assign io_resultNext = accXor;
  always @(posedge clk_peripheral or posedge reset_peripheral) begin
    if(reset_peripheral) begin
      state <= 16'hffff;
    end else begin
      if(io_input_valid) begin
        state <= acc_8;
      end
      if(io_flush) begin
        state <= 16'hffff;
      end
    end
  end


endmodule

module Crc_1 (
  input  wire          io_flush,
  input  wire          io_input_valid,
  input  wire [7:0]    io_input_payload,
  output wire [15:0]   io_result,
  output wire [15:0]   io_resultNext,
  input  wire          clk_peripheral,
  input  wire          reset_peripheral
);

  wire       [15:0]   _zz_acc_1;
  wire       [15:0]   _zz_acc_2;
  wire       [15:0]   _zz_acc_3;
  wire       [15:0]   _zz_acc_4;
  wire       [15:0]   _zz_acc_5;
  wire       [15:0]   _zz_acc_6;
  wire       [15:0]   _zz_acc_7;
  wire       [15:0]   _zz_acc_8;
  wire                _zz_io_result;
  wire       [0:0]    _zz_io_result_1;
  wire       [6:0]    _zz_io_result_2;
  wire                _zz_io_resultNext;
  wire       [0:0]    _zz_io_resultNext_1;
  wire       [6:0]    _zz_io_resultNext_2;
  reg        [15:0]   acc_8;
  reg        [15:0]   acc_7;
  reg        [15:0]   acc_6;
  reg        [15:0]   acc_5;
  reg        [15:0]   acc_4;
  reg        [15:0]   acc_3;
  reg        [15:0]   acc_2;
  reg        [15:0]   acc_1;
  reg        [15:0]   state;
  wire       [15:0]   acc;
  wire       [15:0]   stateXor;
  wire       [15:0]   accXor;

  assign _zz_acc_1 = (acc <<< 1);
  assign _zz_acc_2 = (acc_1 <<< 1);
  assign _zz_acc_3 = (acc_2 <<< 1);
  assign _zz_acc_4 = (acc_3 <<< 1);
  assign _zz_acc_5 = (acc_4 <<< 1);
  assign _zz_acc_6 = (acc_5 <<< 1);
  assign _zz_acc_7 = (acc_6 <<< 1);
  assign _zz_acc_8 = (acc_7 <<< 1);
  assign _zz_io_result = stateXor[7];
  assign _zz_io_result_1 = stateXor[8];
  assign _zz_io_result_2 = {stateXor[9],{stateXor[10],{stateXor[11],{stateXor[12],{stateXor[13],{stateXor[14],stateXor[15]}}}}}};
  assign _zz_io_resultNext = accXor[7];
  assign _zz_io_resultNext_1 = accXor[8];
  assign _zz_io_resultNext_2 = {accXor[9],{accXor[10],{accXor[11],{accXor[12],{accXor[13],{accXor[14],accXor[15]}}}}}};
  always @(*) begin
    acc_8 = acc_7;
    acc_8 = (_zz_acc_8 ^ ((io_input_payload[7] ^ acc_7[15]) ? 16'h8005 : 16'h0));
  end

  always @(*) begin
    acc_7 = acc_6;
    acc_7 = (_zz_acc_7 ^ ((io_input_payload[6] ^ acc_6[15]) ? 16'h8005 : 16'h0));
  end

  always @(*) begin
    acc_6 = acc_5;
    acc_6 = (_zz_acc_6 ^ ((io_input_payload[5] ^ acc_5[15]) ? 16'h8005 : 16'h0));
  end

  always @(*) begin
    acc_5 = acc_4;
    acc_5 = (_zz_acc_5 ^ ((io_input_payload[4] ^ acc_4[15]) ? 16'h8005 : 16'h0));
  end

  always @(*) begin
    acc_4 = acc_3;
    acc_4 = (_zz_acc_4 ^ ((io_input_payload[3] ^ acc_3[15]) ? 16'h8005 : 16'h0));
  end

  always @(*) begin
    acc_3 = acc_2;
    acc_3 = (_zz_acc_3 ^ ((io_input_payload[2] ^ acc_2[15]) ? 16'h8005 : 16'h0));
  end

  always @(*) begin
    acc_2 = acc_1;
    acc_2 = (_zz_acc_2 ^ ((io_input_payload[1] ^ acc_1[15]) ? 16'h8005 : 16'h0));
  end

  always @(*) begin
    acc_1 = acc;
    acc_1 = (_zz_acc_1 ^ ((io_input_payload[0] ^ acc[15]) ? 16'h8005 : 16'h0));
  end

  assign acc = state;
  assign stateXor = (state ^ 16'hffff);
  assign accXor = (acc_8 ^ 16'hffff);
  assign io_result = {stateXor[0],{stateXor[1],{stateXor[2],{stateXor[3],{stateXor[4],{stateXor[5],{stateXor[6],{_zz_io_result,{_zz_io_result_1,_zz_io_result_2}}}}}}}}};
  assign io_resultNext = {accXor[0],{accXor[1],{accXor[2],{accXor[3],{accXor[4],{accXor[5],{accXor[6],{_zz_io_resultNext,{_zz_io_resultNext_1,_zz_io_resultNext_2}}}}}}}}};
  always @(posedge clk_peripheral or posedge reset_peripheral) begin
    if(reset_peripheral) begin
      state <= 16'hffff;
    end else begin
      if(io_input_valid) begin
        state <= acc_8;
      end
      if(io_flush) begin
        state <= 16'hffff;
      end
    end
  end


endmodule

module Crc (
  input  wire          io_flush,
  input  wire          io_input_valid,
  input  wire [10:0]   io_input_payload,
  output wire [4:0]    io_result,
  output wire [4:0]    io_resultNext,
  input  wire          clk_peripheral,
  input  wire          reset_peripheral
);

  wire       [4:0]    _zz_acc_1;
  wire       [4:0]    _zz_acc_2;
  wire       [4:0]    _zz_acc_3;
  wire       [4:0]    _zz_acc_4;
  wire       [4:0]    _zz_acc_5;
  wire       [4:0]    _zz_acc_6;
  wire       [4:0]    _zz_acc_7;
  wire       [4:0]    _zz_acc_8;
  wire       [4:0]    _zz_acc_9;
  wire       [4:0]    _zz_acc_10;
  wire       [4:0]    _zz_acc_11;
  reg        [4:0]    acc_11;
  reg        [4:0]    acc_10;
  reg        [4:0]    acc_9;
  reg        [4:0]    acc_8;
  reg        [4:0]    acc_7;
  reg        [4:0]    acc_6;
  reg        [4:0]    acc_5;
  reg        [4:0]    acc_4;
  reg        [4:0]    acc_3;
  reg        [4:0]    acc_2;
  reg        [4:0]    acc_1;
  reg        [4:0]    state;
  wire       [4:0]    acc;
  wire       [4:0]    stateXor;
  wire       [4:0]    accXor;

  assign _zz_acc_1 = (acc <<< 1);
  assign _zz_acc_2 = (acc_1 <<< 1);
  assign _zz_acc_3 = (acc_2 <<< 1);
  assign _zz_acc_4 = (acc_3 <<< 1);
  assign _zz_acc_5 = (acc_4 <<< 1);
  assign _zz_acc_6 = (acc_5 <<< 1);
  assign _zz_acc_7 = (acc_6 <<< 1);
  assign _zz_acc_8 = (acc_7 <<< 1);
  assign _zz_acc_9 = (acc_8 <<< 1);
  assign _zz_acc_10 = (acc_9 <<< 1);
  assign _zz_acc_11 = (acc_10 <<< 1);
  always @(*) begin
    acc_11 = acc_10;
    acc_11 = (_zz_acc_11 ^ ((io_input_payload[10] ^ acc_10[4]) ? 5'h05 : 5'h0));
  end

  always @(*) begin
    acc_10 = acc_9;
    acc_10 = (_zz_acc_10 ^ ((io_input_payload[9] ^ acc_9[4]) ? 5'h05 : 5'h0));
  end

  always @(*) begin
    acc_9 = acc_8;
    acc_9 = (_zz_acc_9 ^ ((io_input_payload[8] ^ acc_8[4]) ? 5'h05 : 5'h0));
  end

  always @(*) begin
    acc_8 = acc_7;
    acc_8 = (_zz_acc_8 ^ ((io_input_payload[7] ^ acc_7[4]) ? 5'h05 : 5'h0));
  end

  always @(*) begin
    acc_7 = acc_6;
    acc_7 = (_zz_acc_7 ^ ((io_input_payload[6] ^ acc_6[4]) ? 5'h05 : 5'h0));
  end

  always @(*) begin
    acc_6 = acc_5;
    acc_6 = (_zz_acc_6 ^ ((io_input_payload[5] ^ acc_5[4]) ? 5'h05 : 5'h0));
  end

  always @(*) begin
    acc_5 = acc_4;
    acc_5 = (_zz_acc_5 ^ ((io_input_payload[4] ^ acc_4[4]) ? 5'h05 : 5'h0));
  end

  always @(*) begin
    acc_4 = acc_3;
    acc_4 = (_zz_acc_4 ^ ((io_input_payload[3] ^ acc_3[4]) ? 5'h05 : 5'h0));
  end

  always @(*) begin
    acc_3 = acc_2;
    acc_3 = (_zz_acc_3 ^ ((io_input_payload[2] ^ acc_2[4]) ? 5'h05 : 5'h0));
  end

  always @(*) begin
    acc_2 = acc_1;
    acc_2 = (_zz_acc_2 ^ ((io_input_payload[1] ^ acc_1[4]) ? 5'h05 : 5'h0));
  end

  always @(*) begin
    acc_1 = acc;
    acc_1 = (_zz_acc_1 ^ ((io_input_payload[0] ^ acc[4]) ? 5'h05 : 5'h0));
  end

  assign acc = state;
  assign stateXor = (state ^ 5'h1f);
  assign accXor = (acc_11 ^ 5'h1f);
  assign io_result = {stateXor[0],{stateXor[1],{stateXor[2],{stateXor[3],stateXor[4]}}}};
  assign io_resultNext = {accXor[0],{accXor[1],{accXor[2],{accXor[3],accXor[4]}}}};
  always @(posedge clk_peripheral or posedge reset_peripheral) begin
    if(reset_peripheral) begin
      state <= 5'h1f;
    end else begin
      if(io_input_valid) begin
        state <= acc_11;
      end
      if(io_flush) begin
        state <= 5'h1f;
      end
    end
  end


endmodule

module RamAsyncMwReg (
  input  wire          io_writes_0_valid,
  input  wire [4:0]    io_writes_0_payload_address,
  input  wire [0:0]    io_writes_0_payload_data,
  input  wire          io_writes_1_valid,
  input  wire [4:0]    io_writes_1_payload_address,
  input  wire [0:0]    io_writes_1_payload_data,
  input  wire          io_read_0_cmd_valid,
  input  wire [4:0]    io_read_0_cmd_payload,
  output wire [0:0]    io_read_0_rsp,
  input  wire          io_read_1_cmd_valid,
  input  wire [4:0]    io_read_1_cmd_payload,
  output wire [0:0]    io_read_1_rsp,
  input  wire          io_read_2_cmd_valid,
  input  wire [4:0]    io_read_2_cmd_payload,
  output wire [0:0]    io_read_2_rsp,
  input  wire          io_read_3_cmd_valid,
  input  wire [4:0]    io_read_3_cmd_payload,
  output wire [0:0]    io_read_3_rsp,
  input  wire          clk_cpu,
  input  wire          reset_cpu
);

  reg        [0:0]    _zz_io_read_0_rsp;
  reg        [0:0]    _zz_io_read_1_rsp;
  reg        [0:0]    _zz_io_read_2_rsp;
  reg        [0:0]    _zz_io_read_3_rsp;
  reg        [0:0]    ram_0;
  reg        [0:0]    ram_1;
  reg        [0:0]    ram_2;
  reg        [0:0]    ram_3;
  reg        [0:0]    ram_4;
  reg        [0:0]    ram_5;
  reg        [0:0]    ram_6;
  reg        [0:0]    ram_7;
  reg        [0:0]    ram_8;
  reg        [0:0]    ram_9;
  reg        [0:0]    ram_10;
  reg        [0:0]    ram_11;
  reg        [0:0]    ram_12;
  reg        [0:0]    ram_13;
  reg        [0:0]    ram_14;
  reg        [0:0]    ram_15;
  reg        [0:0]    ram_16;
  reg        [0:0]    ram_17;
  reg        [0:0]    ram_18;
  reg        [0:0]    ram_19;
  reg        [0:0]    ram_20;
  reg        [0:0]    ram_21;
  reg        [0:0]    ram_22;
  reg        [0:0]    ram_23;
  reg        [0:0]    ram_24;
  reg        [0:0]    ram_25;
  reg        [0:0]    ram_26;
  reg        [0:0]    ram_27;
  reg        [0:0]    ram_28;
  reg        [0:0]    ram_29;
  reg        [0:0]    ram_30;
  reg        [0:0]    ram_31;
  wire       [31:0]   _zz_1;
  wire       [0:0]    _zz_ram_0;
  wire       [31:0]   _zz_2;
  wire       [0:0]    _zz_ram_0_1;

  initial begin
  `ifndef SYNTHESIS
    ram_0 = {$urandom};
    ram_1 = {$urandom};
    ram_2 = {$urandom};
    ram_3 = {$urandom};
    ram_4 = {$urandom};
    ram_5 = {$urandom};
    ram_6 = {$urandom};
    ram_7 = {$urandom};
    ram_8 = {$urandom};
    ram_9 = {$urandom};
    ram_10 = {$urandom};
    ram_11 = {$urandom};
    ram_12 = {$urandom};
    ram_13 = {$urandom};
    ram_14 = {$urandom};
    ram_15 = {$urandom};
    ram_16 = {$urandom};
    ram_17 = {$urandom};
    ram_18 = {$urandom};
    ram_19 = {$urandom};
    ram_20 = {$urandom};
    ram_21 = {$urandom};
    ram_22 = {$urandom};
    ram_23 = {$urandom};
    ram_24 = {$urandom};
    ram_25 = {$urandom};
    ram_26 = {$urandom};
    ram_27 = {$urandom};
    ram_28 = {$urandom};
    ram_29 = {$urandom};
    ram_30 = {$urandom};
    ram_31 = {$urandom};
  `endif
  end

  always @(*) begin
    case(io_read_0_cmd_payload)
      5'b00000 : _zz_io_read_0_rsp = ram_0;
      5'b00001 : _zz_io_read_0_rsp = ram_1;
      5'b00010 : _zz_io_read_0_rsp = ram_2;
      5'b00011 : _zz_io_read_0_rsp = ram_3;
      5'b00100 : _zz_io_read_0_rsp = ram_4;
      5'b00101 : _zz_io_read_0_rsp = ram_5;
      5'b00110 : _zz_io_read_0_rsp = ram_6;
      5'b00111 : _zz_io_read_0_rsp = ram_7;
      5'b01000 : _zz_io_read_0_rsp = ram_8;
      5'b01001 : _zz_io_read_0_rsp = ram_9;
      5'b01010 : _zz_io_read_0_rsp = ram_10;
      5'b01011 : _zz_io_read_0_rsp = ram_11;
      5'b01100 : _zz_io_read_0_rsp = ram_12;
      5'b01101 : _zz_io_read_0_rsp = ram_13;
      5'b01110 : _zz_io_read_0_rsp = ram_14;
      5'b01111 : _zz_io_read_0_rsp = ram_15;
      5'b10000 : _zz_io_read_0_rsp = ram_16;
      5'b10001 : _zz_io_read_0_rsp = ram_17;
      5'b10010 : _zz_io_read_0_rsp = ram_18;
      5'b10011 : _zz_io_read_0_rsp = ram_19;
      5'b10100 : _zz_io_read_0_rsp = ram_20;
      5'b10101 : _zz_io_read_0_rsp = ram_21;
      5'b10110 : _zz_io_read_0_rsp = ram_22;
      5'b10111 : _zz_io_read_0_rsp = ram_23;
      5'b11000 : _zz_io_read_0_rsp = ram_24;
      5'b11001 : _zz_io_read_0_rsp = ram_25;
      5'b11010 : _zz_io_read_0_rsp = ram_26;
      5'b11011 : _zz_io_read_0_rsp = ram_27;
      5'b11100 : _zz_io_read_0_rsp = ram_28;
      5'b11101 : _zz_io_read_0_rsp = ram_29;
      5'b11110 : _zz_io_read_0_rsp = ram_30;
      default : _zz_io_read_0_rsp = ram_31;
    endcase
  end

  always @(*) begin
    case(io_read_1_cmd_payload)
      5'b00000 : _zz_io_read_1_rsp = ram_0;
      5'b00001 : _zz_io_read_1_rsp = ram_1;
      5'b00010 : _zz_io_read_1_rsp = ram_2;
      5'b00011 : _zz_io_read_1_rsp = ram_3;
      5'b00100 : _zz_io_read_1_rsp = ram_4;
      5'b00101 : _zz_io_read_1_rsp = ram_5;
      5'b00110 : _zz_io_read_1_rsp = ram_6;
      5'b00111 : _zz_io_read_1_rsp = ram_7;
      5'b01000 : _zz_io_read_1_rsp = ram_8;
      5'b01001 : _zz_io_read_1_rsp = ram_9;
      5'b01010 : _zz_io_read_1_rsp = ram_10;
      5'b01011 : _zz_io_read_1_rsp = ram_11;
      5'b01100 : _zz_io_read_1_rsp = ram_12;
      5'b01101 : _zz_io_read_1_rsp = ram_13;
      5'b01110 : _zz_io_read_1_rsp = ram_14;
      5'b01111 : _zz_io_read_1_rsp = ram_15;
      5'b10000 : _zz_io_read_1_rsp = ram_16;
      5'b10001 : _zz_io_read_1_rsp = ram_17;
      5'b10010 : _zz_io_read_1_rsp = ram_18;
      5'b10011 : _zz_io_read_1_rsp = ram_19;
      5'b10100 : _zz_io_read_1_rsp = ram_20;
      5'b10101 : _zz_io_read_1_rsp = ram_21;
      5'b10110 : _zz_io_read_1_rsp = ram_22;
      5'b10111 : _zz_io_read_1_rsp = ram_23;
      5'b11000 : _zz_io_read_1_rsp = ram_24;
      5'b11001 : _zz_io_read_1_rsp = ram_25;
      5'b11010 : _zz_io_read_1_rsp = ram_26;
      5'b11011 : _zz_io_read_1_rsp = ram_27;
      5'b11100 : _zz_io_read_1_rsp = ram_28;
      5'b11101 : _zz_io_read_1_rsp = ram_29;
      5'b11110 : _zz_io_read_1_rsp = ram_30;
      default : _zz_io_read_1_rsp = ram_31;
    endcase
  end

  always @(*) begin
    case(io_read_2_cmd_payload)
      5'b00000 : _zz_io_read_2_rsp = ram_0;
      5'b00001 : _zz_io_read_2_rsp = ram_1;
      5'b00010 : _zz_io_read_2_rsp = ram_2;
      5'b00011 : _zz_io_read_2_rsp = ram_3;
      5'b00100 : _zz_io_read_2_rsp = ram_4;
      5'b00101 : _zz_io_read_2_rsp = ram_5;
      5'b00110 : _zz_io_read_2_rsp = ram_6;
      5'b00111 : _zz_io_read_2_rsp = ram_7;
      5'b01000 : _zz_io_read_2_rsp = ram_8;
      5'b01001 : _zz_io_read_2_rsp = ram_9;
      5'b01010 : _zz_io_read_2_rsp = ram_10;
      5'b01011 : _zz_io_read_2_rsp = ram_11;
      5'b01100 : _zz_io_read_2_rsp = ram_12;
      5'b01101 : _zz_io_read_2_rsp = ram_13;
      5'b01110 : _zz_io_read_2_rsp = ram_14;
      5'b01111 : _zz_io_read_2_rsp = ram_15;
      5'b10000 : _zz_io_read_2_rsp = ram_16;
      5'b10001 : _zz_io_read_2_rsp = ram_17;
      5'b10010 : _zz_io_read_2_rsp = ram_18;
      5'b10011 : _zz_io_read_2_rsp = ram_19;
      5'b10100 : _zz_io_read_2_rsp = ram_20;
      5'b10101 : _zz_io_read_2_rsp = ram_21;
      5'b10110 : _zz_io_read_2_rsp = ram_22;
      5'b10111 : _zz_io_read_2_rsp = ram_23;
      5'b11000 : _zz_io_read_2_rsp = ram_24;
      5'b11001 : _zz_io_read_2_rsp = ram_25;
      5'b11010 : _zz_io_read_2_rsp = ram_26;
      5'b11011 : _zz_io_read_2_rsp = ram_27;
      5'b11100 : _zz_io_read_2_rsp = ram_28;
      5'b11101 : _zz_io_read_2_rsp = ram_29;
      5'b11110 : _zz_io_read_2_rsp = ram_30;
      default : _zz_io_read_2_rsp = ram_31;
    endcase
  end

  always @(*) begin
    case(io_read_3_cmd_payload)
      5'b00000 : _zz_io_read_3_rsp = ram_0;
      5'b00001 : _zz_io_read_3_rsp = ram_1;
      5'b00010 : _zz_io_read_3_rsp = ram_2;
      5'b00011 : _zz_io_read_3_rsp = ram_3;
      5'b00100 : _zz_io_read_3_rsp = ram_4;
      5'b00101 : _zz_io_read_3_rsp = ram_5;
      5'b00110 : _zz_io_read_3_rsp = ram_6;
      5'b00111 : _zz_io_read_3_rsp = ram_7;
      5'b01000 : _zz_io_read_3_rsp = ram_8;
      5'b01001 : _zz_io_read_3_rsp = ram_9;
      5'b01010 : _zz_io_read_3_rsp = ram_10;
      5'b01011 : _zz_io_read_3_rsp = ram_11;
      5'b01100 : _zz_io_read_3_rsp = ram_12;
      5'b01101 : _zz_io_read_3_rsp = ram_13;
      5'b01110 : _zz_io_read_3_rsp = ram_14;
      5'b01111 : _zz_io_read_3_rsp = ram_15;
      5'b10000 : _zz_io_read_3_rsp = ram_16;
      5'b10001 : _zz_io_read_3_rsp = ram_17;
      5'b10010 : _zz_io_read_3_rsp = ram_18;
      5'b10011 : _zz_io_read_3_rsp = ram_19;
      5'b10100 : _zz_io_read_3_rsp = ram_20;
      5'b10101 : _zz_io_read_3_rsp = ram_21;
      5'b10110 : _zz_io_read_3_rsp = ram_22;
      5'b10111 : _zz_io_read_3_rsp = ram_23;
      5'b11000 : _zz_io_read_3_rsp = ram_24;
      5'b11001 : _zz_io_read_3_rsp = ram_25;
      5'b11010 : _zz_io_read_3_rsp = ram_26;
      5'b11011 : _zz_io_read_3_rsp = ram_27;
      5'b11100 : _zz_io_read_3_rsp = ram_28;
      5'b11101 : _zz_io_read_3_rsp = ram_29;
      5'b11110 : _zz_io_read_3_rsp = ram_30;
      default : _zz_io_read_3_rsp = ram_31;
    endcase
  end

  assign _zz_1 = ({31'd0,1'b1} <<< io_writes_0_payload_address);
  assign _zz_ram_0 = io_writes_0_payload_data;
  assign _zz_2 = ({31'd0,1'b1} <<< io_writes_1_payload_address);
  assign _zz_ram_0_1 = io_writes_1_payload_data;
  assign io_read_0_rsp = _zz_io_read_0_rsp;
  assign io_read_1_rsp = _zz_io_read_1_rsp;
  assign io_read_2_rsp = _zz_io_read_2_rsp;
  assign io_read_3_rsp = _zz_io_read_3_rsp;
  always @(posedge clk_cpu) begin
    if(io_writes_0_valid) begin
      if(_zz_1[0]) begin
        ram_0 <= _zz_ram_0;
      end
      if(_zz_1[1]) begin
        ram_1 <= _zz_ram_0;
      end
      if(_zz_1[2]) begin
        ram_2 <= _zz_ram_0;
      end
      if(_zz_1[3]) begin
        ram_3 <= _zz_ram_0;
      end
      if(_zz_1[4]) begin
        ram_4 <= _zz_ram_0;
      end
      if(_zz_1[5]) begin
        ram_5 <= _zz_ram_0;
      end
      if(_zz_1[6]) begin
        ram_6 <= _zz_ram_0;
      end
      if(_zz_1[7]) begin
        ram_7 <= _zz_ram_0;
      end
      if(_zz_1[8]) begin
        ram_8 <= _zz_ram_0;
      end
      if(_zz_1[9]) begin
        ram_9 <= _zz_ram_0;
      end
      if(_zz_1[10]) begin
        ram_10 <= _zz_ram_0;
      end
      if(_zz_1[11]) begin
        ram_11 <= _zz_ram_0;
      end
      if(_zz_1[12]) begin
        ram_12 <= _zz_ram_0;
      end
      if(_zz_1[13]) begin
        ram_13 <= _zz_ram_0;
      end
      if(_zz_1[14]) begin
        ram_14 <= _zz_ram_0;
      end
      if(_zz_1[15]) begin
        ram_15 <= _zz_ram_0;
      end
      if(_zz_1[16]) begin
        ram_16 <= _zz_ram_0;
      end
      if(_zz_1[17]) begin
        ram_17 <= _zz_ram_0;
      end
      if(_zz_1[18]) begin
        ram_18 <= _zz_ram_0;
      end
      if(_zz_1[19]) begin
        ram_19 <= _zz_ram_0;
      end
      if(_zz_1[20]) begin
        ram_20 <= _zz_ram_0;
      end
      if(_zz_1[21]) begin
        ram_21 <= _zz_ram_0;
      end
      if(_zz_1[22]) begin
        ram_22 <= _zz_ram_0;
      end
      if(_zz_1[23]) begin
        ram_23 <= _zz_ram_0;
      end
      if(_zz_1[24]) begin
        ram_24 <= _zz_ram_0;
      end
      if(_zz_1[25]) begin
        ram_25 <= _zz_ram_0;
      end
      if(_zz_1[26]) begin
        ram_26 <= _zz_ram_0;
      end
      if(_zz_1[27]) begin
        ram_27 <= _zz_ram_0;
      end
      if(_zz_1[28]) begin
        ram_28 <= _zz_ram_0;
      end
      if(_zz_1[29]) begin
        ram_29 <= _zz_ram_0;
      end
      if(_zz_1[30]) begin
        ram_30 <= _zz_ram_0;
      end
      if(_zz_1[31]) begin
        ram_31 <= _zz_ram_0;
      end
    end
    if(io_writes_1_valid) begin
      if(_zz_2[0]) begin
        ram_0 <= _zz_ram_0_1;
      end
      if(_zz_2[1]) begin
        ram_1 <= _zz_ram_0_1;
      end
      if(_zz_2[2]) begin
        ram_2 <= _zz_ram_0_1;
      end
      if(_zz_2[3]) begin
        ram_3 <= _zz_ram_0_1;
      end
      if(_zz_2[4]) begin
        ram_4 <= _zz_ram_0_1;
      end
      if(_zz_2[5]) begin
        ram_5 <= _zz_ram_0_1;
      end
      if(_zz_2[6]) begin
        ram_6 <= _zz_ram_0_1;
      end
      if(_zz_2[7]) begin
        ram_7 <= _zz_ram_0_1;
      end
      if(_zz_2[8]) begin
        ram_8 <= _zz_ram_0_1;
      end
      if(_zz_2[9]) begin
        ram_9 <= _zz_ram_0_1;
      end
      if(_zz_2[10]) begin
        ram_10 <= _zz_ram_0_1;
      end
      if(_zz_2[11]) begin
        ram_11 <= _zz_ram_0_1;
      end
      if(_zz_2[12]) begin
        ram_12 <= _zz_ram_0_1;
      end
      if(_zz_2[13]) begin
        ram_13 <= _zz_ram_0_1;
      end
      if(_zz_2[14]) begin
        ram_14 <= _zz_ram_0_1;
      end
      if(_zz_2[15]) begin
        ram_15 <= _zz_ram_0_1;
      end
      if(_zz_2[16]) begin
        ram_16 <= _zz_ram_0_1;
      end
      if(_zz_2[17]) begin
        ram_17 <= _zz_ram_0_1;
      end
      if(_zz_2[18]) begin
        ram_18 <= _zz_ram_0_1;
      end
      if(_zz_2[19]) begin
        ram_19 <= _zz_ram_0_1;
      end
      if(_zz_2[20]) begin
        ram_20 <= _zz_ram_0_1;
      end
      if(_zz_2[21]) begin
        ram_21 <= _zz_ram_0_1;
      end
      if(_zz_2[22]) begin
        ram_22 <= _zz_ram_0_1;
      end
      if(_zz_2[23]) begin
        ram_23 <= _zz_ram_0_1;
      end
      if(_zz_2[24]) begin
        ram_24 <= _zz_ram_0_1;
      end
      if(_zz_2[25]) begin
        ram_25 <= _zz_ram_0_1;
      end
      if(_zz_2[26]) begin
        ram_26 <= _zz_ram_0_1;
      end
      if(_zz_2[27]) begin
        ram_27 <= _zz_ram_0_1;
      end
      if(_zz_2[28]) begin
        ram_28 <= _zz_ram_0_1;
      end
      if(_zz_2[29]) begin
        ram_29 <= _zz_ram_0_1;
      end
      if(_zz_2[30]) begin
        ram_30 <= _zz_ram_0_1;
      end
      if(_zz_2[31]) begin
        ram_31 <= _zz_ram_0_1;
      end
    end
  end


endmodule
