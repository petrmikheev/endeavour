`timescale 1ns/1ps

`define SIMULATION

module testbench;

  parameter CPU_FREQ = 96_000_000;
  parameter UART_BAUD_RATE = 48_000_000;

  defparam system.clocks.RESET_DELAY = 3;
  defparam system.uart_ctrl.OVERRIDE_DIVISOR = CPU_FREQ / UART_BAUD_RATE - 1;

  reg clk100mhz = 0;
  always #5 clk100mhz = ~clk100mhz;

  wire [2:0] leds;

  reg uart_rx = 1;
  wire uart_tx;

  /*wire [15:0] DDR_DQ;
  wire [1:0]  DDR_DQS;
  wire [12:0] DDR_A;
  wire [1:0]  DDR_BA;
  wire [3:0]  DDR_nCS;
  wire        DDR_CK;
  wire        DDR_nCK;
  wire        DDR_CKE;
  wire        DDR_nWE;
  wire        DDR_nCAS;
  wire        DDR_nRAS;
  wire [1:0]  DDR_DM;*/

  wire SD_CLK;
  wire SD_CMD;
  wire [3:0] SD_DATA;

  pullup(SD_CMD);

  EndeavourSoc system(
    .io_clk100mhz(clk100mhz),
    .io_nreset(1'b1),
    .io_keys(2'b0),
    .io_leds(leds),
    .io_uart_rx(uart_rx),
    .io_uart_tx(uart_tx),
    /*.DDR_DQ(DDR_DQ),
    .DDR_DQS(DDR_DQS),
    .DDR_A(DDR_A),
    .DDR_BA(DDR_BA),
    .DDR_nCS(DDR_nCS),
    .DDR_CK(DDR_CK),
    .DDR_nCK(DDR_nCK),
    .DDR_CKE(DDR_CKE),
    .DDR_nWE(DDR_nWE),
    .DDR_nCAS(DDR_nCAS),
    .DDR_nRAS(DDR_nRAS),
    .DDR_DM(DDR_DM)*/
    .io_sdcard_clk(SD_CLK),
    .io_sdcard_cmd(SD_CMD),
    .io_sdcard_data(SD_DATA)
  );

  mdl_sdio #(.OPT_HIGH_CAPACITY(1'b1)) sdcard(
    .sd_clk(SD_CLK),
    .sd_cmd(SD_CMD),
    .sd_dat(SD_DATA)
  );

  // AS4C32M16D1A
  /*micron_ddr_sdram_model #(
    .DEBUG(0),
    .BA_BITS(2),
    .ROW_BITS(13),
    .COL_BITS(10),
    .DQ_LEVEL(2)*/
/*    .tCK(7.5),     // tCK    ns    Nominal Clock Cycle Time
    .tDQSQ(0.4),   // tDQSQ  ns    DQS-DQ skew, DQS to last DQ valid, per group, per access
    .tMRD(10.0),   // tMRD   ns    Load Mode Register command cycle time
    // .tRAP(?),   // tRAP   ns    ACTIVE to READ with Auto precharge command
    .tRAS(40.0),   // tRAS   ns    Active to Precharge command time
    .tRC(55.0),    // tRC    ns    Active to Active/Auto Refresh command time
    .tRFC(70.0),   // tRFC   ns    Refresh to Refresh Command interval time
    .tRCD(15.0),   // tRCD   ns    Active to Read/Write command time
    .tRP(15.0),    // tRP    ns    Precharge command period
    .tRRD(10.0),   // tRRD   ns    Active bank a to Active bank b command time
    .tWR(15.0)     // tWR    ns    Write recovery time*/
  /*) ram (
    .Clk(DDR_CK), .Clk_n(DDR_nCK), .Cke(DDR_CKE),
    .Cs_n(DDR_nCS[3]),
    .Ras_n(DDR_nRAS), .Cas_n(DDR_nCAS), .We_n(DDR_nWE),
    .Ba(DDR_BA), .Addr(DDR_A),
    .Dm(DDR_DM), .Dq(DDR_DQ), .Dqs(DDR_DQS)
  );*/

  wire [31:0] pc_decode = testbench.system.vexRiscv_1.decode_PC;
  wire [31:0] instr_decode = testbench.system.vexRiscv_1.decode_INSTRUCTION;
  wire [31:0] instr_execute = testbench.system.vexRiscv_1.execute_INSTRUCTION;
  wire [31:0] instr_memory = testbench.system.vexRiscv_1.memory_INSTRUCTION;
  wire [31:0] instr_writeBack = testbench.system.vexRiscv_1.writeBack_INSTRUCTION;

  wire [31:0] reg01_ra = testbench.system.vexRiscv_1.RegFilePlugin_regFile[1];
  wire [31:0] reg02_sp = testbench.system.vexRiscv_1.RegFilePlugin_regFile[2];
  wire [31:0] reg03_gp = testbench.system.vexRiscv_1.RegFilePlugin_regFile[3];
  wire [31:0] reg04_tp = testbench.system.vexRiscv_1.RegFilePlugin_regFile[4];
  wire [31:0] reg05_t0 = testbench.system.vexRiscv_1.RegFilePlugin_regFile[5];
  wire [31:0] reg06_t1 = testbench.system.vexRiscv_1.RegFilePlugin_regFile[6];
  wire [31:0] reg07_t2 = testbench.system.vexRiscv_1.RegFilePlugin_regFile[7];
  wire [31:0] reg08_s0 = testbench.system.vexRiscv_1.RegFilePlugin_regFile[8];
  wire [31:0] reg09_s1 = testbench.system.vexRiscv_1.RegFilePlugin_regFile[9];
  wire [31:0] reg10_a0 = testbench.system.vexRiscv_1.RegFilePlugin_regFile[10];
  wire [31:0] reg11_a1 = testbench.system.vexRiscv_1.RegFilePlugin_regFile[11];
  wire [31:0] reg12_a2 = testbench.system.vexRiscv_1.RegFilePlugin_regFile[12];
  wire [31:0] reg13_a3 = testbench.system.vexRiscv_1.RegFilePlugin_regFile[13];
  wire [31:0] reg14_a4 = testbench.system.vexRiscv_1.RegFilePlugin_regFile[14];
  wire [31:0] reg15_a5 = testbench.system.vexRiscv_1.RegFilePlugin_regFile[15];
  wire [31:0] reg16_a6 = testbench.system.vexRiscv_1.RegFilePlugin_regFile[16];
  wire [31:0] reg17_a7 = testbench.system.vexRiscv_1.RegFilePlugin_regFile[17];
  wire [31:0] reg18_s2 = testbench.system.vexRiscv_1.RegFilePlugin_regFile[18];
  wire [31:0] reg19_s3 = testbench.system.vexRiscv_1.RegFilePlugin_regFile[19];
  wire [31:0] reg20_s4 = testbench.system.vexRiscv_1.RegFilePlugin_regFile[20];
  wire [31:0] reg21_s5 = testbench.system.vexRiscv_1.RegFilePlugin_regFile[21];
  wire [31:0] reg22_s6 = testbench.system.vexRiscv_1.RegFilePlugin_regFile[22];
  wire [31:0] reg23_s7 = testbench.system.vexRiscv_1.RegFilePlugin_regFile[23];
  wire [31:0] reg24_s8 = testbench.system.vexRiscv_1.RegFilePlugin_regFile[24];
  wire [31:0] reg25_s9 = testbench.system.vexRiscv_1.RegFilePlugin_regFile[25];
  wire [31:0] reg26_s10 = testbench.system.vexRiscv_1.RegFilePlugin_regFile[26];
  wire [31:0] reg27_s11 = testbench.system.vexRiscv_1.RegFilePlugin_regFile[27];
  wire [31:0] reg28_t3 = testbench.system.vexRiscv_1.RegFilePlugin_regFile[28];
  wire [31:0] reg29_t4 = testbench.system.vexRiscv_1.RegFilePlugin_regFile[29];
  wire [31:0] reg30_t5 = testbench.system.vexRiscv_1.RegFilePlugin_regFile[30];
  wire [31:0] reg31_t6 = testbench.system.vexRiscv_1.RegFilePlugin_regFile[31];

  integer dump_i;
  initial begin
    $dumpfile("dump.vcd");
    $dumpvars(0, testbench);
    // cpu registers
    /*$dumpvars(1,
        // cpu instruction
        testbench.system.core.cpu.decode_PC,
        testbench.system.core.cpu.decode_INSTRUCTION,
        testbench.system.core.cpu.execute_INSTRUCTION,
        testbench.system.core.cpu.memory_INSTRUCTION,
        testbench.system.core.cpu.writeBack_INSTRUCTION,
        // cpu io
        testbench.system.core.cpu.dBus_cmd_valid,
        testbench.system.core.cpu.dBus_cmd_ready,
        testbench.system.core.cpu.dBus_cmd_payload_wr,
        testbench.system.core.cpu.dBus_cmd_payload_uncached,
        testbench.system.core.cpu.dBus_cmd_payload_address,
        testbench.system.core.cpu.dBus_cmd_payload_data,
        testbench.system.core.cpu.dBus_cmd_payload_mask,
        testbench.system.core.cpu.dBus_cmd_payload_size,
        testbench.system.core.cpu.dBus_cmd_payload_last,
        testbench.system.core.cpu.dBus_rsp_valid,
        testbench.system.core.cpu.dBus_rsp_payload_last,
        testbench.system.core.cpu.dBus_rsp_payload_data,
        testbench.system.core.cpu.dBus_rsp_payload_error,
        testbench.system.core.cpu.timerInterrupt,
        testbench.system.core.cpu.externalInterrupt,
        testbench.system.core.cpu.softwareInterrupt,
        testbench.system.core.cpu.iBus_cmd_valid,
        testbench.system.core.cpu.iBus_cmd_ready,
        testbench.system.core.cpu.iBus_cmd_payload_address,
        testbench.system.core.cpu.iBus_cmd_payload_size,
        testbench.system.core.cpu.iBus_rsp_valid,
        testbench.system.core.cpu.iBus_rsp_payload_data,
        testbench.system.core.cpu.iBus_rsp_payload_error,*/
        // ram
        /*testbench.system.ram_ctrl.ddr_in,
        testbench.system.ram_ctrl.ddr_out,
        testbench.system.ram_ctrl.stat*/
        //testbench.system.ram_ctrl
    //);

    #4000000;
    $finish;
  end

  // Initialize sdcard content
  integer sdcard_file;
  reg [511:0] sdcard_file_path;
  initial begin
    if ($value$plusargs("sdcard=%s", sdcard_file_path)) begin
      sdcard_file = $fopen(sdcard_file_path, "rb");
      if (!$fread(sdcard.mem, sdcard_file)) $display("Sdcard content initialization failed");
    end
  end

  // Send uart
  integer uart_send_count = 0;
  integer uart_file = -1;
  integer uart_i;
  reg [511:0] uart_file_path;
  initial begin
    if ($value$plusargs("uart=%s", uart_file_path))
      uart_file = $fopen(uart_file_path, "rb");
  end

  reg [7:0] uart_byte;
  localparam UART_BIT_TIME = 1_000_000_000.0 / UART_BAUD_RATE;
  initial begin
    #500000;
    while (uart_file != -1 && !$feof(uart_file)) begin
      uart_send_count = uart_send_count + 1;
      #UART_BIT_TIME;
      uart_rx = 0; #UART_BIT_TIME;
      uart_byte = $fgetc(uart_file);
      for (uart_i = 0; uart_i < 8; uart_i = uart_i + 1) begin
        uart_rx = uart_byte[uart_i]; #UART_BIT_TIME;
      end
      uart_rx = ^uart_byte;
      // if (uart_send_count == 40) uart_rx = ~uart_rx;  // simulate parity error
      #UART_BIT_TIME;  // parity bit
      /*if (uart_send_count == 57) begin  // simulate framing error
        uart_rx = 0;
        #(UART_BIT_TIME*2/3);
      end*/
      uart_rx = 1; #UART_BIT_TIME;
    end
  end

endmodule
